-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Feb 19 2025 19:26:15

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    CMA : out std_logic_vector(10 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__11942\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \N_969_i\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_7_9_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0_cascade_\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_318_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.BANK0_RNOZ0Z_0_cascade_\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.BANK0_RNOZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.N_361_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_344_cascade_\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.N_253_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\ : std_logic;
signal \U712_CHIP_RAM.N_344\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_1\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0_a3_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_345\ : std_logic;
signal \U712_CHIP_RAM.N_71_i\ : std_logic;
signal \U712_CHIP_RAM.N_71_i_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_49\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_3\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_239_i_0_en_cascade_\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \U712_CYCLE_TERM.N_239_i_0_en_0\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.BANK0_RNOZ0Z_1\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_354_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_414_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_5_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_0_a2_i_1_cascade_\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_230_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a3_1_1\ : std_logic;
signal \U712_CHIP_RAM.N_287_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_217\ : std_logic;
signal \U712_CHIP_RAM.N_22\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_113_tz_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3T4KZ0Z7_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_284_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_230\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_271\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_271_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_347\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_1_0\ : std_logic;
signal \U712_REG_SM.N_304\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.N_340\ : std_logic;
signal \U712_REG_SM.N_52\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \C1_c\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_414_0\ : std_logic;
signal \U712_CHIP_RAM.N_363_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_282\ : std_logic;
signal \U712_CHIP_RAM.N_292\ : std_logic;
signal \U712_CHIP_RAM.N_236_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_274\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_366\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a2_2_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a3_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_252_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_286\ : std_logic;
signal \U712_CHIP_RAM.N_267\ : std_logic;
signal \U712_CHIP_RAM.N_225_i\ : std_logic;
signal \U712_CHIP_RAM.N_236\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_i_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.N_234\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_i_o2_0_1_3_cascade_\ : std_logic;
signal \U712_REG_SM.N_272_cascade_\ : std_logic;
signal \U712_REG_SM.N_270_cascade_\ : std_logic;
signal \N_202_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_242\ : std_logic;
signal \N_188_i\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0\ : std_logic;
signal \N_203_i\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0\ : std_logic;
signal \N_186_i\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_243\ : std_logic;
signal \U712_BYTE_ENABLE.N_244\ : std_logic;
signal \U712_BYTE_ENABLE.N_245\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \DMA_LATCH_EN_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_320_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_414\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_1\ : std_logic;
signal \U712_CHIP_RAM.N_48_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_363\ : std_logic;
signal \U712_CHIP_RAM.N_358_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_a3_1\ : std_logic;
signal \U712_CHIP_RAM.N_357\ : std_logic;
signal \U712_CHIP_RAM.N_413\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \A_c_10\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_269_cascade_\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.DS_EN_RNOZ0Z_0\ : std_logic;
signal \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_cascade_\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.N_313\ : std_logic;
signal \U712_REG_SM.N_220\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.STATE_COUNTc_0_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_266\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_222\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_1\ : std_logic;
signal \U712_REG_SM.N_222_cascade_\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_REG_SM.N_241\ : std_logic;
signal \U712_REG_SM.ASn_0_sqmuxa_1\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \N_243_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \WEn_c\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_358\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.N_333\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.N_367\ : std_logic;
signal \U712_REG_SM.N_374\ : std_logic;
signal \U712_REG_SM.N_226\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \N_182\ : std_logic;
signal \DS_ENm\ : std_logic;
signal \N_184\ : std_logic;
signal \N_245_i\ : std_logic;
signal \N_242_i\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \A_c_0\ : std_logic;
signal \N_244_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \CASn_c\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \WRITE_CYCLEm\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \N_268\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    RAMENn <= \RAMENn_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4066\,
            RESETB => \N__7081\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11942\,
            DIN => \N__11941\,
            DOUT => \N__11940\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11942\,
            PADOUT => \N__11941\,
            PADIN => \N__11940\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5056\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11933\,
            DIN => \N__11932\,
            DOUT => \N__11931\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11933\,
            PADOUT => \N__11932\,
            PADIN => \N__11931\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11924\,
            DIN => \N__11923\,
            DOUT => \N__11922\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11924\,
            PADOUT => \N__11923\,
            PADIN => \N__11922\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8020\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11915\,
            DIN => \N__11914\,
            DOUT => \N__11913\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11915\,
            PADOUT => \N__11914\,
            PADIN => \N__11913\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10834\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11906\,
            DIN => \N__11905\,
            DOUT => \N__11904\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11906\,
            PADOUT => \N__11905\,
            PADIN => \N__11904\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11897\,
            DIN => \N__11896\,
            DOUT => \N__11895\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11897\,
            PADOUT => \N__11896\,
            PADIN => \N__11895\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11888\,
            DIN => \N__11887\,
            DOUT => \N__11886\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11888\,
            PADOUT => \N__11887\,
            PADIN => \N__11886\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11879\,
            DIN => \N__11878\,
            DOUT => \N__11877\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11879\,
            PADOUT => \N__11878\,
            PADIN => \N__11877\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11870\,
            DIN => \N__11869\,
            DOUT => \N__11868\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11870\,
            PADOUT => \N__11869\,
            PADIN => \N__11868\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11861\,
            DIN => \N__11860\,
            DOUT => \N__11859\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11861\,
            PADOUT => \N__11860\,
            PADIN => \N__11859\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11852\,
            DIN => \N__11851\,
            DOUT => \N__11850\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11852\,
            PADOUT => \N__11851\,
            PADIN => \N__11850\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8962\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11843\,
            DIN => \N__11842\,
            DOUT => \N__11841\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11843\,
            PADOUT => \N__11842\,
            PADIN => \N__11841\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8545\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11834\,
            DIN => \N__11833\,
            DOUT => \N__11832\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11834\,
            PADOUT => \N__11833\,
            PADIN => \N__11832\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11825\,
            DIN => \N__11824\,
            DOUT => \N__11823\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11825\,
            PADOUT => \N__11824\,
            PADIN => \N__11823\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11816\,
            DIN => \N__11815\,
            DOUT => \N__11814\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11816\,
            PADOUT => \N__11815\,
            PADIN => \N__11814\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11807\,
            DIN => \N__11806\,
            DOUT => \N__11805\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11807\,
            PADOUT => \N__11806\,
            PADIN => \N__11805\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4657\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11798\,
            DIN => \N__11797\,
            DOUT => \N__11796\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11798\,
            PADOUT => \N__11797\,
            PADIN => \N__11796\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11789\,
            DIN => \N__11788\,
            DOUT => \N__11787\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11789\,
            PADOUT => \N__11788\,
            PADIN => \N__11787\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11780\,
            DIN => \N__11779\,
            DOUT => \N__11778\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11780\,
            PADOUT => \N__11779\,
            PADIN => \N__11778\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9061\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11771\,
            DIN => \N__11770\,
            DOUT => \N__11769\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11771\,
            PADOUT => \N__11770\,
            PADIN => \N__11769\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11762\,
            DIN => \N__11761\,
            DOUT => \N__11760\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11762\,
            PADOUT => \N__11761\,
            PADIN => \N__11760\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8038\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11753\,
            DIN => \N__11752\,
            DOUT => \N__11751\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11753\,
            PADOUT => \N__11752\,
            PADIN => \N__11751\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11744\,
            DIN => \N__11743\,
            DOUT => \N__11742\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11744\,
            PADOUT => \N__11743\,
            PADIN => \N__11742\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8530\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11735\,
            DIN => \N__11734\,
            DOUT => \N__11733\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11735\,
            PADOUT => \N__11734\,
            PADIN => \N__11733\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11726\,
            DIN => \N__11725\,
            DOUT => \N__11724\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11726\,
            PADOUT => \N__11725\,
            PADIN => \N__11724\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11717\,
            DIN => \N__11716\,
            DOUT => \N__11715\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11717\,
            PADOUT => \N__11716\,
            PADIN => \N__11715\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11708\,
            DIN => \N__11707\,
            DOUT => \N__11706\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11708\,
            PADOUT => \N__11707\,
            PADIN => \N__11706\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11699\,
            DIN => \N__11698\,
            DOUT => \N__11697\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11699\,
            PADOUT => \N__11698\,
            PADIN => \N__11697\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11690\,
            DIN => \N__11689\,
            DOUT => \N__11688\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11690\,
            PADOUT => \N__11689\,
            PADIN => \N__11688\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6475\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11681\,
            DIN => \N__11680\,
            DOUT => \N__11679\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11681\,
            PADOUT => \N__11680\,
            PADIN => \N__11679\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11672\,
            DIN => \N__11671\,
            DOUT => \N__11670\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11672\,
            PADOUT => \N__11671\,
            PADIN => \N__11670\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11663\,
            DIN => \N__11662\,
            DOUT => \N__11661\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11663\,
            PADOUT => \N__11662\,
            PADIN => \N__11661\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11654\,
            DIN => \N__11653\,
            DOUT => \N__11652\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11654\,
            PADOUT => \N__11653\,
            PADIN => \N__11652\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11645\,
            DIN => \N__11644\,
            DOUT => \N__11643\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11645\,
            PADOUT => \N__11644\,
            PADIN => \N__11643\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11636\,
            DIN => \N__11635\,
            DOUT => \N__11634\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11636\,
            PADOUT => \N__11635\,
            PADIN => \N__11634\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8101\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11627\,
            DIN => \N__11626\,
            DOUT => \N__11625\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11627\,
            PADOUT => \N__11626\,
            PADIN => \N__11625\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4309\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11618\,
            DIN => \N__11617\,
            DOUT => \N__11616\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11618\,
            PADOUT => \N__11617\,
            PADIN => \N__11616\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9339\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11609\,
            DIN => \N__11608\,
            DOUT => \N__11607\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11609\,
            PADOUT => \N__11608\,
            PADIN => \N__11607\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4081\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11600\,
            DIN => \N__11599\,
            DOUT => \N__11598\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11600\,
            PADOUT => \N__11599\,
            PADIN => \N__11598\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11591\,
            DIN => \N__11590\,
            DOUT => \N__11589\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11591\,
            PADOUT => \N__11590\,
            PADIN => \N__11589\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4198\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11582\,
            DIN => \N__11581\,
            DOUT => \N__11580\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11582\,
            PADOUT => \N__11581\,
            PADIN => \N__11580\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7351\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11573\,
            DIN => \N__11572\,
            DOUT => \N__11571\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11573\,
            PADOUT => \N__11572\,
            PADIN => \N__11571\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11564\,
            DIN => \N__11563\,
            DOUT => \N__11562\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11564\,
            PADOUT => \N__11563\,
            PADIN => \N__11562\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11555\,
            DIN => \N__11554\,
            DOUT => \N__11553\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11555\,
            PADOUT => \N__11554\,
            PADIN => \N__11553\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11546\,
            DIN => \N__11545\,
            DOUT => \N__11544\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11546\,
            PADOUT => \N__11545\,
            PADIN => \N__11544\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11537\,
            DIN => \N__11536\,
            DOUT => \N__11535\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11537\,
            PADOUT => \N__11536\,
            PADIN => \N__11535\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11528\,
            DIN => \N__11527\,
            DOUT => \N__11526\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11528\,
            PADOUT => \N__11527\,
            PADIN => \N__11526\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7045\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11519\,
            DIN => \N__11518\,
            DOUT => \N__11517\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11519\,
            PADOUT => \N__11518\,
            PADIN => \N__11517\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11510\,
            DIN => \N__11509\,
            DOUT => \N__11508\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11510\,
            PADOUT => \N__11509\,
            PADIN => \N__11508\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9338\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11501\,
            DIN => \N__11500\,
            DOUT => \N__11499\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11501\,
            PADOUT => \N__11500\,
            PADIN => \N__11499\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8947\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11492\,
            DIN => \N__11491\,
            DOUT => \N__11490\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11492\,
            PADOUT => \N__11491\,
            PADIN => \N__11490\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9964\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11483\,
            DIN => \N__11482\,
            DOUT => \N__11481\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11483\,
            PADOUT => \N__11482\,
            PADIN => \N__11481\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5737\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11474\,
            DIN => \N__11473\,
            DOUT => \N__11472\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11474\,
            PADOUT => \N__11473\,
            PADIN => \N__11472\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8992\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11465\,
            DIN => \N__11464\,
            DOUT => \N__11463\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11465\,
            PADOUT => \N__11464\,
            PADIN => \N__11463\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7222\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11456\,
            DIN => \N__11455\,
            DOUT => \N__11454\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11456\,
            PADOUT => \N__11455\,
            PADIN => \N__11454\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11447\,
            DIN => \N__11446\,
            DOUT => \N__11445\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11447\,
            PADOUT => \N__11446\,
            PADIN => \N__11445\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11438\,
            DIN => \N__11437\,
            DOUT => \N__11436\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11438\,
            PADOUT => \N__11437\,
            PADIN => \N__11436\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5668\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11429\,
            DIN => \N__11428\,
            DOUT => \N__11427\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11429\,
            PADOUT => \N__11428\,
            PADIN => \N__11427\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7066\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11420\,
            DIN => \N__11419\,
            DOUT => \N__11418\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11420\,
            PADOUT => \N__11419\,
            PADIN => \N__11418\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4480\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11411\,
            DIN => \N__11410\,
            DOUT => \N__11409\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11411\,
            PADOUT => \N__11410\,
            PADIN => \N__11409\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5707\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11402\,
            DIN => \N__11401\,
            DOUT => \N__11400\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11402\,
            PADOUT => \N__11401\,
            PADIN => \N__11400\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11393\,
            DIN => \N__11392\,
            DOUT => \N__11391\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11393\,
            PADOUT => \N__11392\,
            PADIN => \N__11391\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11384\,
            DIN => \N__11383\,
            DOUT => \N__11382\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11384\,
            PADOUT => \N__11383\,
            PADIN => \N__11382\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11375\,
            DIN => \N__11374\,
            DOUT => \N__11373\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11375\,
            PADOUT => \N__11374\,
            PADIN => \N__11373\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11366\,
            DIN => \N__11365\,
            DOUT => \N__11364\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11366\,
            PADOUT => \N__11365\,
            PADIN => \N__11364\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7870\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11357\,
            DIN => \N__11356\,
            DOUT => \N__11355\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11357\,
            PADOUT => \N__11356\,
            PADIN => \N__11355\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8167\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11348\,
            DIN => \N__11347\,
            DOUT => \N__11346\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11348\,
            PADOUT => \N__11347\,
            PADIN => \N__11346\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11339\,
            DIN => \N__11338\,
            DOUT => \N__11337\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11339\,
            PADOUT => \N__11338\,
            PADIN => \N__11337\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5770\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11330\,
            DIN => \N__11329\,
            DOUT => \N__11328\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11330\,
            PADOUT => \N__11329\,
            PADIN => \N__11328\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4156\,
            DIN0 => OPEN,
            DOUT0 => \N__4507\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11321\,
            DIN => \N__11320\,
            DOUT => \N__11319\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11321\,
            PADOUT => \N__11320\,
            PADIN => \N__11319\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7027\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11312\,
            DIN => \N__11311\,
            DOUT => \N__11310\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11312\,
            PADOUT => \N__11311\,
            PADIN => \N__11310\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11303\,
            DIN => \N__11302\,
            DOUT => \N__11301\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11303\,
            PADOUT => \N__11302\,
            PADIN => \N__11301\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11294\,
            DIN => \N__11293\,
            DOUT => \N__11292\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11294\,
            PADOUT => \N__11293\,
            PADIN => \N__11292\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5536\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11285\,
            DIN => \N__11284\,
            DOUT => \N__11283\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11285\,
            PADOUT => \N__11284\,
            PADIN => \N__11283\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11276\,
            DIN => \N__11275\,
            DOUT => \N__11274\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11276\,
            PADOUT => \N__11275\,
            PADIN => \N__11274\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11267\,
            DIN => \N__11266\,
            DOUT => \N__11265\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11267\,
            PADOUT => \N__11266\,
            PADIN => \N__11265\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11258\,
            DIN => \N__11257\,
            DOUT => \N__11256\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11258\,
            PADOUT => \N__11257\,
            PADIN => \N__11256\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11249\,
            DIN => \N__11248\,
            DOUT => \N__11247\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11249\,
            PADOUT => \N__11248\,
            PADIN => \N__11247\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7834\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11240\,
            DIN => \N__11239\,
            DOUT => \N__11238\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11240\,
            PADOUT => \N__11239\,
            PADIN => \N__11238\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8608\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11231\,
            DIN => \N__11230\,
            DOUT => \N__11229\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11231\,
            PADOUT => \N__11230\,
            PADIN => \N__11229\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7102\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11222\,
            DIN => \N__11221\,
            DOUT => \N__11220\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11222\,
            PADOUT => \N__11221\,
            PADIN => \N__11220\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4837\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11213\,
            DIN => \N__11212\,
            DOUT => \N__11211\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11213\,
            PADOUT => \N__11212\,
            PADIN => \N__11211\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11204\,
            DIN => \N__11203\,
            DOUT => \N__11202\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11204\,
            PADOUT => \N__11203\,
            PADIN => \N__11202\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11195\,
            DIN => \N__11194\,
            DOUT => \N__11193\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11195\,
            PADOUT => \N__11194\,
            PADIN => \N__11193\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8815\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11186\,
            DIN => \N__11185\,
            DOUT => \N__11184\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11186\,
            PADOUT => \N__11185\,
            PADIN => \N__11184\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11177\,
            DIN => \N__11176\,
            DOUT => \N__11175\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11177\,
            PADOUT => \N__11176\,
            PADIN => \N__11175\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11168\,
            DIN => \N__11167\,
            DOUT => \N__11166\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11168\,
            PADOUT => \N__11167\,
            PADIN => \N__11166\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4363\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11159\,
            DIN => \N__11158\,
            DOUT => \N__11157\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11159\,
            PADOUT => \N__11158\,
            PADIN => \N__11157\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8560\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11150\,
            DIN => \N__11149\,
            DOUT => \N__11148\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11150\,
            PADOUT => \N__11149\,
            PADIN => \N__11148\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9346\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11141\,
            DIN => \N__11140\,
            DOUT => \N__11139\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11141\,
            PADOUT => \N__11140\,
            PADIN => \N__11139\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2709\ : InMux
    port map (
            O => \N__11122\,
            I => \N__11117\
        );

    \I__2708\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11113\
        );

    \I__2707\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11110\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__11117\,
            I => \N__11107\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11104\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__11113\,
            I => \N__11101\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__11110\,
            I => \N__11098\
        );

    \I__2702\ : Span4Mux_v
    port map (
            O => \N__11107\,
            I => \N__11093\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__11104\,
            I => \N__11093\
        );

    \I__2700\ : Span4Mux_v
    port map (
            O => \N__11101\,
            I => \N__11090\
        );

    \I__2699\ : Span4Mux_v
    port map (
            O => \N__11098\,
            I => \N__11087\
        );

    \I__2698\ : Span4Mux_v
    port map (
            O => \N__11093\,
            I => \N__11084\
        );

    \I__2697\ : Sp12to4
    port map (
            O => \N__11090\,
            I => \N__11081\
        );

    \I__2696\ : Sp12to4
    port map (
            O => \N__11087\,
            I => \N__11076\
        );

    \I__2695\ : Sp12to4
    port map (
            O => \N__11084\,
            I => \N__11076\
        );

    \I__2694\ : Span12Mux_h
    port map (
            O => \N__11081\,
            I => \N__11073\
        );

    \I__2693\ : Span12Mux_h
    port map (
            O => \N__11076\,
            I => \N__11070\
        );

    \I__2692\ : Span12Mux_h
    port map (
            O => \N__11073\,
            I => \N__11067\
        );

    \I__2691\ : Span12Mux_v
    port map (
            O => \N__11070\,
            I => \N__11064\
        );

    \I__2690\ : Odrv12
    port map (
            O => \N__11067\,
            I => \RnW_c\
        );

    \I__2689\ : Odrv12
    port map (
            O => \N__11064\,
            I => \RnW_c\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__11059\,
            I => \N__11055\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__11058\,
            I => \N__11052\
        );

    \I__2686\ : InMux
    port map (
            O => \N__11055\,
            I => \N__11043\
        );

    \I__2685\ : InMux
    port map (
            O => \N__11052\,
            I => \N__11043\
        );

    \I__2684\ : InMux
    port map (
            O => \N__11051\,
            I => \N__11040\
        );

    \I__2683\ : InMux
    port map (
            O => \N__11050\,
            I => \N__11037\
        );

    \I__2682\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11032\
        );

    \I__2681\ : InMux
    port map (
            O => \N__11048\,
            I => \N__11032\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__11043\,
            I => \N__11025\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__11040\,
            I => \N__11025\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__11037\,
            I => \N__11025\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11032\,
            I => \N__11022\
        );

    \I__2676\ : Span12Mux_v
    port map (
            O => \N__11025\,
            I => \N__11019\
        );

    \I__2675\ : Span4Mux_h
    port map (
            O => \N__11022\,
            I => \N__11016\
        );

    \I__2674\ : Span12Mux_h
    port map (
            O => \N__11019\,
            I => \N__11013\
        );

    \I__2673\ : Span4Mux_v
    port map (
            O => \N__11016\,
            I => \N__11010\
        );

    \I__2672\ : Odrv12
    port map (
            O => \N__11013\,
            I => \CASUn_c\
        );

    \I__2671\ : Odrv4
    port map (
            O => \N__11010\,
            I => \CASUn_c\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__11005\,
            I => \N__11002\
        );

    \I__2669\ : InMux
    port map (
            O => \N__11002\,
            I => \N__10999\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__10999\,
            I => \N__10996\
        );

    \I__2667\ : Span4Mux_h
    port map (
            O => \N__10996\,
            I => \N__10993\
        );

    \I__2666\ : Span4Mux_h
    port map (
            O => \N__10993\,
            I => \N__10990\
        );

    \I__2665\ : Span4Mux_h
    port map (
            O => \N__10990\,
            I => \N__10986\
        );

    \I__2664\ : InMux
    port map (
            O => \N__10989\,
            I => \N__10983\
        );

    \I__2663\ : Span4Mux_h
    port map (
            O => \N__10986\,
            I => \N__10977\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__10983\,
            I => \N__10977\
        );

    \I__2661\ : CascadeMux
    port map (
            O => \N__10982\,
            I => \N__10970\
        );

    \I__2660\ : Span4Mux_v
    port map (
            O => \N__10977\,
            I => \N__10967\
        );

    \I__2659\ : InMux
    port map (
            O => \N__10976\,
            I => \N__10964\
        );

    \I__2658\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10961\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__10974\,
            I => \N__10956\
        );

    \I__2656\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10951\
        );

    \I__2655\ : InMux
    port map (
            O => \N__10970\,
            I => \N__10951\
        );

    \I__2654\ : Span4Mux_v
    port map (
            O => \N__10967\,
            I => \N__10944\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__10964\,
            I => \N__10944\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__10961\,
            I => \N__10944\
        );

    \I__2651\ : InMux
    port map (
            O => \N__10960\,
            I => \N__10941\
        );

    \I__2650\ : InMux
    port map (
            O => \N__10959\,
            I => \N__10936\
        );

    \I__2649\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10936\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__10951\,
            I => \N__10932\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__10944\,
            I => \N__10927\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__10941\,
            I => \N__10927\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__10936\,
            I => \N__10923\
        );

    \I__2644\ : InMux
    port map (
            O => \N__10935\,
            I => \N__10920\
        );

    \I__2643\ : Span4Mux_v
    port map (
            O => \N__10932\,
            I => \N__10917\
        );

    \I__2642\ : Span4Mux_h
    port map (
            O => \N__10927\,
            I => \N__10914\
        );

    \I__2641\ : InMux
    port map (
            O => \N__10926\,
            I => \N__10911\
        );

    \I__2640\ : Span4Mux_h
    port map (
            O => \N__10923\,
            I => \N__10908\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__10920\,
            I => \WRITE_CYCLEm\
        );

    \I__2638\ : Odrv4
    port map (
            O => \N__10917\,
            I => \WRITE_CYCLEm\
        );

    \I__2637\ : Odrv4
    port map (
            O => \N__10914\,
            I => \WRITE_CYCLEm\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__10911\,
            I => \WRITE_CYCLEm\
        );

    \I__2635\ : Odrv4
    port map (
            O => \N__10908\,
            I => \WRITE_CYCLEm\
        );

    \I__2634\ : InMux
    port map (
            O => \N__10897\,
            I => \N__10894\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__10894\,
            I => \N__10890\
        );

    \I__2632\ : InMux
    port map (
            O => \N__10893\,
            I => \N__10887\
        );

    \I__2631\ : Span4Mux_v
    port map (
            O => \N__10890\,
            I => \N__10880\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__10887\,
            I => \N__10880\
        );

    \I__2629\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10874\
        );

    \I__2628\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10874\
        );

    \I__2627\ : Span4Mux_v
    port map (
            O => \N__10880\,
            I => \N__10871\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__10879\,
            I => \N__10868\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__10874\,
            I => \N__10864\
        );

    \I__2624\ : Span4Mux_v
    port map (
            O => \N__10871\,
            I => \N__10861\
        );

    \I__2623\ : InMux
    port map (
            O => \N__10868\,
            I => \N__10856\
        );

    \I__2622\ : InMux
    port map (
            O => \N__10867\,
            I => \N__10856\
        );

    \I__2621\ : Span12Mux_h
    port map (
            O => \N__10864\,
            I => \N__10853\
        );

    \I__2620\ : Sp12to4
    port map (
            O => \N__10861\,
            I => \N__10850\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__10856\,
            I => \N__10847\
        );

    \I__2618\ : Span12Mux_v
    port map (
            O => \N__10853\,
            I => \N__10844\
        );

    \I__2617\ : Span12Mux_h
    port map (
            O => \N__10850\,
            I => \N__10839\
        );

    \I__2616\ : Span12Mux_v
    port map (
            O => \N__10847\,
            I => \N__10839\
        );

    \I__2615\ : Odrv12
    port map (
            O => \N__10844\,
            I => \CASLn_c\
        );

    \I__2614\ : Odrv12
    port map (
            O => \N__10839\,
            I => \CASLn_c\
        );

    \I__2613\ : IoInMux
    port map (
            O => \N__10834\,
            I => \N__10831\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__10831\,
            I => \N__10828\
        );

    \I__2611\ : IoSpan4Mux
    port map (
            O => \N__10828\,
            I => \N__10825\
        );

    \I__2610\ : Span4Mux_s3_v
    port map (
            O => \N__10825\,
            I => \N__10822\
        );

    \I__2609\ : Span4Mux_v
    port map (
            O => \N__10822\,
            I => \N__10819\
        );

    \I__2608\ : Odrv4
    port map (
            O => \N__10819\,
            I => \N_268\
        );

    \I__2607\ : InMux
    port map (
            O => \N__10816\,
            I => \N__10809\
        );

    \I__2606\ : InMux
    port map (
            O => \N__10815\,
            I => \N__10809\
        );

    \I__2605\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10806\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__10809\,
            I => \N__10803\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__10806\,
            I => \N__10800\
        );

    \I__2602\ : Span4Mux_v
    port map (
            O => \N__10803\,
            I => \N__10794\
        );

    \I__2601\ : Span4Mux_v
    port map (
            O => \N__10800\,
            I => \N__10794\
        );

    \I__2600\ : InMux
    port map (
            O => \N__10799\,
            I => \N__10791\
        );

    \I__2599\ : Span4Mux_v
    port map (
            O => \N__10794\,
            I => \N__10788\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__10791\,
            I => \N__10785\
        );

    \I__2597\ : Sp12to4
    port map (
            O => \N__10788\,
            I => \N__10780\
        );

    \I__2596\ : Span12Mux_v
    port map (
            O => \N__10785\,
            I => \N__10780\
        );

    \I__2595\ : Span12Mux_h
    port map (
            O => \N__10780\,
            I => \N__10777\
        );

    \I__2594\ : Odrv12
    port map (
            O => \N__10777\,
            I => \DRA_c_6\
        );

    \I__2593\ : InMux
    port map (
            O => \N__10774\,
            I => \N__10771\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__10771\,
            I => \N__10768\
        );

    \I__2591\ : Span4Mux_h
    port map (
            O => \N__10768\,
            I => \N__10765\
        );

    \I__2590\ : Odrv4
    port map (
            O => \N__10765\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2589\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10756\
        );

    \I__2588\ : InMux
    port map (
            O => \N__10761\,
            I => \N__10756\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__10756\,
            I => \N__10753\
        );

    \I__2586\ : Odrv12
    port map (
            O => \N__10753\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__10750\,
            I => \N__10747\
        );

    \I__2584\ : InMux
    port map (
            O => \N__10747\,
            I => \N__10744\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__10744\,
            I => \N__10741\
        );

    \I__2582\ : Odrv12
    port map (
            O => \N__10741\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2581\ : InMux
    port map (
            O => \N__10738\,
            I => \N__10734\
        );

    \I__2580\ : InMux
    port map (
            O => \N__10737\,
            I => \N__10730\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__10734\,
            I => \N__10727\
        );

    \I__2578\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10724\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__10730\,
            I => \N__10716\
        );

    \I__2576\ : Span4Mux_h
    port map (
            O => \N__10727\,
            I => \N__10716\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__10724\,
            I => \N__10716\
        );

    \I__2574\ : InMux
    port map (
            O => \N__10723\,
            I => \N__10713\
        );

    \I__2573\ : Span4Mux_v
    port map (
            O => \N__10716\,
            I => \N__10710\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__10713\,
            I => \N__10707\
        );

    \I__2571\ : Span4Mux_v
    port map (
            O => \N__10710\,
            I => \N__10704\
        );

    \I__2570\ : Span12Mux_v
    port map (
            O => \N__10707\,
            I => \N__10699\
        );

    \I__2569\ : Sp12to4
    port map (
            O => \N__10704\,
            I => \N__10699\
        );

    \I__2568\ : Span12Mux_h
    port map (
            O => \N__10699\,
            I => \N__10696\
        );

    \I__2567\ : Odrv12
    port map (
            O => \N__10696\,
            I => \DRA_c_3\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__10693\,
            I => \N__10690\
        );

    \I__2565\ : InMux
    port map (
            O => \N__10690\,
            I => \N__10687\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__10687\,
            I => \N__10684\
        );

    \I__2563\ : Odrv4
    port map (
            O => \N__10684\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2562\ : InMux
    port map (
            O => \N__10681\,
            I => \N__10678\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__10678\,
            I => \N__10672\
        );

    \I__2560\ : InMux
    port map (
            O => \N__10677\,
            I => \N__10669\
        );

    \I__2559\ : InMux
    port map (
            O => \N__10676\,
            I => \N__10666\
        );

    \I__2558\ : InMux
    port map (
            O => \N__10675\,
            I => \N__10663\
        );

    \I__2557\ : Span4Mux_h
    port map (
            O => \N__10672\,
            I => \N__10658\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__10669\,
            I => \N__10658\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__10666\,
            I => \N__10653\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__10663\,
            I => \N__10653\
        );

    \I__2553\ : Span4Mux_v
    port map (
            O => \N__10658\,
            I => \N__10650\
        );

    \I__2552\ : Span4Mux_h
    port map (
            O => \N__10653\,
            I => \N__10647\
        );

    \I__2551\ : Span4Mux_v
    port map (
            O => \N__10650\,
            I => \N__10644\
        );

    \I__2550\ : Sp12to4
    port map (
            O => \N__10647\,
            I => \N__10641\
        );

    \I__2549\ : Sp12to4
    port map (
            O => \N__10644\,
            I => \N__10638\
        );

    \I__2548\ : Span12Mux_v
    port map (
            O => \N__10641\,
            I => \N__10635\
        );

    \I__2547\ : Span12Mux_h
    port map (
            O => \N__10638\,
            I => \N__10632\
        );

    \I__2546\ : Odrv12
    port map (
            O => \N__10635\,
            I => \DRA_c_2\
        );

    \I__2545\ : Odrv12
    port map (
            O => \N__10632\,
            I => \DRA_c_2\
        );

    \I__2544\ : InMux
    port map (
            O => \N__10627\,
            I => \N__10622\
        );

    \I__2543\ : InMux
    port map (
            O => \N__10626\,
            I => \N__10619\
        );

    \I__2542\ : InMux
    port map (
            O => \N__10625\,
            I => \N__10616\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__10622\,
            I => \N__10613\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__10619\,
            I => \N__10607\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__10616\,
            I => \N__10607\
        );

    \I__2538\ : Span4Mux_v
    port map (
            O => \N__10613\,
            I => \N__10604\
        );

    \I__2537\ : InMux
    port map (
            O => \N__10612\,
            I => \N__10601\
        );

    \I__2536\ : Span4Mux_h
    port map (
            O => \N__10607\,
            I => \N__10598\
        );

    \I__2535\ : Sp12to4
    port map (
            O => \N__10604\,
            I => \N__10593\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__10601\,
            I => \N__10593\
        );

    \I__2533\ : Sp12to4
    port map (
            O => \N__10598\,
            I => \N__10590\
        );

    \I__2532\ : Span12Mux_h
    port map (
            O => \N__10593\,
            I => \N__10587\
        );

    \I__2531\ : Span12Mux_v
    port map (
            O => \N__10590\,
            I => \N__10584\
        );

    \I__2530\ : Span12Mux_v
    port map (
            O => \N__10587\,
            I => \N__10581\
        );

    \I__2529\ : Odrv12
    port map (
            O => \N__10584\,
            I => \DRA_c_1\
        );

    \I__2528\ : Odrv12
    port map (
            O => \N__10581\,
            I => \DRA_c_1\
        );

    \I__2527\ : InMux
    port map (
            O => \N__10576\,
            I => \N__10573\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__10573\,
            I => \N__10570\
        );

    \I__2525\ : Odrv12
    port map (
            O => \N__10570\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__10567\,
            I => \N__10564\
        );

    \I__2523\ : InMux
    port map (
            O => \N__10564\,
            I => \N__10557\
        );

    \I__2522\ : InMux
    port map (
            O => \N__10563\,
            I => \N__10557\
        );

    \I__2521\ : InMux
    port map (
            O => \N__10562\,
            I => \N__10554\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__10557\,
            I => \N__10548\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__10554\,
            I => \N__10548\
        );

    \I__2518\ : InMux
    port map (
            O => \N__10553\,
            I => \N__10545\
        );

    \I__2517\ : Span4Mux_v
    port map (
            O => \N__10548\,
            I => \N__10542\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__10545\,
            I => \N__10539\
        );

    \I__2515\ : Sp12to4
    port map (
            O => \N__10542\,
            I => \N__10534\
        );

    \I__2514\ : Span12Mux_v
    port map (
            O => \N__10539\,
            I => \N__10534\
        );

    \I__2513\ : Span12Mux_h
    port map (
            O => \N__10534\,
            I => \N__10531\
        );

    \I__2512\ : Odrv12
    port map (
            O => \N__10531\,
            I => \DRA_c_7\
        );

    \I__2511\ : InMux
    port map (
            O => \N__10528\,
            I => \N__10524\
        );

    \I__2510\ : InMux
    port map (
            O => \N__10527\,
            I => \N__10521\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__10524\,
            I => \N__10516\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10521\,
            I => \N__10516\
        );

    \I__2507\ : Span4Mux_v
    port map (
            O => \N__10516\,
            I => \N__10511\
        );

    \I__2506\ : InMux
    port map (
            O => \N__10515\,
            I => \N__10508\
        );

    \I__2505\ : InMux
    port map (
            O => \N__10514\,
            I => \N__10505\
        );

    \I__2504\ : Sp12to4
    port map (
            O => \N__10511\,
            I => \N__10498\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10508\,
            I => \N__10498\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__10505\,
            I => \N__10498\
        );

    \I__2501\ : Span12Mux_h
    port map (
            O => \N__10498\,
            I => \N__10495\
        );

    \I__2500\ : Odrv12
    port map (
            O => \N__10495\,
            I => \DRA_c_8\
        );

    \I__2499\ : InMux
    port map (
            O => \N__10492\,
            I => \N__10489\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__10489\,
            I => \N__10486\
        );

    \I__2497\ : Odrv4
    port map (
            O => \N__10486\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2496\ : InMux
    port map (
            O => \N__10483\,
            I => \N__10480\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__10480\,
            I => \N__10475\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10479\,
            I => \N__10462\
        );

    \I__2493\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10459\
        );

    \I__2492\ : Span4Mux_v
    port map (
            O => \N__10475\,
            I => \N__10454\
        );

    \I__2491\ : InMux
    port map (
            O => \N__10474\,
            I => \N__10451\
        );

    \I__2490\ : InMux
    port map (
            O => \N__10473\,
            I => \N__10446\
        );

    \I__2489\ : InMux
    port map (
            O => \N__10472\,
            I => \N__10446\
        );

    \I__2488\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10443\
        );

    \I__2487\ : InMux
    port map (
            O => \N__10470\,
            I => \N__10440\
        );

    \I__2486\ : InMux
    port map (
            O => \N__10469\,
            I => \N__10435\
        );

    \I__2485\ : InMux
    port map (
            O => \N__10468\,
            I => \N__10435\
        );

    \I__2484\ : InMux
    port map (
            O => \N__10467\,
            I => \N__10430\
        );

    \I__2483\ : InMux
    port map (
            O => \N__10466\,
            I => \N__10430\
        );

    \I__2482\ : InMux
    port map (
            O => \N__10465\,
            I => \N__10427\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__10462\,
            I => \N__10422\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__10459\,
            I => \N__10422\
        );

    \I__2479\ : InMux
    port map (
            O => \N__10458\,
            I => \N__10419\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10457\,
            I => \N__10411\
        );

    \I__2477\ : Span4Mux_h
    port map (
            O => \N__10454\,
            I => \N__10407\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__10451\,
            I => \N__10404\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__10446\,
            I => \N__10391\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__10443\,
            I => \N__10391\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__10440\,
            I => \N__10391\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__10435\,
            I => \N__10391\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__10430\,
            I => \N__10391\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__10427\,
            I => \N__10391\
        );

    \I__2469\ : Span4Mux_h
    port map (
            O => \N__10422\,
            I => \N__10386\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__10419\,
            I => \N__10386\
        );

    \I__2467\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10383\
        );

    \I__2466\ : InMux
    port map (
            O => \N__10417\,
            I => \N__10380\
        );

    \I__2465\ : InMux
    port map (
            O => \N__10416\,
            I => \N__10373\
        );

    \I__2464\ : InMux
    port map (
            O => \N__10415\,
            I => \N__10373\
        );

    \I__2463\ : InMux
    port map (
            O => \N__10414\,
            I => \N__10373\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__10411\,
            I => \N__10370\
        );

    \I__2461\ : InMux
    port map (
            O => \N__10410\,
            I => \N__10367\
        );

    \I__2460\ : Span4Mux_h
    port map (
            O => \N__10407\,
            I => \N__10362\
        );

    \I__2459\ : Span4Mux_v
    port map (
            O => \N__10404\,
            I => \N__10362\
        );

    \I__2458\ : Span4Mux_v
    port map (
            O => \N__10391\,
            I => \N__10357\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__10386\,
            I => \N__10357\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__10383\,
            I => \N__10352\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__10380\,
            I => \N__10352\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__10373\,
            I => \N__10345\
        );

    \I__2453\ : Sp12to4
    port map (
            O => \N__10370\,
            I => \N__10345\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__10367\,
            I => \N__10345\
        );

    \I__2451\ : Sp12to4
    port map (
            O => \N__10362\,
            I => \N__10340\
        );

    \I__2450\ : Sp12to4
    port map (
            O => \N__10357\,
            I => \N__10340\
        );

    \I__2449\ : Span12Mux_h
    port map (
            O => \N__10352\,
            I => \N__10337\
        );

    \I__2448\ : Span12Mux_v
    port map (
            O => \N__10345\,
            I => \N__10334\
        );

    \I__2447\ : Span12Mux_h
    port map (
            O => \N__10340\,
            I => \N__10331\
        );

    \I__2446\ : Span12Mux_v
    port map (
            O => \N__10337\,
            I => \N__10326\
        );

    \I__2445\ : Span12Mux_h
    port map (
            O => \N__10334\,
            I => \N__10326\
        );

    \I__2444\ : Span12Mux_v
    port map (
            O => \N__10331\,
            I => \N__10323\
        );

    \I__2443\ : Odrv12
    port map (
            O => \N__10326\,
            I => \AGNUS_REV_c\
        );

    \I__2442\ : Odrv12
    port map (
            O => \N__10323\,
            I => \AGNUS_REV_c\
        );

    \I__2441\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10315\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__10315\,
            I => \N__10312\
        );

    \I__2439\ : Odrv12
    port map (
            O => \N__10312\,
            I => \RAS0n_c\
        );

    \I__2438\ : CascadeMux
    port map (
            O => \N__10309\,
            I => \N__10305\
        );

    \I__2437\ : InMux
    port map (
            O => \N__10308\,
            I => \N__10302\
        );

    \I__2436\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10298\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__10302\,
            I => \N__10295\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10301\,
            I => \N__10292\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__10298\,
            I => \N__10289\
        );

    \I__2432\ : Span4Mux_h
    port map (
            O => \N__10295\,
            I => \N__10284\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__10292\,
            I => \N__10284\
        );

    \I__2430\ : Span4Mux_v
    port map (
            O => \N__10289\,
            I => \N__10280\
        );

    \I__2429\ : Span4Mux_v
    port map (
            O => \N__10284\,
            I => \N__10277\
        );

    \I__2428\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10274\
        );

    \I__2427\ : Sp12to4
    port map (
            O => \N__10280\,
            I => \N__10269\
        );

    \I__2426\ : Sp12to4
    port map (
            O => \N__10277\,
            I => \N__10269\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__10274\,
            I => \N__10266\
        );

    \I__2424\ : Span12Mux_h
    port map (
            O => \N__10269\,
            I => \N__10263\
        );

    \I__2423\ : Span12Mux_v
    port map (
            O => \N__10266\,
            I => \N__10260\
        );

    \I__2422\ : Span12Mux_v
    port map (
            O => \N__10263\,
            I => \N__10257\
        );

    \I__2421\ : Span12Mux_v
    port map (
            O => \N__10260\,
            I => \N__10254\
        );

    \I__2420\ : Odrv12
    port map (
            O => \N__10257\,
            I => \DRA_c_9\
        );

    \I__2419\ : Odrv12
    port map (
            O => \N__10254\,
            I => \DRA_c_9\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10249\,
            I => \N__10246\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__10246\,
            I => \N__10243\
        );

    \I__2416\ : Odrv12
    port map (
            O => \N__10243\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2415\ : ClkMux
    port map (
            O => \N__10240\,
            I => \N__10225\
        );

    \I__2414\ : ClkMux
    port map (
            O => \N__10239\,
            I => \N__10225\
        );

    \I__2413\ : ClkMux
    port map (
            O => \N__10238\,
            I => \N__10225\
        );

    \I__2412\ : ClkMux
    port map (
            O => \N__10237\,
            I => \N__10225\
        );

    \I__2411\ : ClkMux
    port map (
            O => \N__10236\,
            I => \N__10225\
        );

    \I__2410\ : GlobalMux
    port map (
            O => \N__10225\,
            I => \N__10222\
        );

    \I__2409\ : gio2CtrlBuf
    port map (
            O => \N__10222\,
            I => \C3_c_g\
        );

    \I__2408\ : CEMux
    port map (
            O => \N__10219\,
            I => \N__10186\
        );

    \I__2407\ : CEMux
    port map (
            O => \N__10218\,
            I => \N__10186\
        );

    \I__2406\ : CEMux
    port map (
            O => \N__10217\,
            I => \N__10186\
        );

    \I__2405\ : CEMux
    port map (
            O => \N__10216\,
            I => \N__10186\
        );

    \I__2404\ : CEMux
    port map (
            O => \N__10215\,
            I => \N__10186\
        );

    \I__2403\ : CEMux
    port map (
            O => \N__10214\,
            I => \N__10186\
        );

    \I__2402\ : CEMux
    port map (
            O => \N__10213\,
            I => \N__10186\
        );

    \I__2401\ : CEMux
    port map (
            O => \N__10212\,
            I => \N__10186\
        );

    \I__2400\ : CEMux
    port map (
            O => \N__10211\,
            I => \N__10186\
        );

    \I__2399\ : CEMux
    port map (
            O => \N__10210\,
            I => \N__10186\
        );

    \I__2398\ : CEMux
    port map (
            O => \N__10209\,
            I => \N__10186\
        );

    \I__2397\ : GlobalMux
    port map (
            O => \N__10186\,
            I => \N__10183\
        );

    \I__2396\ : gio2CtrlBuf
    port map (
            O => \N__10183\,
            I => \DBRn_c_i_0_g\
        );

    \I__2395\ : InMux
    port map (
            O => \N__10180\,
            I => \N__10172\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10179\,
            I => \N__10169\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10178\,
            I => \N__10166\
        );

    \I__2392\ : InMux
    port map (
            O => \N__10177\,
            I => \N__10163\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10176\,
            I => \N__10160\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10175\,
            I => \N__10157\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__10172\,
            I => \N__10153\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__10169\,
            I => \N__10147\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__10166\,
            I => \N__10144\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__10163\,
            I => \N__10130\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__10160\,
            I => \N__10116\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10157\,
            I => \N__10105\
        );

    \I__2383\ : SRMux
    port map (
            O => \N__10156\,
            I => \N__10015\
        );

    \I__2382\ : Glb2LocalMux
    port map (
            O => \N__10153\,
            I => \N__10015\
        );

    \I__2381\ : SRMux
    port map (
            O => \N__10152\,
            I => \N__10015\
        );

    \I__2380\ : SRMux
    port map (
            O => \N__10151\,
            I => \N__10015\
        );

    \I__2379\ : SRMux
    port map (
            O => \N__10150\,
            I => \N__10015\
        );

    \I__2378\ : Glb2LocalMux
    port map (
            O => \N__10147\,
            I => \N__10015\
        );

    \I__2377\ : Glb2LocalMux
    port map (
            O => \N__10144\,
            I => \N__10015\
        );

    \I__2376\ : SRMux
    port map (
            O => \N__10143\,
            I => \N__10015\
        );

    \I__2375\ : SRMux
    port map (
            O => \N__10142\,
            I => \N__10015\
        );

    \I__2374\ : SRMux
    port map (
            O => \N__10141\,
            I => \N__10015\
        );

    \I__2373\ : SRMux
    port map (
            O => \N__10140\,
            I => \N__10015\
        );

    \I__2372\ : SRMux
    port map (
            O => \N__10139\,
            I => \N__10015\
        );

    \I__2371\ : SRMux
    port map (
            O => \N__10138\,
            I => \N__10015\
        );

    \I__2370\ : SRMux
    port map (
            O => \N__10137\,
            I => \N__10015\
        );

    \I__2369\ : SRMux
    port map (
            O => \N__10136\,
            I => \N__10015\
        );

    \I__2368\ : SRMux
    port map (
            O => \N__10135\,
            I => \N__10015\
        );

    \I__2367\ : SRMux
    port map (
            O => \N__10134\,
            I => \N__10015\
        );

    \I__2366\ : SRMux
    port map (
            O => \N__10133\,
            I => \N__10015\
        );

    \I__2365\ : Glb2LocalMux
    port map (
            O => \N__10130\,
            I => \N__10015\
        );

    \I__2364\ : SRMux
    port map (
            O => \N__10129\,
            I => \N__10015\
        );

    \I__2363\ : SRMux
    port map (
            O => \N__10128\,
            I => \N__10015\
        );

    \I__2362\ : SRMux
    port map (
            O => \N__10127\,
            I => \N__10015\
        );

    \I__2361\ : SRMux
    port map (
            O => \N__10126\,
            I => \N__10015\
        );

    \I__2360\ : SRMux
    port map (
            O => \N__10125\,
            I => \N__10015\
        );

    \I__2359\ : SRMux
    port map (
            O => \N__10124\,
            I => \N__10015\
        );

    \I__2358\ : SRMux
    port map (
            O => \N__10123\,
            I => \N__10015\
        );

    \I__2357\ : SRMux
    port map (
            O => \N__10122\,
            I => \N__10015\
        );

    \I__2356\ : SRMux
    port map (
            O => \N__10121\,
            I => \N__10015\
        );

    \I__2355\ : SRMux
    port map (
            O => \N__10120\,
            I => \N__10015\
        );

    \I__2354\ : SRMux
    port map (
            O => \N__10119\,
            I => \N__10015\
        );

    \I__2353\ : Glb2LocalMux
    port map (
            O => \N__10116\,
            I => \N__10015\
        );

    \I__2352\ : SRMux
    port map (
            O => \N__10115\,
            I => \N__10015\
        );

    \I__2351\ : SRMux
    port map (
            O => \N__10114\,
            I => \N__10015\
        );

    \I__2350\ : SRMux
    port map (
            O => \N__10113\,
            I => \N__10015\
        );

    \I__2349\ : SRMux
    port map (
            O => \N__10112\,
            I => \N__10015\
        );

    \I__2348\ : SRMux
    port map (
            O => \N__10111\,
            I => \N__10015\
        );

    \I__2347\ : SRMux
    port map (
            O => \N__10110\,
            I => \N__10015\
        );

    \I__2346\ : SRMux
    port map (
            O => \N__10109\,
            I => \N__10015\
        );

    \I__2345\ : SRMux
    port map (
            O => \N__10108\,
            I => \N__10015\
        );

    \I__2344\ : Glb2LocalMux
    port map (
            O => \N__10105\,
            I => \N__10015\
        );

    \I__2343\ : SRMux
    port map (
            O => \N__10104\,
            I => \N__10015\
        );

    \I__2342\ : SRMux
    port map (
            O => \N__10103\,
            I => \N__10015\
        );

    \I__2341\ : SRMux
    port map (
            O => \N__10102\,
            I => \N__10015\
        );

    \I__2340\ : GlobalMux
    port map (
            O => \N__10015\,
            I => \N__10012\
        );

    \I__2339\ : gio2CtrlBuf
    port map (
            O => \N__10012\,
            I => \RESETn_c_i_g\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10009\,
            I => \N__10005\
        );

    \I__2337\ : InMux
    port map (
            O => \N__10008\,
            I => \N__10002\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__10005\,
            I => \N__9999\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__10002\,
            I => \N__9995\
        );

    \I__2334\ : Span4Mux_v
    port map (
            O => \N__9999\,
            I => \N__9992\
        );

    \I__2333\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9989\
        );

    \I__2332\ : Span12Mux_s9_v
    port map (
            O => \N__9995\,
            I => \N__9986\
        );

    \I__2331\ : Span4Mux_v
    port map (
            O => \N__9992\,
            I => \N__9983\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__9989\,
            I => \N__9980\
        );

    \I__2329\ : Span12Mux_h
    port map (
            O => \N__9986\,
            I => \N__9977\
        );

    \I__2328\ : Span4Mux_v
    port map (
            O => \N__9983\,
            I => \N__9974\
        );

    \I__2327\ : Span4Mux_v
    port map (
            O => \N__9980\,
            I => \N__9971\
        );

    \I__2326\ : Odrv12
    port map (
            O => \N__9977\,
            I => \REG_CYCLEm\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__9974\,
            I => \REG_CYCLEm\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__9971\,
            I => \REG_CYCLEm\
        );

    \I__2323\ : IoInMux
    port map (
            O => \N__9964\,
            I => \N__9961\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__9961\,
            I => \N__9958\
        );

    \I__2321\ : Span4Mux_s3_v
    port map (
            O => \N__9958\,
            I => \N__9955\
        );

    \I__2320\ : Span4Mux_v
    port map (
            O => \N__9955\,
            I => \N__9952\
        );

    \I__2319\ : Odrv4
    port map (
            O => \N__9952\,
            I => \DRDENn_c\
        );

    \I__2318\ : InMux
    port map (
            O => \N__9949\,
            I => \N__9946\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__9946\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__9943\,
            I => \N__9940\
        );

    \I__2315\ : InMux
    port map (
            O => \N__9940\,
            I => \N__9937\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__9937\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2313\ : InMux
    port map (
            O => \N__9934\,
            I => \N__9931\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__9931\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2311\ : InMux
    port map (
            O => \N__9928\,
            I => \N__9925\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__9925\,
            I => \N__9919\
        );

    \I__2309\ : InMux
    port map (
            O => \N__9924\,
            I => \N__9914\
        );

    \I__2308\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9914\
        );

    \I__2307\ : InMux
    port map (
            O => \N__9922\,
            I => \N__9911\
        );

    \I__2306\ : Span4Mux_h
    port map (
            O => \N__9919\,
            I => \N__9904\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__9914\,
            I => \N__9904\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__9911\,
            I => \N__9904\
        );

    \I__2303\ : Span4Mux_v
    port map (
            O => \N__9904\,
            I => \N__9901\
        );

    \I__2302\ : Span4Mux_v
    port map (
            O => \N__9901\,
            I => \N__9898\
        );

    \I__2301\ : Sp12to4
    port map (
            O => \N__9898\,
            I => \N__9895\
        );

    \I__2300\ : Span12Mux_h
    port map (
            O => \N__9895\,
            I => \N__9892\
        );

    \I__2299\ : Odrv12
    port map (
            O => \N__9892\,
            I => \DRA_c_4\
        );

    \I__2298\ : InMux
    port map (
            O => \N__9889\,
            I => \N__9881\
        );

    \I__2297\ : InMux
    port map (
            O => \N__9888\,
            I => \N__9881\
        );

    \I__2296\ : InMux
    port map (
            O => \N__9887\,
            I => \N__9878\
        );

    \I__2295\ : InMux
    port map (
            O => \N__9886\,
            I => \N__9875\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__9881\,
            I => \N__9868\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__9878\,
            I => \N__9868\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__9875\,
            I => \N__9868\
        );

    \I__2291\ : Span12Mux_v
    port map (
            O => \N__9868\,
            I => \N__9865\
        );

    \I__2290\ : Span12Mux_h
    port map (
            O => \N__9865\,
            I => \N__9862\
        );

    \I__2289\ : Odrv12
    port map (
            O => \N__9862\,
            I => \DRA_c_5\
        );

    \I__2288\ : InMux
    port map (
            O => \N__9859\,
            I => \N__9856\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__9856\,
            I => \N__9853\
        );

    \I__2286\ : Span4Mux_v
    port map (
            O => \N__9853\,
            I => \N__9850\
        );

    \I__2285\ : Odrv4
    port map (
            O => \N__9850\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2284\ : InMux
    port map (
            O => \N__9847\,
            I => \N__9844\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__9844\,
            I => \N__9841\
        );

    \I__2282\ : Span4Mux_h
    port map (
            O => \N__9841\,
            I => \N__9838\
        );

    \I__2281\ : Odrv4
    port map (
            O => \N__9838\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2280\ : InMux
    port map (
            O => \N__9835\,
            I => \N__9832\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__9832\,
            I => \N__9829\
        );

    \I__2278\ : Odrv4
    port map (
            O => \N__9829\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2277\ : InMux
    port map (
            O => \N__9826\,
            I => \N__9822\
        );

    \I__2276\ : InMux
    port map (
            O => \N__9825\,
            I => \N__9819\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__9822\,
            I => \N__9816\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__9819\,
            I => \N__9813\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__9816\,
            I => \N__9808\
        );

    \I__2272\ : Span4Mux_v
    port map (
            O => \N__9813\,
            I => \N__9808\
        );

    \I__2271\ : Sp12to4
    port map (
            O => \N__9808\,
            I => \N__9805\
        );

    \I__2270\ : Span12Mux_v
    port map (
            O => \N__9805\,
            I => \N__9802\
        );

    \I__2269\ : Span12Mux_h
    port map (
            O => \N__9802\,
            I => \N__9799\
        );

    \I__2268\ : Odrv12
    port map (
            O => \N__9799\,
            I => \DRA_c_0\
        );

    \I__2267\ : InMux
    port map (
            O => \N__9796\,
            I => \N__9793\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__9793\,
            I => \N__9790\
        );

    \I__2265\ : Span4Mux_h
    port map (
            O => \N__9790\,
            I => \N__9787\
        );

    \I__2264\ : Span4Mux_h
    port map (
            O => \N__9787\,
            I => \N__9784\
        );

    \I__2263\ : Odrv4
    port map (
            O => \N__9784\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2262\ : InMux
    port map (
            O => \N__9781\,
            I => \N__9778\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__9778\,
            I => \N__9775\
        );

    \I__2260\ : Span4Mux_v
    port map (
            O => \N__9775\,
            I => \N__9772\
        );

    \I__2259\ : Odrv4
    port map (
            O => \N__9772\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2258\ : InMux
    port map (
            O => \N__9769\,
            I => \N__9766\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__9766\,
            I => \N__9763\
        );

    \I__2256\ : Span4Mux_v
    port map (
            O => \N__9763\,
            I => \N__9760\
        );

    \I__2255\ : Sp12to4
    port map (
            O => \N__9760\,
            I => \N__9757\
        );

    \I__2254\ : Span12Mux_h
    port map (
            O => \N__9757\,
            I => \N__9754\
        );

    \I__2253\ : Odrv12
    port map (
            O => \N__9754\,
            I => \A_c_6\
        );

    \I__2252\ : InMux
    port map (
            O => \N__9751\,
            I => \N__9748\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__9748\,
            I => \N__9745\
        );

    \I__2250\ : Span4Mux_v
    port map (
            O => \N__9745\,
            I => \N__9742\
        );

    \I__2249\ : Span4Mux_h
    port map (
            O => \N__9742\,
            I => \N__9739\
        );

    \I__2248\ : Sp12to4
    port map (
            O => \N__9739\,
            I => \N__9736\
        );

    \I__2247\ : Odrv12
    port map (
            O => \N__9736\,
            I => \A_c_13\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__9733\,
            I => \N__9728\
        );

    \I__2245\ : InMux
    port map (
            O => \N__9732\,
            I => \N__9711\
        );

    \I__2244\ : InMux
    port map (
            O => \N__9731\,
            I => \N__9711\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9711\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9727\,
            I => \N__9711\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9726\,
            I => \N__9704\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9725\,
            I => \N__9698\
        );

    \I__2239\ : InMux
    port map (
            O => \N__9724\,
            I => \N__9698\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9723\,
            I => \N__9693\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9722\,
            I => \N__9693\
        );

    \I__2236\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9690\
        );

    \I__2235\ : InMux
    port map (
            O => \N__9720\,
            I => \N__9687\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__9711\,
            I => \N__9684\
        );

    \I__2233\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9681\
        );

    \I__2232\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9678\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__9708\,
            I => \N__9674\
        );

    \I__2230\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9669\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__9704\,
            I => \N__9666\
        );

    \I__2228\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9659\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__9698\,
            I => \N__9656\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__9693\,
            I => \N__9653\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__9690\,
            I => \N__9648\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__9687\,
            I => \N__9648\
        );

    \I__2223\ : Span4Mux_h
    port map (
            O => \N__9684\,
            I => \N__9641\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__9681\,
            I => \N__9641\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__9678\,
            I => \N__9641\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9677\,
            I => \N__9638\
        );

    \I__2219\ : InMux
    port map (
            O => \N__9674\,
            I => \N__9635\
        );

    \I__2218\ : InMux
    port map (
            O => \N__9673\,
            I => \N__9632\
        );

    \I__2217\ : InMux
    port map (
            O => \N__9672\,
            I => \N__9629\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__9669\,
            I => \N__9624\
        );

    \I__2215\ : Span4Mux_h
    port map (
            O => \N__9666\,
            I => \N__9624\
        );

    \I__2214\ : InMux
    port map (
            O => \N__9665\,
            I => \N__9615\
        );

    \I__2213\ : InMux
    port map (
            O => \N__9664\,
            I => \N__9615\
        );

    \I__2212\ : InMux
    port map (
            O => \N__9663\,
            I => \N__9615\
        );

    \I__2211\ : InMux
    port map (
            O => \N__9662\,
            I => \N__9615\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9659\,
            I => \N__9604\
        );

    \I__2209\ : Span4Mux_v
    port map (
            O => \N__9656\,
            I => \N__9604\
        );

    \I__2208\ : Span4Mux_v
    port map (
            O => \N__9653\,
            I => \N__9604\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__9648\,
            I => \N__9604\
        );

    \I__2206\ : Span4Mux_v
    port map (
            O => \N__9641\,
            I => \N__9604\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__9638\,
            I => \CPU_CYCLEm\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__9635\,
            I => \CPU_CYCLEm\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__9632\,
            I => \CPU_CYCLEm\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__9629\,
            I => \CPU_CYCLEm\
        );

    \I__2201\ : Odrv4
    port map (
            O => \N__9624\,
            I => \CPU_CYCLEm\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__9615\,
            I => \CPU_CYCLEm\
        );

    \I__2199\ : Odrv4
    port map (
            O => \N__9604\,
            I => \CPU_CYCLEm\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9580\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__9588\,
            I => \N__9577\
        );

    \I__2196\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9566\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9586\,
            I => \N__9566\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9585\,
            I => \N__9563\
        );

    \I__2193\ : InMux
    port map (
            O => \N__9584\,
            I => \N__9558\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9583\,
            I => \N__9558\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__9580\,
            I => \N__9548\
        );

    \I__2190\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9543\
        );

    \I__2189\ : InMux
    port map (
            O => \N__9576\,
            I => \N__9543\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9540\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9574\,
            I => \N__9537\
        );

    \I__2186\ : InMux
    port map (
            O => \N__9573\,
            I => \N__9532\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9572\,
            I => \N__9532\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9529\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__9566\,
            I => \N__9522\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__9563\,
            I => \N__9517\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9558\,
            I => \N__9517\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9557\,
            I => \N__9508\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9556\,
            I => \N__9508\
        );

    \I__2178\ : InMux
    port map (
            O => \N__9555\,
            I => \N__9508\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9554\,
            I => \N__9508\
        );

    \I__2176\ : InMux
    port map (
            O => \N__9553\,
            I => \N__9501\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9552\,
            I => \N__9501\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9551\,
            I => \N__9501\
        );

    \I__2173\ : Span4Mux_v
    port map (
            O => \N__9548\,
            I => \N__9490\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9543\,
            I => \N__9490\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9540\,
            I => \N__9490\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9537\,
            I => \N__9490\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__9532\,
            I => \N__9490\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__9529\,
            I => \N__9487\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9484\
        );

    \I__2166\ : CascadeMux
    port map (
            O => \N__9527\,
            I => \N__9481\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__9526\,
            I => \N__9478\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9525\,
            I => \N__9475\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__9522\,
            I => \N__9464\
        );

    \I__2162\ : Span4Mux_v
    port map (
            O => \N__9517\,
            I => \N__9464\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__9508\,
            I => \N__9464\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__9501\,
            I => \N__9464\
        );

    \I__2159\ : Span4Mux_v
    port map (
            O => \N__9490\,
            I => \N__9464\
        );

    \I__2158\ : Span4Mux_h
    port map (
            O => \N__9487\,
            I => \N__9459\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9484\,
            I => \N__9459\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9454\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9478\,
            I => \N__9454\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9475\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__9464\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2152\ : Odrv4
    port map (
            O => \N__9459\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__9454\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__9445\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9442\,
            I => \N__9439\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9439\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9436\,
            I => \N__9433\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__9433\,
            I => \N__9429\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9432\,
            I => \N__9426\
        );

    \I__2144\ : Span4Mux_h
    port map (
            O => \N__9429\,
            I => \N__9423\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9426\,
            I => \N__9420\
        );

    \I__2142\ : Span4Mux_h
    port map (
            O => \N__9423\,
            I => \N__9415\
        );

    \I__2141\ : Span4Mux_v
    port map (
            O => \N__9420\,
            I => \N__9415\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__9415\,
            I => \DBRn_c_i\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9409\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9409\,
            I => \N__9406\
        );

    \I__2137\ : Span4Mux_h
    port map (
            O => \N__9406\,
            I => \N__9402\
        );

    \I__2136\ : InMux
    port map (
            O => \N__9405\,
            I => \N__9399\
        );

    \I__2135\ : Span4Mux_h
    port map (
            O => \N__9402\,
            I => \N__9396\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9399\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2133\ : Odrv4
    port map (
            O => \N__9396\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__9391\,
            I => \N__9388\
        );

    \I__2131\ : InMux
    port map (
            O => \N__9388\,
            I => \N__9385\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__9385\,
            I => \N__9381\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__9384\,
            I => \N__9377\
        );

    \I__2128\ : Span4Mux_h
    port map (
            O => \N__9381\,
            I => \N__9373\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9380\,
            I => \N__9368\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9377\,
            I => \N__9368\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9376\,
            I => \N__9365\
        );

    \I__2124\ : Span4Mux_h
    port map (
            O => \N__9373\,
            I => \N__9362\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__9368\,
            I => \N__9359\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9365\,
            I => \N__9352\
        );

    \I__2121\ : Sp12to4
    port map (
            O => \N__9362\,
            I => \N__9352\
        );

    \I__2120\ : Span12Mux_h
    port map (
            O => \N__9359\,
            I => \N__9352\
        );

    \I__2119\ : Span12Mux_v
    port map (
            O => \N__9352\,
            I => \N__9349\
        );

    \I__2118\ : Odrv12
    port map (
            O => \N__9349\,
            I => \CLK40_PLL_i\
        );

    \I__2117\ : IoInMux
    port map (
            O => \N__9346\,
            I => \N__9343\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__9343\,
            I => \N__9340\
        );

    \I__2115\ : Span4Mux_s0_v
    port map (
            O => \N__9340\,
            I => \N__9335\
        );

    \I__2114\ : IoInMux
    port map (
            O => \N__9339\,
            I => \N__9332\
        );

    \I__2113\ : IoInMux
    port map (
            O => \N__9338\,
            I => \N__9329\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__9335\,
            I => \N__9326\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__9332\,
            I => \N__9323\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9329\,
            I => \N__9320\
        );

    \I__2109\ : Sp12to4
    port map (
            O => \N__9326\,
            I => \N__9315\
        );

    \I__2108\ : Span12Mux_s4_v
    port map (
            O => \N__9323\,
            I => \N__9315\
        );

    \I__2107\ : Span12Mux_s4_h
    port map (
            O => \N__9320\,
            I => \N__9312\
        );

    \I__2106\ : Span12Mux_h
    port map (
            O => \N__9315\,
            I => \N__9307\
        );

    \I__2105\ : Span12Mux_h
    port map (
            O => \N__9312\,
            I => \N__9307\
        );

    \I__2104\ : Odrv12
    port map (
            O => \N__9307\,
            I => \CLK40_PLL_i_i\
        );

    \I__2103\ : InMux
    port map (
            O => \N__9304\,
            I => \N__9289\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9303\,
            I => \N__9289\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9302\,
            I => \N__9289\
        );

    \I__2100\ : InMux
    port map (
            O => \N__9301\,
            I => \N__9282\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9300\,
            I => \N__9282\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9299\,
            I => \N__9282\
        );

    \I__2097\ : InMux
    port map (
            O => \N__9298\,
            I => \N__9277\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9277\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9272\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__9289\,
            I => \N__9267\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__9282\,
            I => \N__9267\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__9277\,
            I => \N__9263\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9276\,
            I => \N__9260\
        );

    \I__2090\ : InMux
    port map (
            O => \N__9275\,
            I => \N__9256\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__9272\,
            I => \N__9251\
        );

    \I__2088\ : Span4Mux_v
    port map (
            O => \N__9267\,
            I => \N__9248\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9266\,
            I => \N__9245\
        );

    \I__2086\ : Span4Mux_h
    port map (
            O => \N__9263\,
            I => \N__9237\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__9260\,
            I => \N__9237\
        );

    \I__2084\ : InMux
    port map (
            O => \N__9259\,
            I => \N__9234\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__9256\,
            I => \N__9231\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9255\,
            I => \N__9228\
        );

    \I__2081\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9225\
        );

    \I__2080\ : Span4Mux_h
    port map (
            O => \N__9251\,
            I => \N__9222\
        );

    \I__2079\ : Span4Mux_h
    port map (
            O => \N__9248\,
            I => \N__9219\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__9245\,
            I => \N__9216\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9244\,
            I => \N__9213\
        );

    \I__2076\ : InMux
    port map (
            O => \N__9243\,
            I => \N__9208\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9242\,
            I => \N__9208\
        );

    \I__2074\ : Span4Mux_h
    port map (
            O => \N__9237\,
            I => \N__9203\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__9234\,
            I => \N__9203\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__9231\,
            I => \N__9198\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__9228\,
            I => \N__9198\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__9225\,
            I => \N__9195\
        );

    \I__2069\ : Span4Mux_h
    port map (
            O => \N__9222\,
            I => \N__9185\
        );

    \I__2068\ : Span4Mux_v
    port map (
            O => \N__9219\,
            I => \N__9180\
        );

    \I__2067\ : Span4Mux_v
    port map (
            O => \N__9216\,
            I => \N__9180\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__9213\,
            I => \N__9175\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9208\,
            I => \N__9175\
        );

    \I__2064\ : Span4Mux_v
    port map (
            O => \N__9203\,
            I => \N__9168\
        );

    \I__2063\ : Span4Mux_v
    port map (
            O => \N__9198\,
            I => \N__9168\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__9195\,
            I => \N__9168\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9194\,
            I => \N__9161\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9193\,
            I => \N__9161\
        );

    \I__2059\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9161\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9191\,
            I => \N__9158\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9190\,
            I => \N__9153\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9189\,
            I => \N__9153\
        );

    \I__2055\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9150\
        );

    \I__2054\ : Sp12to4
    port map (
            O => \N__9185\,
            I => \N__9147\
        );

    \I__2053\ : Sp12to4
    port map (
            O => \N__9180\,
            I => \N__9132\
        );

    \I__2052\ : Span12Mux_v
    port map (
            O => \N__9175\,
            I => \N__9132\
        );

    \I__2051\ : Sp12to4
    port map (
            O => \N__9168\,
            I => \N__9132\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__9161\,
            I => \N__9132\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9158\,
            I => \N__9132\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9153\,
            I => \N__9132\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9150\,
            I => \N__9132\
        );

    \I__2046\ : Span12Mux_v
    port map (
            O => \N__9147\,
            I => \N__9127\
        );

    \I__2045\ : Span12Mux_h
    port map (
            O => \N__9132\,
            I => \N__9127\
        );

    \I__2044\ : Odrv12
    port map (
            O => \N__9127\,
            I => \RESETn_c\
        );

    \I__2043\ : IoInMux
    port map (
            O => \N__9124\,
            I => \N__9121\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9121\,
            I => \N__9118\
        );

    \I__2041\ : Span12Mux_s9_v
    port map (
            O => \N__9118\,
            I => \N__9115\
        );

    \I__2040\ : Odrv12
    port map (
            O => \N__9115\,
            I => \RESETn_c_i\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9112\,
            I => \N__9109\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__9109\,
            I => \N__9106\
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__9106\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9103\,
            I => \N__9100\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__9100\,
            I => \N__9097\
        );

    \I__2034\ : Odrv4
    port map (
            O => \N__9097\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9091\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9091\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2031\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9082\
        );

    \I__2030\ : InMux
    port map (
            O => \N__9087\,
            I => \N__9082\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__9082\,
            I => \N__9079\
        );

    \I__2028\ : Span4Mux_v
    port map (
            O => \N__9079\,
            I => \N__9076\
        );

    \I__2027\ : Odrv4
    port map (
            O => \N__9076\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__9073\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\
        );

    \I__2025\ : CascadeMux
    port map (
            O => \N__9070\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0_cascade_\
        );

    \I__2024\ : InMux
    port map (
            O => \N__9067\,
            I => \N__9064\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9064\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__2022\ : IoInMux
    port map (
            O => \N__9061\,
            I => \N__9058\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9058\,
            I => \N__9055\
        );

    \I__2020\ : Span4Mux_s3_v
    port map (
            O => \N__9055\,
            I => \N__9052\
        );

    \I__2019\ : Span4Mux_v
    port map (
            O => \N__9052\,
            I => \N__9049\
        );

    \I__2018\ : Span4Mux_v
    port map (
            O => \N__9049\,
            I => \N__9046\
        );

    \I__2017\ : Span4Mux_h
    port map (
            O => \N__9046\,
            I => \N__9043\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__9043\,
            I => \CMA_c_0\
        );

    \I__2015\ : InMux
    port map (
            O => \N__9040\,
            I => \N__9037\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__9037\,
            I => \N__9034\
        );

    \I__2013\ : Span4Mux_v
    port map (
            O => \N__9034\,
            I => \N__9031\
        );

    \I__2012\ : Sp12to4
    port map (
            O => \N__9031\,
            I => \N__9028\
        );

    \I__2011\ : Span12Mux_h
    port map (
            O => \N__9028\,
            I => \N__9025\
        );

    \I__2010\ : Span12Mux_v
    port map (
            O => \N__9025\,
            I => \N__9022\
        );

    \I__2009\ : Odrv12
    port map (
            O => \N__9022\,
            I => \A_c_19\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__9019\,
            I => \N__9014\
        );

    \I__2007\ : InMux
    port map (
            O => \N__9018\,
            I => \N__9011\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__9017\,
            I => \N__9008\
        );

    \I__2005\ : InMux
    port map (
            O => \N__9014\,
            I => \N__9005\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__9011\,
            I => \N__9002\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9008\,
            I => \N__8999\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9005\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__2001\ : Odrv4
    port map (
            O => \N__9002\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__8999\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1999\ : IoInMux
    port map (
            O => \N__8992\,
            I => \N__8989\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__8989\,
            I => \N__8986\
        );

    \I__1997\ : Span4Mux_s3_h
    port map (
            O => \N__8986\,
            I => \N__8983\
        );

    \I__1996\ : Sp12to4
    port map (
            O => \N__8983\,
            I => \N__8980\
        );

    \I__1995\ : Span12Mux_s11_v
    port map (
            O => \N__8980\,
            I => \N__8977\
        );

    \I__1994\ : Span12Mux_h
    port map (
            O => \N__8977\,
            I => \N__8974\
        );

    \I__1993\ : Odrv12
    port map (
            O => \N__8974\,
            I => \CMA_c_9\
        );

    \I__1992\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8968\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__8968\,
            I => \N__8965\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__8965\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1989\ : IoInMux
    port map (
            O => \N__8962\,
            I => \N__8959\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__8959\,
            I => \N__8956\
        );

    \I__1987\ : Span12Mux_s3_h
    port map (
            O => \N__8956\,
            I => \N__8953\
        );

    \I__1986\ : Span12Mux_h
    port map (
            O => \N__8953\,
            I => \N__8950\
        );

    \I__1985\ : Odrv12
    port map (
            O => \N__8950\,
            I => \CMA_c_7\
        );

    \I__1984\ : IoInMux
    port map (
            O => \N__8947\,
            I => \N__8944\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__8944\,
            I => \N__8941\
        );

    \I__1982\ : IoSpan4Mux
    port map (
            O => \N__8941\,
            I => \N__8938\
        );

    \I__1981\ : Sp12to4
    port map (
            O => \N__8938\,
            I => \N__8935\
        );

    \I__1980\ : Span12Mux_s7_v
    port map (
            O => \N__8935\,
            I => \N__8932\
        );

    \I__1979\ : Span12Mux_h
    port map (
            O => \N__8932\,
            I => \N__8929\
        );

    \I__1978\ : Odrv12
    port map (
            O => \N__8929\,
            I => \CMA_c_4\
        );

    \I__1977\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8923\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__8923\,
            I => \N__8920\
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__8920\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1974\ : InMux
    port map (
            O => \N__8917\,
            I => \N__8912\
        );

    \I__1973\ : InMux
    port map (
            O => \N__8916\,
            I => \N__8909\
        );

    \I__1972\ : InMux
    port map (
            O => \N__8915\,
            I => \N__8904\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__8912\,
            I => \N__8899\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__8909\,
            I => \N__8899\
        );

    \I__1969\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8894\
        );

    \I__1968\ : InMux
    port map (
            O => \N__8907\,
            I => \N__8894\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__8904\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__8899\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__8894\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__8887\,
            I => \N__8880\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8886\,
            I => \N__8877\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__8885\,
            I => \N__8874\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__8884\,
            I => \N__8869\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__8883\,
            I => \N__8866\
        );

    \I__1959\ : InMux
    port map (
            O => \N__8880\,
            I => \N__8862\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__8877\,
            I => \N__8859\
        );

    \I__1957\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8856\
        );

    \I__1956\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8853\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8872\,
            I => \N__8850\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8869\,
            I => \N__8847\
        );

    \I__1953\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8844\
        );

    \I__1952\ : InMux
    port map (
            O => \N__8865\,
            I => \N__8841\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__8862\,
            I => \N__8838\
        );

    \I__1950\ : Span4Mux_v
    port map (
            O => \N__8859\,
            I => \N__8833\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__8856\,
            I => \N__8833\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__8853\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__8850\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__8847\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__8844\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__8841\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__8838\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1942\ : Odrv4
    port map (
            O => \N__8833\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__8818\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_\
        );

    \I__1940\ : IoInMux
    port map (
            O => \N__8815\,
            I => \N__8812\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__8812\,
            I => \N__8809\
        );

    \I__1938\ : IoSpan4Mux
    port map (
            O => \N__8809\,
            I => \N__8806\
        );

    \I__1937\ : Span4Mux_s1_h
    port map (
            O => \N__8806\,
            I => \N__8803\
        );

    \I__1936\ : Sp12to4
    port map (
            O => \N__8803\,
            I => \N__8800\
        );

    \I__1935\ : Span12Mux_h
    port map (
            O => \N__8800\,
            I => \N__8797\
        );

    \I__1934\ : Odrv12
    port map (
            O => \N__8797\,
            I => \CMA_c_6\
        );

    \I__1933\ : InMux
    port map (
            O => \N__8794\,
            I => \N__8791\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__8791\,
            I => \N__8769\
        );

    \I__1931\ : ClkMux
    port map (
            O => \N__8790\,
            I => \N__8671\
        );

    \I__1930\ : ClkMux
    port map (
            O => \N__8789\,
            I => \N__8671\
        );

    \I__1929\ : ClkMux
    port map (
            O => \N__8788\,
            I => \N__8671\
        );

    \I__1928\ : ClkMux
    port map (
            O => \N__8787\,
            I => \N__8671\
        );

    \I__1927\ : ClkMux
    port map (
            O => \N__8786\,
            I => \N__8671\
        );

    \I__1926\ : ClkMux
    port map (
            O => \N__8785\,
            I => \N__8671\
        );

    \I__1925\ : ClkMux
    port map (
            O => \N__8784\,
            I => \N__8671\
        );

    \I__1924\ : ClkMux
    port map (
            O => \N__8783\,
            I => \N__8671\
        );

    \I__1923\ : ClkMux
    port map (
            O => \N__8782\,
            I => \N__8671\
        );

    \I__1922\ : ClkMux
    port map (
            O => \N__8781\,
            I => \N__8671\
        );

    \I__1921\ : ClkMux
    port map (
            O => \N__8780\,
            I => \N__8671\
        );

    \I__1920\ : ClkMux
    port map (
            O => \N__8779\,
            I => \N__8671\
        );

    \I__1919\ : ClkMux
    port map (
            O => \N__8778\,
            I => \N__8671\
        );

    \I__1918\ : ClkMux
    port map (
            O => \N__8777\,
            I => \N__8671\
        );

    \I__1917\ : ClkMux
    port map (
            O => \N__8776\,
            I => \N__8671\
        );

    \I__1916\ : ClkMux
    port map (
            O => \N__8775\,
            I => \N__8671\
        );

    \I__1915\ : ClkMux
    port map (
            O => \N__8774\,
            I => \N__8671\
        );

    \I__1914\ : ClkMux
    port map (
            O => \N__8773\,
            I => \N__8671\
        );

    \I__1913\ : ClkMux
    port map (
            O => \N__8772\,
            I => \N__8671\
        );

    \I__1912\ : Glb2LocalMux
    port map (
            O => \N__8769\,
            I => \N__8671\
        );

    \I__1911\ : ClkMux
    port map (
            O => \N__8768\,
            I => \N__8671\
        );

    \I__1910\ : ClkMux
    port map (
            O => \N__8767\,
            I => \N__8671\
        );

    \I__1909\ : ClkMux
    port map (
            O => \N__8766\,
            I => \N__8671\
        );

    \I__1908\ : ClkMux
    port map (
            O => \N__8765\,
            I => \N__8671\
        );

    \I__1907\ : ClkMux
    port map (
            O => \N__8764\,
            I => \N__8671\
        );

    \I__1906\ : ClkMux
    port map (
            O => \N__8763\,
            I => \N__8671\
        );

    \I__1905\ : ClkMux
    port map (
            O => \N__8762\,
            I => \N__8671\
        );

    \I__1904\ : ClkMux
    port map (
            O => \N__8761\,
            I => \N__8671\
        );

    \I__1903\ : ClkMux
    port map (
            O => \N__8760\,
            I => \N__8671\
        );

    \I__1902\ : ClkMux
    port map (
            O => \N__8759\,
            I => \N__8671\
        );

    \I__1901\ : ClkMux
    port map (
            O => \N__8758\,
            I => \N__8671\
        );

    \I__1900\ : ClkMux
    port map (
            O => \N__8757\,
            I => \N__8671\
        );

    \I__1899\ : ClkMux
    port map (
            O => \N__8756\,
            I => \N__8671\
        );

    \I__1898\ : ClkMux
    port map (
            O => \N__8755\,
            I => \N__8671\
        );

    \I__1897\ : ClkMux
    port map (
            O => \N__8754\,
            I => \N__8671\
        );

    \I__1896\ : ClkMux
    port map (
            O => \N__8753\,
            I => \N__8671\
        );

    \I__1895\ : ClkMux
    port map (
            O => \N__8752\,
            I => \N__8671\
        );

    \I__1894\ : ClkMux
    port map (
            O => \N__8751\,
            I => \N__8671\
        );

    \I__1893\ : ClkMux
    port map (
            O => \N__8750\,
            I => \N__8671\
        );

    \I__1892\ : GlobalMux
    port map (
            O => \N__8671\,
            I => \CLK80_PLL\
        );

    \I__1891\ : CEMux
    port map (
            O => \N__8668\,
            I => \N__8664\
        );

    \I__1890\ : CEMux
    port map (
            O => \N__8667\,
            I => \N__8661\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__8664\,
            I => \N__8657\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8661\,
            I => \N__8654\
        );

    \I__1887\ : CEMux
    port map (
            O => \N__8660\,
            I => \N__8651\
        );

    \I__1886\ : Span4Mux_h
    port map (
            O => \N__8657\,
            I => \N__8647\
        );

    \I__1885\ : Span12Mux_h
    port map (
            O => \N__8654\,
            I => \N__8641\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__8651\,
            I => \N__8638\
        );

    \I__1883\ : CEMux
    port map (
            O => \N__8650\,
            I => \N__8635\
        );

    \I__1882\ : Span4Mux_h
    port map (
            O => \N__8647\,
            I => \N__8632\
        );

    \I__1881\ : CEMux
    port map (
            O => \N__8646\,
            I => \N__8629\
        );

    \I__1880\ : CEMux
    port map (
            O => \N__8645\,
            I => \N__8626\
        );

    \I__1879\ : CEMux
    port map (
            O => \N__8644\,
            I => \N__8623\
        );

    \I__1878\ : Odrv12
    port map (
            O => \N__8641\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1877\ : Odrv12
    port map (
            O => \N__8638\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8635\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1875\ : Odrv4
    port map (
            O => \N__8632\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__8629\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__8626\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8623\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1871\ : IoInMux
    port map (
            O => \N__8608\,
            I => \N__8605\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8605\,
            I => \N__8602\
        );

    \I__1869\ : Span12Mux_s8_v
    port map (
            O => \N__8602\,
            I => \N__8599\
        );

    \I__1868\ : Odrv12
    port map (
            O => \N__8599\,
            I => \N_182\
        );

    \I__1867\ : InMux
    port map (
            O => \N__8596\,
            I => \N__8592\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8589\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8592\,
            I => \N__8586\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8589\,
            I => \N__8583\
        );

    \I__1863\ : Span4Mux_v
    port map (
            O => \N__8586\,
            I => \N__8580\
        );

    \I__1862\ : Span4Mux_h
    port map (
            O => \N__8583\,
            I => \N__8577\
        );

    \I__1861\ : Span4Mux_v
    port map (
            O => \N__8580\,
            I => \N__8573\
        );

    \I__1860\ : Sp12to4
    port map (
            O => \N__8577\,
            I => \N__8570\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8567\
        );

    \I__1858\ : Odrv4
    port map (
            O => \N__8573\,
            I => \DS_ENm\
        );

    \I__1857\ : Odrv12
    port map (
            O => \N__8570\,
            I => \DS_ENm\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8567\,
            I => \DS_ENm\
        );

    \I__1855\ : IoInMux
    port map (
            O => \N__8560\,
            I => \N__8557\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8557\,
            I => \N__8554\
        );

    \I__1853\ : Span12Mux_s0_v
    port map (
            O => \N__8554\,
            I => \N__8551\
        );

    \I__1852\ : Span12Mux_h
    port map (
            O => \N__8551\,
            I => \N__8548\
        );

    \I__1851\ : Odrv12
    port map (
            O => \N__8548\,
            I => \N_184\
        );

    \I__1850\ : IoInMux
    port map (
            O => \N__8545\,
            I => \N__8542\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8542\,
            I => \N__8539\
        );

    \I__1848\ : Span4Mux_s2_v
    port map (
            O => \N__8539\,
            I => \N__8536\
        );

    \I__1847\ : Span4Mux_v
    port map (
            O => \N__8536\,
            I => \N__8533\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__8533\,
            I => \N_245_i\
        );

    \I__1845\ : IoInMux
    port map (
            O => \N__8530\,
            I => \N__8527\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__8527\,
            I => \N__8524\
        );

    \I__1843\ : Span12Mux_s6_v
    port map (
            O => \N__8524\,
            I => \N__8521\
        );

    \I__1842\ : Odrv12
    port map (
            O => \N__8521\,
            I => \N_242_i\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8518\,
            I => \N__8509\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8509\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8509\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8509\,
            I => \N__8503\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8508\,
            I => \N__8500\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__8507\,
            I => \N__8497\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8506\,
            I => \N__8492\
        );

    \I__1834\ : Span4Mux_h
    port map (
            O => \N__8503\,
            I => \N__8487\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__8500\,
            I => \N__8487\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8497\,
            I => \N__8484\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8481\
        );

    \I__1830\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8478\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__8492\,
            I => \N__8475\
        );

    \I__1828\ : Span4Mux_h
    port map (
            O => \N__8487\,
            I => \N__8472\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8484\,
            I => \N__8463\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__8481\,
            I => \N__8463\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__8478\,
            I => \N__8463\
        );

    \I__1824\ : Sp12to4
    port map (
            O => \N__8475\,
            I => \N__8463\
        );

    \I__1823\ : Span4Mux_v
    port map (
            O => \N__8472\,
            I => \N__8460\
        );

    \I__1822\ : Span12Mux_v
    port map (
            O => \N__8463\,
            I => \N__8457\
        );

    \I__1821\ : Span4Mux_h
    port map (
            O => \N__8460\,
            I => \N__8454\
        );

    \I__1820\ : Span12Mux_h
    port map (
            O => \N__8457\,
            I => \N__8451\
        );

    \I__1819\ : Span4Mux_h
    port map (
            O => \N__8454\,
            I => \N__8448\
        );

    \I__1818\ : Odrv12
    port map (
            O => \N__8451\,
            I => \SIZ_c_1\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__8448\,
            I => \SIZ_c_1\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8443\,
            I => \N__8437\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8442\,
            I => \N__8432\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8441\,
            I => \N__8432\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8440\,
            I => \N__8429\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8437\,
            I => \N__8425\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8432\,
            I => \N__8417\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8429\,
            I => \N__8417\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8428\,
            I => \N__8414\
        );

    \I__1808\ : Span4Mux_v
    port map (
            O => \N__8425\,
            I => \N__8411\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8424\,
            I => \N__8404\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8404\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8404\
        );

    \I__1804\ : Span4Mux_v
    port map (
            O => \N__8417\,
            I => \N__8401\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8414\,
            I => \N__8398\
        );

    \I__1802\ : Span4Mux_v
    port map (
            O => \N__8411\,
            I => \N__8395\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8404\,
            I => \N__8392\
        );

    \I__1800\ : Span4Mux_v
    port map (
            O => \N__8401\,
            I => \N__8387\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__8398\,
            I => \N__8387\
        );

    \I__1798\ : Sp12to4
    port map (
            O => \N__8395\,
            I => \N__8380\
        );

    \I__1797\ : Span12Mux_s7_v
    port map (
            O => \N__8392\,
            I => \N__8380\
        );

    \I__1796\ : Sp12to4
    port map (
            O => \N__8387\,
            I => \N__8380\
        );

    \I__1795\ : Span12Mux_h
    port map (
            O => \N__8380\,
            I => \N__8377\
        );

    \I__1794\ : Odrv12
    port map (
            O => \N__8377\,
            I => \A_c_1\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__8374\,
            I => \N__8370\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8373\,
            I => \N__8365\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8365\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8365\,
            I => \N__8356\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__8364\,
            I => \N__8353\
        );

    \I__1788\ : InMux
    port map (
            O => \N__8363\,
            I => \N__8350\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8362\,
            I => \N__8347\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8361\,
            I => \N__8344\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__8360\,
            I => \N__8340\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__8359\,
            I => \N__8336\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__8356\,
            I => \N__8333\
        );

    \I__1782\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8330\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__8350\,
            I => \N__8327\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8347\,
            I => \N__8322\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8344\,
            I => \N__8322\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8315\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8340\,
            I => \N__8315\
        );

    \I__1776\ : InMux
    port map (
            O => \N__8339\,
            I => \N__8315\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8336\,
            I => \N__8312\
        );

    \I__1774\ : Span4Mux_v
    port map (
            O => \N__8333\,
            I => \N__8309\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__8330\,
            I => \N__8306\
        );

    \I__1772\ : Span4Mux_v
    port map (
            O => \N__8327\,
            I => \N__8303\
        );

    \I__1771\ : Span4Mux_v
    port map (
            O => \N__8322\,
            I => \N__8296\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8315\,
            I => \N__8296\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__8312\,
            I => \N__8296\
        );

    \I__1768\ : Span4Mux_v
    port map (
            O => \N__8309\,
            I => \N__8293\
        );

    \I__1767\ : Span4Mux_h
    port map (
            O => \N__8306\,
            I => \N__8290\
        );

    \I__1766\ : Span4Mux_v
    port map (
            O => \N__8303\,
            I => \N__8285\
        );

    \I__1765\ : Span4Mux_h
    port map (
            O => \N__8296\,
            I => \N__8285\
        );

    \I__1764\ : Span4Mux_h
    port map (
            O => \N__8293\,
            I => \N__8282\
        );

    \I__1763\ : Sp12to4
    port map (
            O => \N__8290\,
            I => \N__8279\
        );

    \I__1762\ : Span4Mux_v
    port map (
            O => \N__8285\,
            I => \N__8276\
        );

    \I__1761\ : Sp12to4
    port map (
            O => \N__8282\,
            I => \N__8269\
        );

    \I__1760\ : Span12Mux_v
    port map (
            O => \N__8279\,
            I => \N__8269\
        );

    \I__1759\ : Sp12to4
    port map (
            O => \N__8276\,
            I => \N__8269\
        );

    \I__1758\ : Odrv12
    port map (
            O => \N__8269\,
            I => \SIZ_c_0\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__8266\,
            I => \N__8257\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__8265\,
            I => \N__8253\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8264\,
            I => \N__8248\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8245\
        );

    \I__1753\ : InMux
    port map (
            O => \N__8262\,
            I => \N__8242\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8239\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__8260\,
            I => \N__8236\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8229\
        );

    \I__1749\ : InMux
    port map (
            O => \N__8256\,
            I => \N__8229\
        );

    \I__1748\ : InMux
    port map (
            O => \N__8253\,
            I => \N__8229\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8252\,
            I => \N__8226\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8251\,
            I => \N__8223\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8248\,
            I => \N__8220\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__8245\,
            I => \N__8217\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8242\,
            I => \N__8212\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__8239\,
            I => \N__8212\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8209\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__8229\,
            I => \N__8202\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8226\,
            I => \N__8202\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8223\,
            I => \N__8202\
        );

    \I__1737\ : Span4Mux_v
    port map (
            O => \N__8220\,
            I => \N__8197\
        );

    \I__1736\ : Span4Mux_v
    port map (
            O => \N__8217\,
            I => \N__8197\
        );

    \I__1735\ : Span4Mux_v
    port map (
            O => \N__8212\,
            I => \N__8194\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__8209\,
            I => \N__8191\
        );

    \I__1733\ : Span12Mux_s10_v
    port map (
            O => \N__8202\,
            I => \N__8188\
        );

    \I__1732\ : Span4Mux_h
    port map (
            O => \N__8197\,
            I => \N__8183\
        );

    \I__1731\ : Span4Mux_h
    port map (
            O => \N__8194\,
            I => \N__8183\
        );

    \I__1730\ : Span4Mux_v
    port map (
            O => \N__8191\,
            I => \N__8180\
        );

    \I__1729\ : Span12Mux_h
    port map (
            O => \N__8188\,
            I => \N__8177\
        );

    \I__1728\ : Sp12to4
    port map (
            O => \N__8183\,
            I => \N__8172\
        );

    \I__1727\ : Sp12to4
    port map (
            O => \N__8180\,
            I => \N__8172\
        );

    \I__1726\ : Odrv12
    port map (
            O => \N__8177\,
            I => \A_c_0\
        );

    \I__1725\ : Odrv12
    port map (
            O => \N__8172\,
            I => \A_c_0\
        );

    \I__1724\ : IoInMux
    port map (
            O => \N__8167\,
            I => \N__8164\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8164\,
            I => \N__8161\
        );

    \I__1722\ : Span4Mux_s3_v
    port map (
            O => \N__8161\,
            I => \N__8158\
        );

    \I__1721\ : Span4Mux_h
    port map (
            O => \N__8158\,
            I => \N__8155\
        );

    \I__1720\ : Odrv4
    port map (
            O => \N__8155\,
            I => \N_244_i\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8149\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__8149\,
            I => \N__8145\
        );

    \I__1717\ : InMux
    port map (
            O => \N__8148\,
            I => \N__8142\
        );

    \I__1716\ : Span4Mux_h
    port map (
            O => \N__8145\,
            I => \N__8139\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8142\,
            I => \N__8131\
        );

    \I__1714\ : Span4Mux_v
    port map (
            O => \N__8139\,
            I => \N__8131\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8138\,
            I => \N__8126\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8137\,
            I => \N__8126\
        );

    \I__1711\ : InMux
    port map (
            O => \N__8136\,
            I => \N__8121\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__8131\,
            I => \N__8118\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__8126\,
            I => \N__8115\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8110\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8110\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8121\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__8118\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1704\ : Odrv12
    port map (
            O => \N__8115\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__8110\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1702\ : IoInMux
    port map (
            O => \N__8101\,
            I => \N__8098\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8098\,
            I => \N__8095\
        );

    \I__1700\ : Span4Mux_s2_v
    port map (
            O => \N__8095\,
            I => \N__8092\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__8092\,
            I => \N__8089\
        );

    \I__1698\ : Span4Mux_h
    port map (
            O => \N__8089\,
            I => \N__8086\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__8086\,
            I => \RASn_c\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__8083\,
            I => \N__8080\
        );

    \I__1695\ : InMux
    port map (
            O => \N__8080\,
            I => \N__8076\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8079\,
            I => \N__8073\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8076\,
            I => \N__8069\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__8073\,
            I => \N__8066\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8072\,
            I => \N__8061\
        );

    \I__1690\ : Span4Mux_h
    port map (
            O => \N__8069\,
            I => \N__8058\
        );

    \I__1689\ : Span12Mux_v
    port map (
            O => \N__8066\,
            I => \N__8055\
        );

    \I__1688\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8052\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8049\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8061\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__8058\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1684\ : Odrv12
    port map (
            O => \N__8055\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8052\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__8049\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1681\ : IoInMux
    port map (
            O => \N__8038\,
            I => \N__8035\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__8035\,
            I => \N__8032\
        );

    \I__1679\ : Span4Mux_s3_v
    port map (
            O => \N__8032\,
            I => \N__8029\
        );

    \I__1678\ : Span4Mux_v
    port map (
            O => \N__8029\,
            I => \N__8026\
        );

    \I__1677\ : Sp12to4
    port map (
            O => \N__8026\,
            I => \N__8023\
        );

    \I__1676\ : Odrv12
    port map (
            O => \N__8023\,
            I => \CRCSn_c\
        );

    \I__1675\ : IoInMux
    port map (
            O => \N__8020\,
            I => \N__8017\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8017\,
            I => \N__8014\
        );

    \I__1673\ : IoSpan4Mux
    port map (
            O => \N__8014\,
            I => \N__8011\
        );

    \I__1672\ : Sp12to4
    port map (
            O => \N__8011\,
            I => \N__8008\
        );

    \I__1671\ : Span12Mux_s9_v
    port map (
            O => \N__8008\,
            I => \N__8005\
        );

    \I__1670\ : Odrv12
    port map (
            O => \N__8005\,
            I => \CASn_c\
        );

    \I__1669\ : InMux
    port map (
            O => \N__8002\,
            I => \N__7999\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__7999\,
            I => \N__7996\
        );

    \I__1667\ : Sp12to4
    port map (
            O => \N__7996\,
            I => \N__7993\
        );

    \I__1666\ : Span12Mux_v
    port map (
            O => \N__7993\,
            I => \N__7990\
        );

    \I__1665\ : Span12Mux_h
    port map (
            O => \N__7990\,
            I => \N__7987\
        );

    \I__1664\ : Odrv12
    port map (
            O => \N__7987\,
            I => \A_c_16\
        );

    \I__1663\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7981\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7981\,
            I => \N__7978\
        );

    \I__1661\ : Sp12to4
    port map (
            O => \N__7978\,
            I => \N__7975\
        );

    \I__1660\ : Span12Mux_v
    port map (
            O => \N__7975\,
            I => \N__7972\
        );

    \I__1659\ : Span12Mux_h
    port map (
            O => \N__7972\,
            I => \N__7969\
        );

    \I__1658\ : Odrv12
    port map (
            O => \N__7969\,
            I => \A_c_18\
        );

    \I__1657\ : InMux
    port map (
            O => \N__7966\,
            I => \N__7963\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__7963\,
            I => \N__7959\
        );

    \I__1655\ : InMux
    port map (
            O => \N__7962\,
            I => \N__7956\
        );

    \I__1654\ : Span4Mux_h
    port map (
            O => \N__7959\,
            I => \N__7948\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__7956\,
            I => \N__7948\
        );

    \I__1652\ : InMux
    port map (
            O => \N__7955\,
            I => \N__7943\
        );

    \I__1651\ : InMux
    port map (
            O => \N__7954\,
            I => \N__7943\
        );

    \I__1650\ : InMux
    port map (
            O => \N__7953\,
            I => \N__7938\
        );

    \I__1649\ : Span4Mux_v
    port map (
            O => \N__7948\,
            I => \N__7933\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__7943\,
            I => \N__7933\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7942\,
            I => \N__7930\
        );

    \I__1646\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7927\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__7938\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__7933\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7930\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__7927\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__7918\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\
        );

    \I__1640\ : InMux
    port map (
            O => \N__7915\,
            I => \N__7909\
        );

    \I__1639\ : InMux
    port map (
            O => \N__7914\,
            I => \N__7909\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__7909\,
            I => \N__7906\
        );

    \I__1637\ : Span4Mux_v
    port map (
            O => \N__7906\,
            I => \N__7903\
        );

    \I__1636\ : Sp12to4
    port map (
            O => \N__7903\,
            I => \N__7900\
        );

    \I__1635\ : Span12Mux_h
    port map (
            O => \N__7900\,
            I => \N__7897\
        );

    \I__1634\ : Span12Mux_v
    port map (
            O => \N__7897\,
            I => \N__7894\
        );

    \I__1633\ : Odrv12
    port map (
            O => \N__7894\,
            I => \A_c_14\
        );

    \I__1632\ : InMux
    port map (
            O => \N__7891\,
            I => \N__7888\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__7888\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\
        );

    \I__1630\ : InMux
    port map (
            O => \N__7885\,
            I => \N__7882\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__7882\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__7879\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\
        );

    \I__1627\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7873\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__7873\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1625\ : IoInMux
    port map (
            O => \N__7870\,
            I => \N__7867\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7867\,
            I => \N__7864\
        );

    \I__1623\ : Span12Mux_s8_v
    port map (
            O => \N__7864\,
            I => \N__7861\
        );

    \I__1622\ : Odrv12
    port map (
            O => \N__7861\,
            I => \CMA_c_1\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__7858\,
            I => \N__7855\
        );

    \I__1620\ : InMux
    port map (
            O => \N__7855\,
            I => \N__7852\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7852\,
            I => \U712_CHIP_RAM.N_333\
        );

    \I__1618\ : InMux
    port map (
            O => \N__7849\,
            I => \N__7846\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__7846\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__7843\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5_cascade_\
        );

    \I__1615\ : InMux
    port map (
            O => \N__7840\,
            I => \N__7837\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__7837\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1613\ : IoInMux
    port map (
            O => \N__7834\,
            I => \N__7831\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__7831\,
            I => \N__7828\
        );

    \I__1611\ : Span12Mux_s7_h
    port map (
            O => \N__7828\,
            I => \N__7825\
        );

    \I__1610\ : Span12Mux_v
    port map (
            O => \N__7825\,
            I => \N__7822\
        );

    \I__1609\ : Odrv12
    port map (
            O => \N__7822\,
            I => \CMA_c_5\
        );

    \I__1608\ : CascadeMux
    port map (
            O => \N__7819\,
            I => \N__7814\
        );

    \I__1607\ : InMux
    port map (
            O => \N__7818\,
            I => \N__7811\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7817\,
            I => \N__7808\
        );

    \I__1605\ : InMux
    port map (
            O => \N__7814\,
            I => \N__7805\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__7811\,
            I => \N__7796\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__7808\,
            I => \N__7796\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__7805\,
            I => \N__7793\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7804\,
            I => \N__7788\
        );

    \I__1600\ : InMux
    port map (
            O => \N__7803\,
            I => \N__7788\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7802\,
            I => \N__7785\
        );

    \I__1598\ : InMux
    port map (
            O => \N__7801\,
            I => \N__7782\
        );

    \I__1597\ : Odrv4
    port map (
            O => \N__7796\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__7793\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7788\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__7785\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__7782\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1592\ : InMux
    port map (
            O => \N__7771\,
            I => \N__7768\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__7768\,
            I => \N__7764\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7767\,
            I => \N__7761\
        );

    \I__1589\ : Span4Mux_h
    port map (
            O => \N__7764\,
            I => \N__7753\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__7761\,
            I => \N__7753\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7760\,
            I => \N__7750\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7759\,
            I => \N__7747\
        );

    \I__1585\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7744\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__7753\,
            I => \U712_REG_SM.N_367\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__7750\,
            I => \U712_REG_SM.N_367\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7747\,
            I => \U712_REG_SM.N_367\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__7744\,
            I => \U712_REG_SM.N_367\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__7735\,
            I => \N__7731\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7734\,
            I => \N__7728\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7731\,
            I => \N__7725\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7728\,
            I => \N__7722\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__7725\,
            I => \U712_REG_SM.N_374\
        );

    \I__1575\ : Odrv12
    port map (
            O => \N__7722\,
            I => \U712_REG_SM.N_374\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7717\,
            I => \N__7713\
        );

    \I__1573\ : InMux
    port map (
            O => \N__7716\,
            I => \N__7710\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__7713\,
            I => \U712_REG_SM.N_226\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__7710\,
            I => \U712_REG_SM.N_226\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7705\,
            I => \N__7701\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7704\,
            I => \N__7698\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7701\,
            I => \N__7695\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__7698\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1566\ : Odrv12
    port map (
            O => \N__7695\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1565\ : CascadeMux
    port map (
            O => \N__7690\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7687\,
            I => \N__7684\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__7684\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7681\,
            I => \N__7678\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7678\,
            I => \N__7675\
        );

    \I__1560\ : Span4Mux_v
    port map (
            O => \N__7675\,
            I => \N__7672\
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__7672\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__7669\,
            I => \N__7664\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__7668\,
            I => \N__7656\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__7667\,
            I => \N__7653\
        );

    \I__1555\ : InMux
    port map (
            O => \N__7664\,
            I => \N__7642\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7663\,
            I => \N__7635\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7662\,
            I => \N__7635\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7635\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__7660\,
            I => \N__7632\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7659\,
            I => \N__7627\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7656\,
            I => \N__7627\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7653\,
            I => \N__7622\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7652\,
            I => \N__7622\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__7651\,
            I => \N__7619\
        );

    \I__1545\ : CascadeMux
    port map (
            O => \N__7650\,
            I => \N__7616\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7649\,
            I => \N__7613\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__7648\,
            I => \N__7609\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7647\,
            I => \N__7605\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7646\,
            I => \N__7602\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7645\,
            I => \N__7599\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__7642\,
            I => \N__7594\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7635\,
            I => \N__7594\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7632\,
            I => \N__7591\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__7627\,
            I => \N__7586\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__7622\,
            I => \N__7586\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7619\,
            I => \N__7581\
        );

    \I__1533\ : InMux
    port map (
            O => \N__7616\,
            I => \N__7581\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__7613\,
            I => \N__7578\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7573\
        );

    \I__1530\ : InMux
    port map (
            O => \N__7609\,
            I => \N__7573\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7608\,
            I => \N__7570\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7605\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7602\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__7599\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__7594\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7591\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1523\ : Odrv4
    port map (
            O => \N__7586\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7581\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1521\ : Odrv4
    port map (
            O => \N__7578\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7573\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7570\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__7549\,
            I => \N__7542\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7548\,
            I => \N__7537\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__7547\,
            I => \N__7534\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7546\,
            I => \N__7527\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7520\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7542\,
            I => \N__7520\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7541\,
            I => \N__7520\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7540\,
            I => \N__7517\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7537\,
            I => \N__7512\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7534\,
            I => \N__7509\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7533\,
            I => \N__7502\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7532\,
            I => \N__7499\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7531\,
            I => \N__7496\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7530\,
            I => \N__7493\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7527\,
            I => \N__7488\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7520\,
            I => \N__7488\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7517\,
            I => \N__7485\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7480\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7515\,
            I => \N__7480\
        );

    \I__1499\ : Span4Mux_v
    port map (
            O => \N__7512\,
            I => \N__7475\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7509\,
            I => \N__7475\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7508\,
            I => \N__7470\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7507\,
            I => \N__7470\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7467\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7505\,
            I => \N__7464\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__7502\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7499\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7496\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__7493\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1489\ : Odrv4
    port map (
            O => \N__7488\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__7485\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7480\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1486\ : Odrv4
    port map (
            O => \N__7475\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7470\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7467\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7464\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7435\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7440\,
            I => \N__7429\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7439\,
            I => \N__7426\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7438\,
            I => \N__7423\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7435\,
            I => \N__7420\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7434\,
            I => \N__7417\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7433\,
            I => \N__7413\
        );

    \I__1475\ : CascadeMux
    port map (
            O => \N__7432\,
            I => \N__7409\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7429\,
            I => \N__7397\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7426\,
            I => \N__7397\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__7423\,
            I => \N__7397\
        );

    \I__1471\ : Span4Mux_v
    port map (
            O => \N__7420\,
            I => \N__7397\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7417\,
            I => \N__7397\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7416\,
            I => \N__7394\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7413\,
            I => \N__7391\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7412\,
            I => \N__7388\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7409\,
            I => \N__7385\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7408\,
            I => \N__7382\
        );

    \I__1464\ : Span4Mux_v
    port map (
            O => \N__7397\,
            I => \N__7379\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7394\,
            I => \N__7376\
        );

    \I__1462\ : Odrv12
    port map (
            O => \N__7391\,
            I => \U712_CHIP_RAM.N_358\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__7388\,
            I => \U712_CHIP_RAM.N_358\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__7385\,
            I => \U712_CHIP_RAM.N_358\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7382\,
            I => \U712_CHIP_RAM.N_358\
        );

    \I__1458\ : Odrv4
    port map (
            O => \N__7379\,
            I => \U712_CHIP_RAM.N_358\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__7376\,
            I => \U712_CHIP_RAM.N_358\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7363\,
            I => \N__7360\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7360\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_a3_0\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7357\,
            I => \N__7354\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7354\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1452\ : IoInMux
    port map (
            O => \N__7351\,
            I => \N__7348\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7348\,
            I => \N__7345\
        );

    \I__1450\ : Span12Mux_s8_h
    port map (
            O => \N__7345\,
            I => \N__7342\
        );

    \I__1449\ : Span12Mux_v
    port map (
            O => \N__7342\,
            I => \N__7339\
        );

    \I__1448\ : Odrv12
    port map (
            O => \N__7339\,
            I => \CMA_c_3\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7336\,
            I => \N__7333\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7333\,
            I => \N__7330\
        );

    \I__1445\ : Span12Mux_v
    port map (
            O => \N__7330\,
            I => \N__7327\
        );

    \I__1444\ : Span12Mux_h
    port map (
            O => \N__7327\,
            I => \N__7324\
        );

    \I__1443\ : Odrv12
    port map (
            O => \N__7324\,
            I => \A_c_7\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7321\,
            I => \N__7318\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7318\,
            I => \N__7315\
        );

    \I__1440\ : Odrv4
    port map (
            O => \N__7315\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i\
        );

    \I__1439\ : CascadeMux
    port map (
            O => \N__7312\,
            I => \U712_CHIP_RAM.CMA_5_0_8_cascade_\
        );

    \I__1438\ : CascadeMux
    port map (
            O => \N__7309\,
            I => \U712_REG_SM.N_222_cascade_\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7306\,
            I => \N__7301\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7305\,
            I => \N__7298\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7295\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__7301\,
            I => \N__7287\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7298\,
            I => \N__7280\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7295\,
            I => \N__7277\
        );

    \I__1431\ : ClkMux
    port map (
            O => \N__7294\,
            I => \N__7252\
        );

    \I__1430\ : ClkMux
    port map (
            O => \N__7293\,
            I => \N__7252\
        );

    \I__1429\ : ClkMux
    port map (
            O => \N__7292\,
            I => \N__7252\
        );

    \I__1428\ : ClkMux
    port map (
            O => \N__7291\,
            I => \N__7252\
        );

    \I__1427\ : ClkMux
    port map (
            O => \N__7290\,
            I => \N__7252\
        );

    \I__1426\ : Glb2LocalMux
    port map (
            O => \N__7287\,
            I => \N__7252\
        );

    \I__1425\ : ClkMux
    port map (
            O => \N__7286\,
            I => \N__7252\
        );

    \I__1424\ : ClkMux
    port map (
            O => \N__7285\,
            I => \N__7252\
        );

    \I__1423\ : ClkMux
    port map (
            O => \N__7284\,
            I => \N__7252\
        );

    \I__1422\ : ClkMux
    port map (
            O => \N__7283\,
            I => \N__7252\
        );

    \I__1421\ : Glb2LocalMux
    port map (
            O => \N__7280\,
            I => \N__7252\
        );

    \I__1420\ : Glb2LocalMux
    port map (
            O => \N__7277\,
            I => \N__7252\
        );

    \I__1419\ : GlobalMux
    port map (
            O => \N__7252\,
            I => \N__7249\
        );

    \I__1418\ : gio2CtrlBuf
    port map (
            O => \N__7249\,
            I => \C1_c_g\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7246\,
            I => \N__7243\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7243\,
            I => \N__7239\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7242\,
            I => \N__7236\
        );

    \I__1414\ : Odrv12
    port map (
            O => \N__7239\,
            I => \U712_REG_SM.N_241\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__7236\,
            I => \U712_REG_SM.N_241\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__7231\,
            I => \N__7228\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7228\,
            I => \N__7225\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__7225\,
            I => \U712_REG_SM.ASn_0_sqmuxa_1\
        );

    \I__1409\ : IoInMux
    port map (
            O => \N__7222\,
            I => \N__7219\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__7219\,
            I => \N__7216\
        );

    \I__1407\ : IoSpan4Mux
    port map (
            O => \N__7216\,
            I => \N__7213\
        );

    \I__1406\ : Span4Mux_s2_v
    port map (
            O => \N__7213\,
            I => \N__7209\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7212\,
            I => \N__7206\
        );

    \I__1404\ : Sp12to4
    port map (
            O => \N__7209\,
            I => \N__7203\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7206\,
            I => \N__7199\
        );

    \I__1402\ : Span12Mux_v
    port map (
            O => \N__7203\,
            I => \N__7196\
        );

    \I__1401\ : InMux
    port map (
            O => \N__7202\,
            I => \N__7193\
        );

    \I__1400\ : Span4Mux_v
    port map (
            O => \N__7199\,
            I => \N__7190\
        );

    \I__1399\ : Odrv12
    port map (
            O => \N__7196\,
            I => \REGENn_c\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__7193\,
            I => \REGENn_c\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__7190\,
            I => \REGENn_c\
        );

    \I__1396\ : InMux
    port map (
            O => \N__7183\,
            I => \N__7180\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7180\,
            I => \N__7176\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7179\,
            I => \N__7173\
        );

    \I__1393\ : Span4Mux_v
    port map (
            O => \N__7176\,
            I => \N__7170\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7173\,
            I => \N__7167\
        );

    \I__1391\ : Span4Mux_v
    port map (
            O => \N__7170\,
            I => \N__7164\
        );

    \I__1390\ : Span4Mux_v
    port map (
            O => \N__7167\,
            I => \N__7161\
        );

    \I__1389\ : Span4Mux_v
    port map (
            O => \N__7164\,
            I => \N__7156\
        );

    \I__1388\ : Span4Mux_v
    port map (
            O => \N__7161\,
            I => \N__7156\
        );

    \I__1387\ : Sp12to4
    port map (
            O => \N__7156\,
            I => \N__7153\
        );

    \I__1386\ : Span12Mux_h
    port map (
            O => \N__7153\,
            I => \N__7150\
        );

    \I__1385\ : Odrv12
    port map (
            O => \N__7150\,
            I => \TSn_c\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__7147\,
            I => \N__7144\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7144\,
            I => \N__7141\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__7141\,
            I => \N__7138\
        );

    \I__1381\ : Span4Mux_v
    port map (
            O => \N__7138\,
            I => \N__7135\
        );

    \I__1380\ : Sp12to4
    port map (
            O => \N__7135\,
            I => \N__7132\
        );

    \I__1379\ : Span12Mux_h
    port map (
            O => \N__7132\,
            I => \N__7129\
        );

    \I__1378\ : Span12Mux_v
    port map (
            O => \N__7129\,
            I => \N__7126\
        );

    \I__1377\ : Odrv12
    port map (
            O => \N__7126\,
            I => \REGSPACEn_c\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__7123\,
            I => \N__7119\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7122\,
            I => \N__7115\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7119\,
            I => \N__7112\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7109\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7115\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7112\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__7109\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1369\ : IoInMux
    port map (
            O => \N__7102\,
            I => \N__7099\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7099\,
            I => \N__7096\
        );

    \I__1367\ : IoSpan4Mux
    port map (
            O => \N__7096\,
            I => \N__7093\
        );

    \I__1366\ : IoSpan4Mux
    port map (
            O => \N__7093\,
            I => \N__7090\
        );

    \I__1365\ : Span4Mux_s2_v
    port map (
            O => \N__7090\,
            I => \N__7087\
        );

    \I__1364\ : Span4Mux_v
    port map (
            O => \N__7087\,
            I => \N__7084\
        );

    \I__1363\ : Odrv4
    port map (
            O => \N__7084\,
            I => \N_243_i\
        );

    \I__1362\ : IoInMux
    port map (
            O => \N__7081\,
            I => \N__7078\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__7078\,
            I => \N__7075\
        );

    \I__1360\ : Span4Mux_s3_v
    port map (
            O => \N__7075\,
            I => \N__7072\
        );

    \I__1359\ : Span4Mux_h
    port map (
            O => \N__7072\,
            I => \N__7069\
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__7069\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1357\ : IoInMux
    port map (
            O => \N__7066\,
            I => \N__7063\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7063\,
            I => \N__7060\
        );

    \I__1355\ : Span4Mux_s2_h
    port map (
            O => \N__7060\,
            I => \N__7057\
        );

    \I__1354\ : Span4Mux_h
    port map (
            O => \N__7057\,
            I => \N__7054\
        );

    \I__1353\ : Sp12to4
    port map (
            O => \N__7054\,
            I => \N__7051\
        );

    \I__1352\ : Span12Mux_s10_v
    port map (
            O => \N__7051\,
            I => \N__7048\
        );

    \I__1351\ : Odrv12
    port map (
            O => \N__7048\,
            I => \WEn_c\
        );

    \I__1350\ : IoInMux
    port map (
            O => \N__7045\,
            I => \N__7042\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__7042\,
            I => \N__7039\
        );

    \I__1348\ : Span4Mux_s0_v
    port map (
            O => \N__7039\,
            I => \N__7036\
        );

    \I__1347\ : Sp12to4
    port map (
            O => \N__7036\,
            I => \N__7033\
        );

    \I__1346\ : Span12Mux_h
    port map (
            O => \N__7033\,
            I => \N__7030\
        );

    \I__1345\ : Odrv12
    port map (
            O => \N__7030\,
            I => \CMA_c_10\
        );

    \I__1344\ : IoInMux
    port map (
            O => \N__7027\,
            I => \N__7024\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__7024\,
            I => \N__7021\
        );

    \I__1342\ : Span4Mux_s3_v
    port map (
            O => \N__7021\,
            I => \N__7018\
        );

    \I__1341\ : Span4Mux_v
    port map (
            O => \N__7018\,
            I => \N__7015\
        );

    \I__1340\ : Span4Mux_v
    port map (
            O => \N__7015\,
            I => \N__7012\
        );

    \I__1339\ : Odrv4
    port map (
            O => \N__7012\,
            I => \CMA_c_2\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7009\,
            I => \N__7006\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__7006\,
            I => \N__7003\
        );

    \I__1336\ : Span12Mux_v
    port map (
            O => \N__7003\,
            I => \N__7000\
        );

    \I__1335\ : Span12Mux_h
    port map (
            O => \N__7000\,
            I => \N__6997\
        );

    \I__1334\ : Odrv12
    port map (
            O => \N__6997\,
            I => \A_c_11\
        );

    \I__1333\ : InMux
    port map (
            O => \N__6994\,
            I => \N__6991\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6991\,
            I => \N__6988\
        );

    \I__1331\ : Span4Mux_v
    port map (
            O => \N__6988\,
            I => \N__6985\
        );

    \I__1330\ : Span4Mux_v
    port map (
            O => \N__6985\,
            I => \N__6982\
        );

    \I__1329\ : Sp12to4
    port map (
            O => \N__6982\,
            I => \N__6979\
        );

    \I__1328\ : Span12Mux_h
    port map (
            O => \N__6979\,
            I => \N__6976\
        );

    \I__1327\ : Odrv12
    port map (
            O => \N__6976\,
            I => \A_c_4\
        );

    \I__1326\ : IoInMux
    port map (
            O => \N__6973\,
            I => \N__6970\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__6970\,
            I => \N__6967\
        );

    \I__1324\ : IoSpan4Mux
    port map (
            O => \N__6967\,
            I => \N__6964\
        );

    \I__1323\ : IoSpan4Mux
    port map (
            O => \N__6964\,
            I => \N__6961\
        );

    \I__1322\ : Span4Mux_s3_h
    port map (
            O => \N__6961\,
            I => \N__6957\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6960\,
            I => \N__6954\
        );

    \I__1320\ : Span4Mux_h
    port map (
            O => \N__6957\,
            I => \N__6951\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6954\,
            I => \N__6948\
        );

    \I__1318\ : Sp12to4
    port map (
            O => \N__6951\,
            I => \N__6945\
        );

    \I__1317\ : Sp12to4
    port map (
            O => \N__6948\,
            I => \N__6942\
        );

    \I__1316\ : Span12Mux_h
    port map (
            O => \N__6945\,
            I => \N__6937\
        );

    \I__1315\ : Span12Mux_v
    port map (
            O => \N__6942\,
            I => \N__6937\
        );

    \I__1314\ : Span12Mux_h
    port map (
            O => \N__6937\,
            I => \N__6934\
        );

    \I__1313\ : Odrv12
    port map (
            O => \N__6934\,
            I => \C3_c\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6931\,
            I => \N__6928\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__6928\,
            I => \U712_REG_SM.N_313\
        );

    \I__1310\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6916\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6924\,
            I => \N__6916\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6913\
        );

    \I__1307\ : InMux
    port map (
            O => \N__6922\,
            I => \N__6908\
        );

    \I__1306\ : InMux
    port map (
            O => \N__6921\,
            I => \N__6908\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6916\,
            I => \U712_REG_SM.N_220\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__6913\,
            I => \U712_REG_SM.N_220\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6908\,
            I => \U712_REG_SM.N_220\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6901\,
            I => \N__6892\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6889\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6899\,
            I => \N__6886\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6898\,
            I => \N__6883\
        );

    \I__1298\ : InMux
    port map (
            O => \N__6897\,
            I => \N__6880\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6896\,
            I => \N__6875\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6895\,
            I => \N__6875\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__6892\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6889\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6886\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__6883\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__6880\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__6875\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__6862\,
            I => \U712_REG_SM.STATE_COUNTc_0_0_cascade_\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__6859\,
            I => \N__6856\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6856\,
            I => \N__6853\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__6853\,
            I => \N__6849\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6852\,
            I => \N__6846\
        );

    \I__1284\ : Span4Mux_v
    port map (
            O => \N__6849\,
            I => \N__6843\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6846\,
            I => \U712_REG_SM.N_266\
        );

    \I__1282\ : Odrv4
    port map (
            O => \N__6843\,
            I => \U712_REG_SM.N_266\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__6838\,
            I => \N__6835\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6830\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6834\,
            I => \N__6826\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6833\,
            I => \N__6823\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6830\,
            I => \N__6820\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6829\,
            I => \N__6817\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6826\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__6823\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1273\ : Odrv4
    port map (
            O => \N__6820\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6817\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1271\ : InMux
    port map (
            O => \N__6808\,
            I => \N__6804\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6807\,
            I => \N__6801\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__6804\,
            I => \N__6793\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6801\,
            I => \N__6793\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6800\,
            I => \N__6790\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6799\,
            I => \N__6785\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6798\,
            I => \N__6785\
        );

    \I__1264\ : Span4Mux_v
    port map (
            O => \N__6793\,
            I => \N__6782\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__6790\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__6785\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1261\ : Odrv4
    port map (
            O => \N__6782\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6762\
        );

    \I__1259\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6762\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6762\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6759\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6771\,
            I => \N__6756\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6770\,
            I => \N__6751\
        );

    \I__1254\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6751\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__6762\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__6759\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__6756\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6751\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6742\,
            I => \N__6739\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6739\,
            I => \U712_REG_SM.N_222\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__6736\,
            I => \N__6733\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6733\,
            I => \N__6728\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6732\,
            I => \N__6722\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6719\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__6728\,
            I => \N__6716\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6727\,
            I => \N__6713\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6726\,
            I => \N__6708\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6725\,
            I => \N__6708\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__6722\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6719\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__6716\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6713\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6708\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6697\,
            I => \N__6694\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6694\,
            I => \N__6691\
        );

    \I__1232\ : Sp12to4
    port map (
            O => \N__6691\,
            I => \N__6688\
        );

    \I__1231\ : Span12Mux_v
    port map (
            O => \N__6688\,
            I => \N__6685\
        );

    \I__1230\ : Span12Mux_h
    port map (
            O => \N__6685\,
            I => \N__6682\
        );

    \I__1229\ : Odrv12
    port map (
            O => \N__6682\,
            I => \A_c_5\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6676\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6676\,
            I => \N__6673\
        );

    \I__1226\ : Span4Mux_v
    port map (
            O => \N__6673\,
            I => \N__6670\
        );

    \I__1225\ : Sp12to4
    port map (
            O => \N__6670\,
            I => \N__6667\
        );

    \I__1224\ : Span12Mux_h
    port map (
            O => \N__6667\,
            I => \N__6664\
        );

    \I__1223\ : Odrv12
    port map (
            O => \N__6664\,
            I => \A_c_12\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__6661\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6658\,
            I => \N__6655\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6655\,
            I => \N__6652\
        );

    \I__1219\ : Span4Mux_v
    port map (
            O => \N__6652\,
            I => \N__6649\
        );

    \I__1218\ : Sp12to4
    port map (
            O => \N__6649\,
            I => \N__6646\
        );

    \I__1217\ : Span12Mux_h
    port map (
            O => \N__6646\,
            I => \N__6643\
        );

    \I__1216\ : Odrv12
    port map (
            O => \N__6643\,
            I => \A_c_10\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6637\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6637\,
            I => \N__6634\
        );

    \I__1213\ : Span4Mux_v
    port map (
            O => \N__6634\,
            I => \N__6631\
        );

    \I__1212\ : Sp12to4
    port map (
            O => \N__6631\,
            I => \N__6628\
        );

    \I__1211\ : Span12Mux_h
    port map (
            O => \N__6628\,
            I => \N__6625\
        );

    \I__1210\ : Span12Mux_v
    port map (
            O => \N__6625\,
            I => \N__6622\
        );

    \I__1209\ : Odrv12
    port map (
            O => \N__6622\,
            I => \A_c_3\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6616\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6616\,
            I => \N__6613\
        );

    \I__1206\ : Span4Mux_v
    port map (
            O => \N__6613\,
            I => \N__6610\
        );

    \I__1205\ : Sp12to4
    port map (
            O => \N__6610\,
            I => \N__6607\
        );

    \I__1204\ : Span12Mux_h
    port map (
            O => \N__6607\,
            I => \N__6604\
        );

    \I__1203\ : Span12Mux_v
    port map (
            O => \N__6604\,
            I => \N__6601\
        );

    \I__1202\ : Odrv12
    port map (
            O => \N__6601\,
            I => \A_c_15\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6598\,
            I => \N__6595\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6595\,
            I => \N__6592\
        );

    \I__1199\ : Span4Mux_v
    port map (
            O => \N__6592\,
            I => \N__6589\
        );

    \I__1198\ : Sp12to4
    port map (
            O => \N__6589\,
            I => \N__6586\
        );

    \I__1197\ : Span12Mux_h
    port map (
            O => \N__6586\,
            I => \N__6583\
        );

    \I__1196\ : Odrv12
    port map (
            O => \N__6583\,
            I => \A_c_8\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6580\,
            I => \N__6574\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6579\,
            I => \N__6569\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6578\,
            I => \N__6569\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6566\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__6574\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__6569\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__6566\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__6559\,
            I => \U712_REG_SM.N_269_cascade_\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6552\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__6555\,
            I => \N__6546\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6552\,
            I => \N__6543\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__6551\,
            I => \N__6540\
        );

    \I__1183\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6533\
        );

    \I__1182\ : InMux
    port map (
            O => \N__6549\,
            I => \N__6533\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6546\,
            I => \N__6533\
        );

    \I__1180\ : Span4Mux_h
    port map (
            O => \N__6543\,
            I => \N__6530\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6540\,
            I => \N__6527\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6533\,
            I => \N__6524\
        );

    \I__1177\ : Odrv4
    port map (
            O => \N__6530\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__6527\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1175\ : Odrv4
    port map (
            O => \N__6524\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6517\,
            I => \N__6514\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__6514\,
            I => \U712_REG_SM.DS_EN_RNOZ0Z_0\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__6511\,
            I => \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_cascade_\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6508\,
            I => \N__6504\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6507\,
            I => \N__6501\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6504\,
            I => \N__6496\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6501\,
            I => \N__6496\
        );

    \I__1167\ : Span4Mux_v
    port map (
            O => \N__6496\,
            I => \N__6493\
        );

    \I__1166\ : Span4Mux_v
    port map (
            O => \N__6493\,
            I => \N__6489\
        );

    \I__1165\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6486\
        );

    \I__1164\ : Sp12to4
    port map (
            O => \N__6489\,
            I => \N__6481\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6486\,
            I => \N__6481\
        );

    \I__1162\ : Span12Mux_h
    port map (
            O => \N__6481\,
            I => \N__6478\
        );

    \I__1161\ : Odrv12
    port map (
            O => \N__6478\,
            I => \DBRn_c\
        );

    \I__1160\ : IoInMux
    port map (
            O => \N__6475\,
            I => \N__6472\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6472\,
            I => \N__6469\
        );

    \I__1158\ : IoSpan4Mux
    port map (
            O => \N__6469\,
            I => \N__6466\
        );

    \I__1157\ : IoSpan4Mux
    port map (
            O => \N__6466\,
            I => \N__6463\
        );

    \I__1156\ : Span4Mux_s3_v
    port map (
            O => \N__6463\,
            I => \N__6460\
        );

    \I__1155\ : Span4Mux_v
    port map (
            O => \N__6460\,
            I => \N__6457\
        );

    \I__1154\ : Odrv4
    port map (
            O => \N__6457\,
            I => \DMA_LATCH_EN_c\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__6454\,
            I => \N__6449\
        );

    \I__1152\ : InMux
    port map (
            O => \N__6453\,
            I => \N__6441\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6452\,
            I => \N__6441\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6449\,
            I => \N__6436\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6448\,
            I => \N__6425\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6447\,
            I => \N__6425\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6425\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6441\,
            I => \N__6420\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6440\,
            I => \N__6409\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6439\,
            I => \N__6409\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6436\,
            I => \N__6406\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6435\,
            I => \N__6403\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6434\,
            I => \N__6396\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6433\,
            I => \N__6396\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6432\,
            I => \N__6396\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__6425\,
            I => \N__6393\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6424\,
            I => \N__6390\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6423\,
            I => \N__6387\
        );

    \I__1135\ : Span4Mux_h
    port map (
            O => \N__6420\,
            I => \N__6384\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6419\,
            I => \N__6381\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6378\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6417\,
            I => \N__6369\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6416\,
            I => \N__6369\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6415\,
            I => \N__6369\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6414\,
            I => \N__6369\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6409\,
            I => \N__6366\
        );

    \I__1127\ : Span4Mux_h
    port map (
            O => \N__6406\,
            I => \N__6357\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6403\,
            I => \N__6357\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6396\,
            I => \N__6357\
        );

    \I__1124\ : Span4Mux_h
    port map (
            O => \N__6393\,
            I => \N__6357\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6390\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6387\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1121\ : Odrv4
    port map (
            O => \N__6384\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__6381\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6378\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6369\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__6366\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1116\ : Odrv4
    port map (
            O => \N__6357\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__6340\,
            I => \N__6336\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6339\,
            I => \N__6330\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6327\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6321\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6334\,
            I => \N__6318\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6333\,
            I => \N__6315\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6330\,
            I => \N__6312\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6327\,
            I => \N__6305\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6302\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__6325\,
            I => \N__6299\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6324\,
            I => \N__6295\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6321\,
            I => \N__6286\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__6318\,
            I => \N__6286\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6315\,
            I => \N__6286\
        );

    \I__1101\ : Span4Mux_h
    port map (
            O => \N__6312\,
            I => \N__6286\
        );

    \I__1100\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6281\
        );

    \I__1099\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6281\
        );

    \I__1098\ : InMux
    port map (
            O => \N__6309\,
            I => \N__6276\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6308\,
            I => \N__6276\
        );

    \I__1096\ : Span4Mux_v
    port map (
            O => \N__6305\,
            I => \N__6271\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__6302\,
            I => \N__6271\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6299\,
            I => \N__6266\
        );

    \I__1093\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6266\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__6295\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\
        );

    \I__1091\ : Odrv4
    port map (
            O => \N__6286\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__6281\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__6276\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__6271\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__6266\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__6253\,
            I => \U712_CHIP_RAM.N_320_cascade_\
        );

    \I__1085\ : CascadeMux
    port map (
            O => \N__6250\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6244\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__6244\,
            I => \N__6240\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6237\
        );

    \I__1081\ : Span4Mux_v
    port map (
            O => \N__6240\,
            I => \N__6234\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__6237\,
            I => \U712_CHIP_RAM.N_414\
        );

    \I__1079\ : Odrv4
    port map (
            O => \N__6234\,
            I => \U712_CHIP_RAM.N_414\
        );

    \I__1078\ : CascadeMux
    port map (
            O => \N__6229\,
            I => \N__6226\
        );

    \I__1077\ : InMux
    port map (
            O => \N__6226\,
            I => \N__6223\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__6223\,
            I => \N__6220\
        );

    \I__1075\ : Odrv12
    port map (
            O => \N__6220\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_1\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6208\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6216\,
            I => \N__6208\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6215\,
            I => \N__6208\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__6208\,
            I => \N__6200\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6207\,
            I => \N__6197\
        );

    \I__1069\ : InMux
    port map (
            O => \N__6206\,
            I => \N__6194\
        );

    \I__1068\ : InMux
    port map (
            O => \N__6205\,
            I => \N__6187\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6187\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6187\
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__6200\,
            I => \U712_CHIP_RAM.N_48_0\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__6197\,
            I => \U712_CHIP_RAM.N_48_0\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__6194\,
            I => \U712_CHIP_RAM.N_48_0\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__6187\,
            I => \U712_CHIP_RAM.N_48_0\
        );

    \I__1061\ : CEMux
    port map (
            O => \N__6178\,
            I => \N__6174\
        );

    \I__1060\ : CEMux
    port map (
            O => \N__6177\,
            I => \N__6170\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6174\,
            I => \N__6167\
        );

    \I__1058\ : CEMux
    port map (
            O => \N__6173\,
            I => \N__6164\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6170\,
            I => \N__6161\
        );

    \I__1056\ : Sp12to4
    port map (
            O => \N__6167\,
            I => \N__6156\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__6164\,
            I => \N__6156\
        );

    \I__1054\ : Odrv12
    port map (
            O => \N__6161\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__1053\ : Odrv12
    port map (
            O => \N__6156\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__1052\ : InMux
    port map (
            O => \N__6151\,
            I => \N__6147\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__6150\,
            I => \N__6143\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6147\,
            I => \N__6139\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6146\,
            I => \N__6136\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6130\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6142\,
            I => \N__6126\
        );

    \I__1046\ : Span4Mux_h
    port map (
            O => \N__6139\,
            I => \N__6122\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__6136\,
            I => \N__6119\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__6135\,
            I => \N__6116\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6134\,
            I => \N__6111\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6111\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__6130\,
            I => \N__6108\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6129\,
            I => \N__6105\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__6126\,
            I => \N__6102\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6125\,
            I => \N__6094\
        );

    \I__1037\ : Span4Mux_v
    port map (
            O => \N__6122\,
            I => \N__6091\
        );

    \I__1036\ : Span4Mux_h
    port map (
            O => \N__6119\,
            I => \N__6088\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6116\,
            I => \N__6085\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6111\,
            I => \N__6078\
        );

    \I__1033\ : Span4Mux_h
    port map (
            O => \N__6108\,
            I => \N__6078\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6105\,
            I => \N__6078\
        );

    \I__1031\ : Span4Mux_h
    port map (
            O => \N__6102\,
            I => \N__6075\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6101\,
            I => \N__6066\
        );

    \I__1029\ : InMux
    port map (
            O => \N__6100\,
            I => \N__6066\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6099\,
            I => \N__6066\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6098\,
            I => \N__6066\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6063\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__6094\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1024\ : Odrv4
    port map (
            O => \N__6091\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1023\ : Odrv4
    port map (
            O => \N__6088\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6085\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__6078\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1020\ : Odrv4
    port map (
            O => \N__6075\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6066\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__6063\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6046\,
            I => \N__6043\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__6043\,
            I => \N__6038\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6042\,
            I => \N__6035\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6041\,
            I => \N__6032\
        );

    \I__1013\ : Odrv4
    port map (
            O => \N__6038\,
            I => \U712_CHIP_RAM.N_363\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6035\,
            I => \U712_CHIP_RAM.N_363\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__6032\,
            I => \U712_CHIP_RAM.N_363\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__6025\,
            I => \U712_CHIP_RAM.N_358_cascade_\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6022\,
            I => \N__6019\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6019\,
            I => \N__6016\
        );

    \I__1007\ : Odrv4
    port map (
            O => \N__6016\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_a3_1\
        );

    \I__1006\ : InMux
    port map (
            O => \N__6013\,
            I => \N__6007\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6012\,
            I => \N__5999\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6011\,
            I => \N__5995\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6010\,
            I => \N__5992\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6007\,
            I => \N__5988\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6006\,
            I => \N__5985\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6005\,
            I => \N__5978\
        );

    \I__999\ : InMux
    port map (
            O => \N__6004\,
            I => \N__5978\
        );

    \I__998\ : InMux
    port map (
            O => \N__6003\,
            I => \N__5978\
        );

    \I__997\ : InMux
    port map (
            O => \N__6002\,
            I => \N__5972\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5999\,
            I => \N__5969\
        );

    \I__995\ : InMux
    port map (
            O => \N__5998\,
            I => \N__5966\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5995\,
            I => \N__5963\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5992\,
            I => \N__5960\
        );

    \I__992\ : InMux
    port map (
            O => \N__5991\,
            I => \N__5957\
        );

    \I__991\ : Span4Mux_v
    port map (
            O => \N__5988\,
            I => \N__5950\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__5985\,
            I => \N__5950\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__5978\,
            I => \N__5950\
        );

    \I__988\ : InMux
    port map (
            O => \N__5977\,
            I => \N__5943\
        );

    \I__987\ : InMux
    port map (
            O => \N__5976\,
            I => \N__5943\
        );

    \I__986\ : InMux
    port map (
            O => \N__5975\,
            I => \N__5943\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__5972\,
            I => \U712_CHIP_RAM.N_357\
        );

    \I__984\ : Odrv4
    port map (
            O => \N__5969\,
            I => \U712_CHIP_RAM.N_357\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5966\,
            I => \U712_CHIP_RAM.N_357\
        );

    \I__982\ : Odrv4
    port map (
            O => \N__5963\,
            I => \U712_CHIP_RAM.N_357\
        );

    \I__981\ : Odrv4
    port map (
            O => \N__5960\,
            I => \U712_CHIP_RAM.N_357\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__5957\,
            I => \U712_CHIP_RAM.N_357\
        );

    \I__979\ : Odrv4
    port map (
            O => \N__5950\,
            I => \U712_CHIP_RAM.N_357\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5943\,
            I => \U712_CHIP_RAM.N_357\
        );

    \I__977\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5922\
        );

    \I__976\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5919\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__5922\,
            I => \N__5916\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__5919\,
            I => \N__5913\
        );

    \I__973\ : Span4Mux_h
    port map (
            O => \N__5916\,
            I => \N__5909\
        );

    \I__972\ : Span4Mux_h
    port map (
            O => \N__5913\,
            I => \N__5906\
        );

    \I__971\ : InMux
    port map (
            O => \N__5912\,
            I => \N__5903\
        );

    \I__970\ : Odrv4
    port map (
            O => \N__5909\,
            I => \U712_CHIP_RAM.N_413\
        );

    \I__969\ : Odrv4
    port map (
            O => \N__5906\,
            I => \U712_CHIP_RAM.N_413\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5903\,
            I => \U712_CHIP_RAM.N_413\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__5896\,
            I => \N__5892\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__5895\,
            I => \N__5885\
        );

    \I__965\ : InMux
    port map (
            O => \N__5892\,
            I => \N__5876\
        );

    \I__964\ : InMux
    port map (
            O => \N__5891\,
            I => \N__5876\
        );

    \I__963\ : InMux
    port map (
            O => \N__5890\,
            I => \N__5873\
        );

    \I__962\ : InMux
    port map (
            O => \N__5889\,
            I => \N__5870\
        );

    \I__961\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5866\
        );

    \I__960\ : InMux
    port map (
            O => \N__5885\,
            I => \N__5863\
        );

    \I__959\ : InMux
    port map (
            O => \N__5884\,
            I => \N__5856\
        );

    \I__958\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5856\
        );

    \I__957\ : InMux
    port map (
            O => \N__5882\,
            I => \N__5856\
        );

    \I__956\ : InMux
    port map (
            O => \N__5881\,
            I => \N__5853\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5876\,
            I => \N__5848\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5873\,
            I => \N__5843\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5870\,
            I => \N__5843\
        );

    \I__952\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5840\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__5866\,
            I => \N__5835\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5863\,
            I => \N__5835\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5856\,
            I => \N__5832\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5853\,
            I => \N__5826\
        );

    \I__947\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5822\
        );

    \I__946\ : InMux
    port map (
            O => \N__5851\,
            I => \N__5819\
        );

    \I__945\ : Span4Mux_h
    port map (
            O => \N__5848\,
            I => \N__5810\
        );

    \I__944\ : Span4Mux_v
    port map (
            O => \N__5843\,
            I => \N__5810\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__5840\,
            I => \N__5810\
        );

    \I__942\ : Span4Mux_v
    port map (
            O => \N__5835\,
            I => \N__5810\
        );

    \I__941\ : Span4Mux_h
    port map (
            O => \N__5832\,
            I => \N__5807\
        );

    \I__940\ : InMux
    port map (
            O => \N__5831\,
            I => \N__5800\
        );

    \I__939\ : InMux
    port map (
            O => \N__5830\,
            I => \N__5800\
        );

    \I__938\ : InMux
    port map (
            O => \N__5829\,
            I => \N__5800\
        );

    \I__937\ : Span4Mux_h
    port map (
            O => \N__5826\,
            I => \N__5797\
        );

    \I__936\ : InMux
    port map (
            O => \N__5825\,
            I => \N__5794\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__5822\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5819\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__5810\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__932\ : Odrv4
    port map (
            O => \N__5807\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5800\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__930\ : Odrv4
    port map (
            O => \N__5797\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5794\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__928\ : CEMux
    port map (
            O => \N__5779\,
            I => \N__5776\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__5776\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0\
        );

    \I__926\ : CascadeMux
    port map (
            O => \N__5773\,
            I => \U712_REG_SM.N_270_cascade_\
        );

    \I__925\ : IoInMux
    port map (
            O => \N__5770\,
            I => \N__5767\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5767\,
            I => \N__5764\
        );

    \I__923\ : Span4Mux_s3_h
    port map (
            O => \N__5764\,
            I => \N__5761\
        );

    \I__922\ : Span4Mux_v
    port map (
            O => \N__5761\,
            I => \N__5758\
        );

    \I__921\ : Span4Mux_v
    port map (
            O => \N__5758\,
            I => \N__5755\
        );

    \I__920\ : Sp12to4
    port map (
            O => \N__5755\,
            I => \N__5752\
        );

    \I__919\ : Span12Mux_s11_h
    port map (
            O => \N__5752\,
            I => \N__5749\
        );

    \I__918\ : Odrv12
    port map (
            O => \N__5749\,
            I => \N_202_i\
        );

    \I__917\ : InMux
    port map (
            O => \N__5746\,
            I => \N__5743\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5743\,
            I => \N__5740\
        );

    \I__915\ : Odrv4
    port map (
            O => \N__5740\,
            I => \U712_BYTE_ENABLE.N_242\
        );

    \I__914\ : IoInMux
    port map (
            O => \N__5737\,
            I => \N__5734\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5734\,
            I => \N__5731\
        );

    \I__912\ : IoSpan4Mux
    port map (
            O => \N__5731\,
            I => \N__5728\
        );

    \I__911\ : Sp12to4
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__910\ : Span12Mux_s7_v
    port map (
            O => \N__5725\,
            I => \N__5722\
        );

    \I__909\ : Odrv12
    port map (
            O => \N__5722\,
            I => \N_188_i\
        );

    \I__908\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5713\
        );

    \I__907\ : InMux
    port map (
            O => \N__5718\,
            I => \N__5713\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5713\,
            I => \N__5710\
        );

    \I__905\ : Odrv4
    port map (
            O => \N__5710\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0\
        );

    \I__904\ : IoInMux
    port map (
            O => \N__5707\,
            I => \N__5704\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5704\,
            I => \N__5701\
        );

    \I__902\ : Span4Mux_s1_h
    port map (
            O => \N__5701\,
            I => \N__5698\
        );

    \I__901\ : Sp12to4
    port map (
            O => \N__5698\,
            I => \N__5695\
        );

    \I__900\ : Span12Mux_s5_v
    port map (
            O => \N__5695\,
            I => \N__5692\
        );

    \I__899\ : Span12Mux_h
    port map (
            O => \N__5692\,
            I => \N__5689\
        );

    \I__898\ : Span12Mux_v
    port map (
            O => \N__5689\,
            I => \N__5686\
        );

    \I__897\ : Odrv12
    port map (
            O => \N__5686\,
            I => \N_203_i\
        );

    \I__896\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5677\
        );

    \I__895\ : InMux
    port map (
            O => \N__5682\,
            I => \N__5677\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__5677\,
            I => \N__5674\
        );

    \I__893\ : Span4Mux_v
    port map (
            O => \N__5674\,
            I => \N__5671\
        );

    \I__892\ : Odrv4
    port map (
            O => \N__5671\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0\
        );

    \I__891\ : IoInMux
    port map (
            O => \N__5668\,
            I => \N__5665\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5665\,
            I => \N__5662\
        );

    \I__889\ : Span4Mux_s2_h
    port map (
            O => \N__5662\,
            I => \N__5659\
        );

    \I__888\ : Span4Mux_h
    port map (
            O => \N__5659\,
            I => \N__5656\
        );

    \I__887\ : Sp12to4
    port map (
            O => \N__5656\,
            I => \N__5653\
        );

    \I__886\ : Span12Mux_s10_v
    port map (
            O => \N__5653\,
            I => \N__5650\
        );

    \I__885\ : Span12Mux_h
    port map (
            O => \N__5650\,
            I => \N__5647\
        );

    \I__884\ : Odrv12
    port map (
            O => \N__5647\,
            I => \N_186_i\
        );

    \I__883\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5638\
        );

    \I__882\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5638\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5638\,
            I => \N__5635\
        );

    \I__880\ : Span4Mux_h
    port map (
            O => \N__5635\,
            I => \N__5632\
        );

    \I__879\ : Span4Mux_v
    port map (
            O => \N__5632\,
            I => \N__5629\
        );

    \I__878\ : Odrv4
    port map (
            O => \N__5629\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__5626\,
            I => \N__5623\
        );

    \I__876\ : InMux
    port map (
            O => \N__5623\,
            I => \N__5620\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5620\,
            I => \U712_BYTE_ENABLE.N_243\
        );

    \I__874\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5614\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5614\,
            I => \U712_BYTE_ENABLE.N_244\
        );

    \I__872\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5608\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5608\,
            I => \N__5605\
        );

    \I__870\ : Odrv4
    port map (
            O => \N__5605\,
            I => \U712_BYTE_ENABLE.N_245\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__5602\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_i_o2_0_1_3_cascade_\
        );

    \I__868\ : CascadeMux
    port map (
            O => \N__5599\,
            I => \U712_REG_SM.N_272_cascade_\
        );

    \I__867\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5593\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5593\,
            I => \U712_CHIP_RAM.N_236\
        );

    \I__865\ : InMux
    port map (
            O => \N__5590\,
            I => \N__5587\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5587\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__5584\,
            I => \N__5581\
        );

    \I__862\ : InMux
    port map (
            O => \N__5581\,
            I => \N__5578\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5578\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_i_0_i_0\
        );

    \I__860\ : InMux
    port map (
            O => \N__5575\,
            I => \N__5566\
        );

    \I__859\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5566\
        );

    \I__858\ : InMux
    port map (
            O => \N__5573\,
            I => \N__5566\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__5566\,
            I => \U712_CHIP_RAM.N_234\
        );

    \I__856\ : SRMux
    port map (
            O => \N__5563\,
            I => \N__5560\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__5560\,
            I => \N__5557\
        );

    \I__854\ : Odrv12
    port map (
            O => \N__5557\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__853\ : InMux
    port map (
            O => \N__5554\,
            I => \N__5551\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5551\,
            I => \N__5548\
        );

    \I__851\ : Span4Mux_h
    port map (
            O => \N__5548\,
            I => \N__5545\
        );

    \I__850\ : Sp12to4
    port map (
            O => \N__5545\,
            I => \N__5542\
        );

    \I__849\ : Span12Mux_v
    port map (
            O => \N__5542\,
            I => \N__5539\
        );

    \I__848\ : Odrv12
    port map (
            O => \N__5539\,
            I => \A_c_17\
        );

    \I__847\ : IoInMux
    port map (
            O => \N__5536\,
            I => \N__5533\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5533\,
            I => \N__5530\
        );

    \I__845\ : IoSpan4Mux
    port map (
            O => \N__5530\,
            I => \N__5527\
        );

    \I__844\ : Sp12to4
    port map (
            O => \N__5527\,
            I => \N__5524\
        );

    \I__843\ : Span12Mux_s9_h
    port map (
            O => \N__5524\,
            I => \N__5521\
        );

    \I__842\ : Span12Mux_v
    port map (
            O => \N__5521\,
            I => \N__5518\
        );

    \I__841\ : Odrv12
    port map (
            O => \N__5518\,
            I => \CMA_c_8\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__5515\,
            I => \N__5512\
        );

    \I__839\ : InMux
    port map (
            O => \N__5512\,
            I => \N__5509\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5509\,
            I => \N__5506\
        );

    \I__837\ : Span4Mux_v
    port map (
            O => \N__5506\,
            I => \N__5499\
        );

    \I__836\ : InMux
    port map (
            O => \N__5505\,
            I => \N__5494\
        );

    \I__835\ : InMux
    port map (
            O => \N__5504\,
            I => \N__5494\
        );

    \I__834\ : InMux
    port map (
            O => \N__5503\,
            I => \N__5489\
        );

    \I__833\ : InMux
    port map (
            O => \N__5502\,
            I => \N__5489\
        );

    \I__832\ : Odrv4
    port map (
            O => \N__5499\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5494\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5489\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__829\ : InMux
    port map (
            O => \N__5482\,
            I => \N__5479\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5479\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_0\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__5476\,
            I => \N__5471\
        );

    \I__826\ : InMux
    port map (
            O => \N__5475\,
            I => \N__5466\
        );

    \I__825\ : InMux
    port map (
            O => \N__5474\,
            I => \N__5466\
        );

    \I__824\ : InMux
    port map (
            O => \N__5471\,
            I => \N__5463\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__5466\,
            I => \N__5456\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5463\,
            I => \N__5456\
        );

    \I__821\ : InMux
    port map (
            O => \N__5462\,
            I => \N__5451\
        );

    \I__820\ : InMux
    port map (
            O => \N__5461\,
            I => \N__5451\
        );

    \I__819\ : Span4Mux_h
    port map (
            O => \N__5456\,
            I => \N__5448\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5451\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__817\ : Odrv4
    port map (
            O => \N__5448\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__5443\,
            I => \N__5439\
        );

    \I__815\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5434\
        );

    \I__814\ : InMux
    port map (
            O => \N__5439\,
            I => \N__5434\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5434\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__5431\,
            I => \U712_CHIP_RAM.N_236_cascade_\
        );

    \I__811\ : InMux
    port map (
            O => \N__5428\,
            I => \N__5425\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__5425\,
            I => \N__5421\
        );

    \I__809\ : InMux
    port map (
            O => \N__5424\,
            I => \N__5417\
        );

    \I__808\ : Span4Mux_h
    port map (
            O => \N__5421\,
            I => \N__5414\
        );

    \I__807\ : InMux
    port map (
            O => \N__5420\,
            I => \N__5411\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5417\,
            I => \U712_CHIP_RAM.N_274\
        );

    \I__805\ : Odrv4
    port map (
            O => \N__5414\,
            I => \U712_CHIP_RAM.N_274\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5411\,
            I => \U712_CHIP_RAM.N_274\
        );

    \I__803\ : CascadeMux
    port map (
            O => \N__5404\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\
        );

    \I__802\ : InMux
    port map (
            O => \N__5401\,
            I => \N__5398\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5398\,
            I => \N__5394\
        );

    \I__800\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5391\
        );

    \I__799\ : Span4Mux_v
    port map (
            O => \N__5394\,
            I => \N__5388\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5391\,
            I => \N__5385\
        );

    \I__797\ : Odrv4
    port map (
            O => \N__5388\,
            I => \U712_CHIP_RAM.N_366\
        );

    \I__796\ : Odrv4
    port map (
            O => \N__5385\,
            I => \U712_CHIP_RAM.N_366\
        );

    \I__795\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5377\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__5377\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a2_2_0_a3_0\
        );

    \I__793\ : InMux
    port map (
            O => \N__5374\,
            I => \N__5371\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5371\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__791\ : InMux
    port map (
            O => \N__5368\,
            I => \N__5365\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5365\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a3_0_1\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__5362\,
            I => \U712_CHIP_RAM.N_252_cascade_\
        );

    \I__788\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5356\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5356\,
            I => \U712_CHIP_RAM.N_286\
        );

    \I__786\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5350\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5350\,
            I => \N__5347\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__5347\,
            I => \U712_CHIP_RAM.N_267\
        );

    \I__783\ : InMux
    port map (
            O => \N__5344\,
            I => \N__5338\
        );

    \I__782\ : InMux
    port map (
            O => \N__5343\,
            I => \N__5338\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5338\,
            I => \U712_CHIP_RAM.N_225_i\
        );

    \I__780\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5332\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5332\,
            I => \U712_REG_SM.N_52\
        );

    \I__778\ : InMux
    port map (
            O => \N__5329\,
            I => \N__5326\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5326\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\
        );

    \I__776\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5319\
        );

    \I__775\ : InMux
    port map (
            O => \N__5322\,
            I => \N__5316\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5319\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__5316\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__5311\,
            I => \N__5306\
        );

    \I__771\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5303\
        );

    \I__770\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5299\
        );

    \I__769\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5296\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5303\,
            I => \N__5293\
        );

    \I__767\ : InMux
    port map (
            O => \N__5302\,
            I => \N__5290\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5299\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__5296\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__764\ : Odrv4
    port map (
            O => \N__5293\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__5290\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__762\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5277\
        );

    \I__761\ : InMux
    port map (
            O => \N__5280\,
            I => \N__5274\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__5277\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5274\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__5269\,
            I => \N__5264\
        );

    \I__757\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5260\
        );

    \I__756\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5257\
        );

    \I__755\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5254\
        );

    \I__754\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5251\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5260\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__5257\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__5254\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__5251\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__749\ : InMux
    port map (
            O => \N__5242\,
            I => \N__5239\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5239\,
            I => \N__5235\
        );

    \I__747\ : IoInMux
    port map (
            O => \N__5238\,
            I => \N__5232\
        );

    \I__746\ : Span4Mux_v
    port map (
            O => \N__5235\,
            I => \N__5229\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__5232\,
            I => \N__5226\
        );

    \I__744\ : Sp12to4
    port map (
            O => \N__5229\,
            I => \N__5223\
        );

    \I__743\ : IoSpan4Mux
    port map (
            O => \N__5226\,
            I => \N__5220\
        );

    \I__742\ : Span12Mux_h
    port map (
            O => \N__5223\,
            I => \N__5217\
        );

    \I__741\ : IoSpan4Mux
    port map (
            O => \N__5220\,
            I => \N__5214\
        );

    \I__740\ : Span12Mux_v
    port map (
            O => \N__5217\,
            I => \N__5211\
        );

    \I__739\ : IoSpan4Mux
    port map (
            O => \N__5214\,
            I => \N__5208\
        );

    \I__738\ : Odrv12
    port map (
            O => \N__5211\,
            I => \C1_c\
        );

    \I__737\ : Odrv4
    port map (
            O => \N__5208\,
            I => \C1_c\
        );

    \I__736\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5199\
        );

    \I__735\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5196\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__5199\,
            I => \N__5193\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5196\,
            I => \N__5190\
        );

    \I__732\ : Span4Mux_v
    port map (
            O => \N__5193\,
            I => \N__5187\
        );

    \I__731\ : Span4Mux_v
    port map (
            O => \N__5190\,
            I => \N__5184\
        );

    \I__730\ : Sp12to4
    port map (
            O => \N__5187\,
            I => \N__5181\
        );

    \I__729\ : Span4Mux_h
    port map (
            O => \N__5184\,
            I => \N__5178\
        );

    \I__728\ : Span12Mux_h
    port map (
            O => \N__5181\,
            I => \N__5175\
        );

    \I__727\ : Sp12to4
    port map (
            O => \N__5178\,
            I => \N__5172\
        );

    \I__726\ : Span12Mux_v
    port map (
            O => \N__5175\,
            I => \N__5169\
        );

    \I__725\ : Span12Mux_v
    port map (
            O => \N__5172\,
            I => \N__5166\
        );

    \I__724\ : Odrv12
    port map (
            O => \N__5169\,
            I => \AWEn_c\
        );

    \I__723\ : Odrv12
    port map (
            O => \N__5166\,
            I => \AWEn_c\
        );

    \I__722\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5155\
        );

    \I__721\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5152\
        );

    \I__720\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5149\
        );

    \I__719\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5139\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5155\,
            I => \N__5136\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5152\,
            I => \N__5131\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5149\,
            I => \N__5131\
        );

    \I__715\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5126\
        );

    \I__714\ : InMux
    port map (
            O => \N__5147\,
            I => \N__5126\
        );

    \I__713\ : InMux
    port map (
            O => \N__5146\,
            I => \N__5121\
        );

    \I__712\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5121\
        );

    \I__711\ : InMux
    port map (
            O => \N__5144\,
            I => \N__5114\
        );

    \I__710\ : InMux
    port map (
            O => \N__5143\,
            I => \N__5114\
        );

    \I__709\ : InMux
    port map (
            O => \N__5142\,
            I => \N__5114\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__5139\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__707\ : Odrv4
    port map (
            O => \N__5136\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__706\ : Odrv12
    port map (
            O => \N__5131\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5126\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5121\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__5114\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__702\ : CEMux
    port map (
            O => \N__5101\,
            I => \N__5098\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5098\,
            I => \N__5095\
        );

    \I__700\ : Span4Mux_v
    port map (
            O => \N__5095\,
            I => \N__5092\
        );

    \I__699\ : Odrv4
    port map (
            O => \N__5092\,
            I => \U712_CHIP_RAM.N_414_0\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__5089\,
            I => \U712_CHIP_RAM.N_363_cascade_\
        );

    \I__697\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5082\
        );

    \I__696\ : InMux
    port map (
            O => \N__5085\,
            I => \N__5079\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__5082\,
            I => \U712_CHIP_RAM.N_282\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__5079\,
            I => \U712_CHIP_RAM.N_282\
        );

    \I__693\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5071\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5071\,
            I => \U712_CHIP_RAM.N_292\
        );

    \I__691\ : InMux
    port map (
            O => \N__5068\,
            I => \N__5065\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__5065\,
            I => \U712_CHIP_RAM.N_347\
        );

    \I__689\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5059\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__5059\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0\
        );

    \I__687\ : IoInMux
    port map (
            O => \N__5056\,
            I => \N__5053\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5053\,
            I => \N__5050\
        );

    \I__685\ : Span12Mux_s2_v
    port map (
            O => \N__5050\,
            I => \N__5047\
        );

    \I__684\ : Span12Mux_v
    port map (
            O => \N__5047\,
            I => \N__5041\
        );

    \I__683\ : InMux
    port map (
            O => \N__5046\,
            I => \N__5038\
        );

    \I__682\ : InMux
    port map (
            O => \N__5045\,
            I => \N__5035\
        );

    \I__681\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5032\
        );

    \I__680\ : Odrv12
    port map (
            O => \N__5041\,
            I => \DBENn_c\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5038\,
            I => \DBENn_c\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__5035\,
            I => \DBENn_c\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5032\,
            I => \DBENn_c\
        );

    \I__676\ : InMux
    port map (
            O => \N__5023\,
            I => \N__5018\
        );

    \I__675\ : InMux
    port map (
            O => \N__5022\,
            I => \N__5013\
        );

    \I__674\ : InMux
    port map (
            O => \N__5021\,
            I => \N__5013\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__5018\,
            I => \N__5010\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__5013\,
            I => \N__5006\
        );

    \I__671\ : Span4Mux_v
    port map (
            O => \N__5010\,
            I => \N__5001\
        );

    \I__670\ : InMux
    port map (
            O => \N__5009\,
            I => \N__4998\
        );

    \I__669\ : Span4Mux_v
    port map (
            O => \N__5006\,
            I => \N__4995\
        );

    \I__668\ : InMux
    port map (
            O => \N__5005\,
            I => \N__4992\
        );

    \I__667\ : InMux
    port map (
            O => \N__5004\,
            I => \N__4989\
        );

    \I__666\ : Odrv4
    port map (
            O => \N__5001\,
            I => \DMA_CYCLEm\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4998\,
            I => \DMA_CYCLEm\
        );

    \I__664\ : Odrv4
    port map (
            O => \N__4995\,
            I => \DMA_CYCLEm\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4992\,
            I => \DMA_CYCLEm\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__4989\,
            I => \DMA_CYCLEm\
        );

    \I__661\ : InMux
    port map (
            O => \N__4978\,
            I => \N__4975\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4975\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_1_0\
        );

    \I__659\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4969\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4969\,
            I => \U712_REG_SM.N_304\
        );

    \I__657\ : InMux
    port map (
            O => \N__4966\,
            I => \N__4960\
        );

    \I__656\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4960\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__4960\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__654\ : InMux
    port map (
            O => \N__4957\,
            I => \N__4954\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4954\,
            I => \N__4950\
        );

    \I__652\ : InMux
    port map (
            O => \N__4953\,
            I => \N__4946\
        );

    \I__651\ : Span4Mux_h
    port map (
            O => \N__4950\,
            I => \N__4943\
        );

    \I__650\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4940\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__4946\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__648\ : Odrv4
    port map (
            O => \N__4943\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__4940\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__646\ : InMux
    port map (
            O => \N__4933\,
            I => \N__4930\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4930\,
            I => \U712_CYCLE_TERM.N_340\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__4927\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3T4KZ0Z7_cascade_\
        );

    \I__643\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4921\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__4921\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__4918\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__4915\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_0_cascade_\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__4912\,
            I => \U712_CHIP_RAM.N_284_cascade_\
        );

    \I__638\ : InMux
    port map (
            O => \N__4909\,
            I => \N__4906\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4906\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_2\
        );

    \I__636\ : InMux
    port map (
            O => \N__4903\,
            I => \N__4900\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4900\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2\
        );

    \I__634\ : InMux
    port map (
            O => \N__4897\,
            I => \N__4892\
        );

    \I__633\ : InMux
    port map (
            O => \N__4896\,
            I => \N__4887\
        );

    \I__632\ : InMux
    port map (
            O => \N__4895\,
            I => \N__4887\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4892\,
            I => \N__4884\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4887\,
            I => \N__4881\
        );

    \I__629\ : Odrv4
    port map (
            O => \N__4884\,
            I => \U712_CHIP_RAM.N_230\
        );

    \I__628\ : Odrv4
    port map (
            O => \N__4881\,
            I => \U712_CHIP_RAM.N_230\
        );

    \I__627\ : CascadeMux
    port map (
            O => \N__4876\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2_cascade_\
        );

    \I__626\ : InMux
    port map (
            O => \N__4873\,
            I => \N__4870\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4870\,
            I => \U712_CHIP_RAM.N_271\
        );

    \I__624\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4862\
        );

    \I__623\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4857\
        );

    \I__622\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4857\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__4862\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__4857\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__4852\,
            I => \U712_CHIP_RAM.N_271_cascade_\
        );

    \I__618\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4846\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__4846\,
            I => \N__4843\
        );

    \I__616\ : Odrv4
    port map (
            O => \N__4843\,
            I => \U712_CHIP_RAM.CLK_EN_5_0\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__4840\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_0_a2_i_1_cascade_\
        );

    \I__614\ : IoInMux
    port map (
            O => \N__4837\,
            I => \N__4834\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__4834\,
            I => \N__4831\
        );

    \I__612\ : Span4Mux_s2_h
    port map (
            O => \N__4831\,
            I => \N__4828\
        );

    \I__611\ : Span4Mux_v
    port map (
            O => \N__4828\,
            I => \N__4825\
        );

    \I__610\ : Span4Mux_v
    port map (
            O => \N__4825\,
            I => \N__4822\
        );

    \I__609\ : Sp12to4
    port map (
            O => \N__4822\,
            I => \N__4819\
        );

    \I__608\ : Span12Mux_h
    port map (
            O => \N__4819\,
            I => \N__4815\
        );

    \I__607\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4812\
        );

    \I__606\ : Odrv12
    port map (
            O => \N__4815\,
            I => \CLK_EN_c\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4812\,
            I => \CLK_EN_c\
        );

    \I__604\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4803\
        );

    \I__603\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4800\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4803\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__4800\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__600\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4791\
        );

    \I__599\ : InMux
    port map (
            O => \N__4794\,
            I => \N__4788\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__4791\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4788\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__4783\,
            I => \N__4779\
        );

    \I__595\ : InMux
    port map (
            O => \N__4782\,
            I => \N__4776\
        );

    \I__594\ : InMux
    port map (
            O => \N__4779\,
            I => \N__4773\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4776\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4773\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__591\ : InMux
    port map (
            O => \N__4768\,
            I => \N__4764\
        );

    \I__590\ : InMux
    port map (
            O => \N__4767\,
            I => \N__4761\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4764\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4761\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__4756\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7_cascade_\
        );

    \I__586\ : CascadeMux
    port map (
            O => \N__4753\,
            I => \U712_CHIP_RAM.N_230_cascade_\
        );

    \I__585\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4747\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4747\,
            I => \N__4744\
        );

    \I__583\ : Odrv4
    port map (
            O => \N__4744\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a3_1_1\
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__4741\,
            I => \U712_CHIP_RAM.N_287_cascade_\
        );

    \I__581\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4735\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4735\,
            I => \U712_CHIP_RAM.N_217\
        );

    \I__579\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4729\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4729\,
            I => \U712_CHIP_RAM.N_22\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__4726\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_113_tz_0_cascade_\
        );

    \I__576\ : InMux
    port map (
            O => \N__4723\,
            I => \bfn_9_7_0_\
        );

    \I__575\ : InMux
    port map (
            O => \N__4720\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__574\ : InMux
    port map (
            O => \N__4717\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__573\ : InMux
    port map (
            O => \N__4714\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__572\ : InMux
    port map (
            O => \N__4711\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__571\ : InMux
    port map (
            O => \N__4708\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__570\ : InMux
    port map (
            O => \N__4705\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__569\ : InMux
    port map (
            O => \N__4702\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__568\ : CEMux
    port map (
            O => \N__4699\,
            I => \N__4696\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4696\,
            I => \N__4693\
        );

    \I__566\ : Span4Mux_v
    port map (
            O => \N__4693\,
            I => \N__4690\
        );

    \I__565\ : Span4Mux_h
    port map (
            O => \N__4690\,
            I => \N__4687\
        );

    \I__564\ : Odrv4
    port map (
            O => \N__4687\,
            I => \U712_CYCLE_TERM.N_239_i_0_en_0\
        );

    \I__563\ : InMux
    port map (
            O => \N__4684\,
            I => \N__4681\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4681\,
            I => \N__4678\
        );

    \I__561\ : Span4Mux_v
    port map (
            O => \N__4678\,
            I => \N__4675\
        );

    \I__560\ : Sp12to4
    port map (
            O => \N__4675\,
            I => \N__4672\
        );

    \I__559\ : Span12Mux_h
    port map (
            O => \N__4672\,
            I => \N__4669\
        );

    \I__558\ : Odrv12
    port map (
            O => \N__4669\,
            I => \A_c_20\
        );

    \I__557\ : InMux
    port map (
            O => \N__4666\,
            I => \N__4663\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4663\,
            I => \N__4660\
        );

    \I__555\ : Odrv12
    port map (
            O => \N__4660\,
            I => \U712_CHIP_RAM.BANK0_RNOZ0Z_1\
        );

    \I__554\ : IoInMux
    port map (
            O => \N__4657\,
            I => \N__4654\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__4654\,
            I => \N__4651\
        );

    \I__552\ : Span4Mux_s3_v
    port map (
            O => \N__4651\,
            I => \N__4648\
        );

    \I__551\ : Span4Mux_v
    port map (
            O => \N__4648\,
            I => \N__4645\
        );

    \I__550\ : Span4Mux_v
    port map (
            O => \N__4645\,
            I => \N__4642\
        );

    \I__549\ : Odrv4
    port map (
            O => \N__4642\,
            I => \VBENn_c\
        );

    \I__548\ : InMux
    port map (
            O => \N__4639\,
            I => \N__4636\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4636\,
            I => \N__4632\
        );

    \I__546\ : InMux
    port map (
            O => \N__4635\,
            I => \N__4629\
        );

    \I__545\ : Span4Mux_h
    port map (
            O => \N__4632\,
            I => \N__4626\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4629\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__543\ : Odrv4
    port map (
            O => \N__4626\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__4621\,
            I => \N__4618\
        );

    \I__541\ : InMux
    port map (
            O => \N__4618\,
            I => \N__4615\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4615\,
            I => \N__4612\
        );

    \I__539\ : Span4Mux_v
    port map (
            O => \N__4612\,
            I => \N__4609\
        );

    \I__538\ : Odrv4
    port map (
            O => \N__4609\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__537\ : InMux
    port map (
            O => \N__4606\,
            I => \N__4603\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4603\,
            I => \N__4600\
        );

    \I__535\ : Span4Mux_h
    port map (
            O => \N__4600\,
            I => \N__4597\
        );

    \I__534\ : Odrv4
    port map (
            O => \N__4597\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__533\ : CascadeMux
    port map (
            O => \N__4594\,
            I => \U712_CHIP_RAM.N_354_cascade_\
        );

    \I__532\ : CascadeMux
    port map (
            O => \N__4591\,
            I => \U712_CHIP_RAM.N_414_cascade_\
        );

    \I__531\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4580\
        );

    \I__530\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4580\
        );

    \I__529\ : InMux
    port map (
            O => \N__4586\,
            I => \N__4575\
        );

    \I__528\ : InMux
    port map (
            O => \N__4585\,
            I => \N__4575\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4580\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4575\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__525\ : InMux
    port map (
            O => \N__4570\,
            I => \N__4567\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4567\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_3\
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__4564\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_2_cascade_\
        );

    \I__522\ : InMux
    port map (
            O => \N__4561\,
            I => \N__4558\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4558\,
            I => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\
        );

    \I__520\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4548\
        );

    \I__519\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4548\
        );

    \I__518\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4545\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4548\,
            I => \CPU_TACKm\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4545\,
            I => \CPU_TACKm\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__4540\,
            I => \N__4537\
        );

    \I__514\ : InMux
    port map (
            O => \N__4537\,
            I => \N__4530\
        );

    \I__513\ : InMux
    port map (
            O => \N__4536\,
            I => \N__4530\
        );

    \I__512\ : InMux
    port map (
            O => \N__4535\,
            I => \N__4527\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4530\,
            I => \REG_TACK\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__4527\,
            I => \REG_TACK\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__4522\,
            I => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\
        );

    \I__508\ : CascadeMux
    port map (
            O => \N__4519\,
            I => \U712_CYCLE_TERM.N_239_i_0_en_cascade_\
        );

    \I__507\ : InMux
    port map (
            O => \N__4516\,
            I => \N__4513\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4513\,
            I => \N__4510\
        );

    \I__505\ : Odrv12
    port map (
            O => \N__4510\,
            I => \TACK_EN_i_ess\
        );

    \I__504\ : IoInMux
    port map (
            O => \N__4507\,
            I => \N__4504\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4504\,
            I => \N__4501\
        );

    \I__502\ : Span12Mux_s5_h
    port map (
            O => \N__4501\,
            I => \N__4498\
        );

    \I__501\ : Span12Mux_v
    port map (
            O => \N__4498\,
            I => \N__4494\
        );

    \I__500\ : InMux
    port map (
            O => \N__4497\,
            I => \N__4491\
        );

    \I__499\ : Odrv12
    port map (
            O => \N__4494\,
            I => \TACK_OUTn\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4491\,
            I => \TACK_OUTn\
        );

    \I__497\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4483\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__4483\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__495\ : IoInMux
    port map (
            O => \N__4480\,
            I => \N__4477\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4477\,
            I => \N__4474\
        );

    \I__493\ : Span4Mux_s2_v
    port map (
            O => \N__4474\,
            I => \N__4471\
        );

    \I__492\ : Span4Mux_v
    port map (
            O => \N__4471\,
            I => \N__4468\
        );

    \I__491\ : Span4Mux_v
    port map (
            O => \N__4468\,
            I => \N__4465\
        );

    \I__490\ : Span4Mux_v
    port map (
            O => \N__4465\,
            I => \N__4461\
        );

    \I__489\ : InMux
    port map (
            O => \N__4464\,
            I => \N__4458\
        );

    \I__488\ : Odrv4
    port map (
            O => \N__4461\,
            I => \DBDIR_c\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4458\,
            I => \DBDIR_c\
        );

    \I__486\ : CascadeMux
    port map (
            O => \N__4453\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0_a3_0_0_cascade_\
        );

    \I__485\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4447\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4447\,
            I => \U712_CHIP_RAM.N_345\
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__4444\,
            I => \N__4441\
        );

    \I__482\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4438\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4438\,
            I => \U712_CHIP_RAM.N_71_i\
        );

    \I__480\ : CascadeMux
    port map (
            O => \N__4435\,
            I => \U712_CHIP_RAM.N_71_i_cascade_\
        );

    \I__479\ : InMux
    port map (
            O => \N__4432\,
            I => \N__4429\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4429\,
            I => \U712_CHIP_RAM.N_49\
        );

    \I__477\ : CascadeMux
    port map (
            O => \N__4426\,
            I => \U712_CHIP_RAM.N_361_cascade_\
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__4423\,
            I => \U712_CHIP_RAM.N_344_cascade_\
        );

    \I__475\ : InMux
    port map (
            O => \N__4420\,
            I => \N__4417\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4417\,
            I => \N__4414\
        );

    \I__473\ : Span12Mux_v
    port map (
            O => \N__4414\,
            I => \N__4411\
        );

    \I__472\ : Odrv12
    port map (
            O => \N__4411\,
            I => \A_c_9\
        );

    \I__471\ : InMux
    port map (
            O => \N__4408\,
            I => \N__4405\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4405\,
            I => \N__4402\
        );

    \I__469\ : Sp12to4
    port map (
            O => \N__4402\,
            I => \N__4399\
        );

    \I__468\ : Span12Mux_v
    port map (
            O => \N__4399\,
            I => \N__4396\
        );

    \I__467\ : Odrv12
    port map (
            O => \N__4396\,
            I => \A_c_2\
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__4393\,
            I => \U712_CHIP_RAM.N_253_cascade_\
        );

    \I__465\ : InMux
    port map (
            O => \N__4390\,
            I => \N__4387\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4387\,
            I => \N__4383\
        );

    \I__463\ : InMux
    port map (
            O => \N__4386\,
            I => \N__4380\
        );

    \I__462\ : Odrv4
    port map (
            O => \N__4383\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4380\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__4375\,
            I => \N__4372\
        );

    \I__459\ : InMux
    port map (
            O => \N__4372\,
            I => \N__4369\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4369\,
            I => \N__4366\
        );

    \I__457\ : Odrv4
    port map (
            O => \N__4366\,
            I => \U712_CHIP_RAM.N_344\
        );

    \I__456\ : IoInMux
    port map (
            O => \N__4363\,
            I => \N__4360\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4360\,
            I => \N__4357\
        );

    \I__454\ : Span12Mux_s5_v
    port map (
            O => \N__4357\,
            I => \N__4354\
        );

    \I__453\ : Span12Mux_v
    port map (
            O => \N__4354\,
            I => \N__4350\
        );

    \I__452\ : InMux
    port map (
            O => \N__4353\,
            I => \N__4347\
        );

    \I__451\ : Odrv12
    port map (
            O => \N__4350\,
            I => \LATCH_CLK_c\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4347\,
            I => \LATCH_CLK_c\
        );

    \I__449\ : InMux
    port map (
            O => \N__4342\,
            I => \N__4339\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4339\,
            I => \N__4336\
        );

    \I__447\ : Span4Mux_v
    port map (
            O => \N__4336\,
            I => \N__4333\
        );

    \I__446\ : Sp12to4
    port map (
            O => \N__4333\,
            I => \N__4330\
        );

    \I__445\ : Span12Mux_s10_h
    port map (
            O => \N__4330\,
            I => \N__4327\
        );

    \I__444\ : Span12Mux_v
    port map (
            O => \N__4327\,
            I => \N__4324\
        );

    \I__443\ : Odrv12
    port map (
            O => \N__4324\,
            I => \RAMSPACEn_c\
        );

    \I__442\ : CascadeMux
    port map (
            O => \N__4321\,
            I => \U712_CHIP_RAM.N_318_cascade_\
        );

    \I__441\ : InMux
    port map (
            O => \N__4318\,
            I => \N__4315\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4315\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__4312\,
            I => \U712_CHIP_RAM.BANK0_RNOZ0Z_0_cascade_\
        );

    \I__438\ : IoInMux
    port map (
            O => \N__4309\,
            I => \N__4306\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__4306\,
            I => \N__4303\
        );

    \I__436\ : Span4Mux_s1_v
    port map (
            O => \N__4303\,
            I => \N__4300\
        );

    \I__435\ : Span4Mux_v
    port map (
            O => \N__4300\,
            I => \N__4297\
        );

    \I__434\ : Span4Mux_v
    port map (
            O => \N__4297\,
            I => \N__4294\
        );

    \I__433\ : Span4Mux_h
    port map (
            O => \N__4294\,
            I => \N__4290\
        );

    \I__432\ : InMux
    port map (
            O => \N__4293\,
            I => \N__4287\
        );

    \I__431\ : Odrv4
    port map (
            O => \N__4290\,
            I => \BANK0_c\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__4287\,
            I => \BANK0_c\
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__4282\,
            I => \N__4279\
        );

    \I__428\ : InMux
    port map (
            O => \N__4279\,
            I => \N__4276\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__4276\,
            I => \N__4273\
        );

    \I__426\ : Odrv4
    port map (
            O => \N__4273\,
            I => \U712_CHIP_RAM.BANK0_RNOZ0Z_2\
        );

    \I__425\ : InMux
    port map (
            O => \N__4270\,
            I => \N__4267\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__4267\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\
        );

    \I__423\ : InMux
    port map (
            O => \N__4264\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__4261\,
            I => \N__4257\
        );

    \I__421\ : InMux
    port map (
            O => \N__4260\,
            I => \N__4254\
        );

    \I__420\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4251\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__4254\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__4251\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__417\ : InMux
    port map (
            O => \N__4246\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__416\ : InMux
    port map (
            O => \N__4243\,
            I => \N__4239\
        );

    \I__415\ : InMux
    port map (
            O => \N__4242\,
            I => \N__4236\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__4239\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__4236\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__412\ : InMux
    port map (
            O => \N__4231\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__411\ : InMux
    port map (
            O => \N__4228\,
            I => \N__4224\
        );

    \I__410\ : InMux
    port map (
            O => \N__4227\,
            I => \N__4221\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__4224\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__4221\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__407\ : InMux
    port map (
            O => \N__4216\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__406\ : InMux
    port map (
            O => \N__4213\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__405\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4206\
        );

    \I__404\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4203\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__4206\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__4203\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__401\ : IoInMux
    port map (
            O => \N__4198\,
            I => \N__4195\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__4195\,
            I => \N__4192\
        );

    \I__399\ : Span4Mux_s2_v
    port map (
            O => \N__4192\,
            I => \N__4189\
        );

    \I__398\ : Span4Mux_h
    port map (
            O => \N__4189\,
            I => \N__4186\
        );

    \I__397\ : Span4Mux_v
    port map (
            O => \N__4186\,
            I => \N__4183\
        );

    \I__396\ : Sp12to4
    port map (
            O => \N__4183\,
            I => \N__4180\
        );

    \I__395\ : Span12Mux_h
    port map (
            O => \N__4180\,
            I => \N__4176\
        );

    \I__394\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4173\
        );

    \I__393\ : Odrv12
    port map (
            O => \N__4176\,
            I => \ASn_c\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__4173\,
            I => \ASn_c\
        );

    \I__391\ : CascadeMux
    port map (
            O => \N__4168\,
            I => \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0_cascade_\
        );

    \I__390\ : IoInMux
    port map (
            O => \N__4165\,
            I => \N__4162\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__4162\,
            I => \N__4159\
        );

    \I__388\ : Odrv12
    port map (
            O => \N__4159\,
            I => \DBRn_c_i_0\
        );

    \I__387\ : IoInMux
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__4153\,
            I => \N__4150\
        );

    \I__385\ : Span4Mux_s2_h
    port map (
            O => \N__4150\,
            I => \N__4147\
        );

    \I__384\ : Span4Mux_h
    port map (
            O => \N__4147\,
            I => \N__4144\
        );

    \I__383\ : Sp12to4
    port map (
            O => \N__4144\,
            I => \N__4141\
        );

    \I__382\ : Odrv12
    port map (
            O => \N__4141\,
            I => \N_969_i\
        );

    \I__381\ : CEMux
    port map (
            O => \N__4138\,
            I => \N__4135\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__4135\,
            I => \N__4132\
        );

    \I__379\ : Span4Mux_h
    port map (
            O => \N__4132\,
            I => \N__4129\
        );

    \I__378\ : Odrv4
    port map (
            O => \N__4129\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0\
        );

    \I__377\ : InMux
    port map (
            O => \N__4126\,
            I => \N__4122\
        );

    \I__376\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4119\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__4122\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__4119\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__373\ : InMux
    port map (
            O => \N__4114\,
            I => \bfn_7_9_0_\
        );

    \I__372\ : InMux
    port map (
            O => \N__4111\,
            I => \N__4107\
        );

    \I__371\ : InMux
    port map (
            O => \N__4110\,
            I => \N__4104\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__4107\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__4104\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__368\ : InMux
    port map (
            O => \N__4099\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__367\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4092\
        );

    \I__366\ : InMux
    port map (
            O => \N__4095\,
            I => \N__4089\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__4092\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__4089\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__363\ : InMux
    port map (
            O => \N__4084\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__362\ : IoInMux
    port map (
            O => \N__4081\,
            I => \N__4078\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__4078\,
            I => \N__4075\
        );

    \I__360\ : IoSpan4Mux
    port map (
            O => \N__4075\,
            I => \N__4072\
        );

    \I__359\ : Span4Mux_s3_v
    port map (
            O => \N__4072\,
            I => \N__4069\
        );

    \I__358\ : Odrv4
    port map (
            O => \N__4069\,
            I => \CLK80_PLL_i_i\
        );

    \I__357\ : IoInMux
    port map (
            O => \N__4066\,
            I => \N__4063\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__4063\,
            I => \N__4060\
        );

    \I__355\ : Span4Mux_s0_v
    port map (
            O => \N__4060\,
            I => \N__4057\
        );

    \I__354\ : Span4Mux_v
    port map (
            O => \N__4057\,
            I => \N__4054\
        );

    \I__353\ : Sp12to4
    port map (
            O => \N__4054\,
            I => \N__4051\
        );

    \I__352\ : Span12Mux_h
    port map (
            O => \N__4051\,
            I => \N__4048\
        );

    \I__351\ : Span12Mux_v
    port map (
            O => \N__4048\,
            I => \N__4045\
        );

    \I__350\ : Odrv12
    port map (
            O => \N__4045\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__7292\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__7293\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__7286\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__7291\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__7284\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__7285\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__7290\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__7283\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_7_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_9_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9124\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5238\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4165\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6973\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8794\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10180\,
            in2 => \_gnd_net_\,
            in3 => \N__9436\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4516\,
            lcout => \N_969_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5158\,
            in1 => \N__7433\,
            in2 => \_gnd_net_\,
            in3 => \N__6002\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8776\,
            ce => \N__4138\,
            sr => \N__10150\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4209\,
            in1 => \N__4227\,
            in2 => \_gnd_net_\,
            in3 => \N__4242\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10178\,
            in2 => \_gnd_net_\,
            in3 => \N__4386\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__4095\,
            in1 => \N__4125\,
            in2 => \N__4261\,
            in3 => \N__4110\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4126\,
            in2 => \_gnd_net_\,
            in3 => \N__4114\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_7_9_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__7294\,
            ce => 'H',
            sr => \N__5563\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4111\,
            in2 => \_gnd_net_\,
            in3 => \N__4099\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__7294\,
            ce => 'H',
            sr => \N__5563\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4096\,
            in2 => \_gnd_net_\,
            in3 => \N__4084\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__7294\,
            ce => 'H',
            sr => \N__5563\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4635\,
            in2 => \_gnd_net_\,
            in3 => \N__4264\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__7294\,
            ce => 'H',
            sr => \N__5563\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4260\,
            in2 => \_gnd_net_\,
            in3 => \N__4246\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__7294\,
            ce => 'H',
            sr => \N__5563\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4243\,
            in2 => \_gnd_net_\,
            in3 => \N__4231\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__7294\,
            ce => 'H',
            sr => \N__5563\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4228\,
            in2 => \_gnd_net_\,
            in3 => \N__4216\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__7294\,
            ce => 'H',
            sr => \N__5563\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4210\,
            in2 => \_gnd_net_\,
            in3 => \N__4213\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7294\,
            ce => 'H',
            sr => \N__5563\
        );

    \U712_REG_SM.ASn_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__4179\,
            in1 => \N__7771\,
            in2 => \N__7819\,
            in3 => \N__7246\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8788\,
            ce => 'H',
            sr => \N__10126\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4318\,
            in2 => \_gnd_net_\,
            in3 => \N__5643\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011101010"
        )
    port map (
            in0 => \N__5144\,
            in1 => \N__9304\,
            in2 => \N__4168\,
            in3 => \N__5009\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9726\,
            in2 => \_gnd_net_\,
            in3 => \N__5503\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_318_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__4342\,
            in1 => \N__7183\,
            in2 => \N__4321\,
            in3 => \N__9303\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIRILU_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4586\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5142\,
            lcout => \U712_CHIP_RAM.N_366\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5644\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9302\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8764\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIR9VE1_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4585\,
            in1 => \N__5143\,
            in2 => \N__5476\,
            in3 => \N__5502\,
            lcout => \U712_CHIP_RAM.N_413\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100100010"
        )
    port map (
            in0 => \N__4270\,
            in1 => \N__4666\,
            in2 => \N__4282\,
            in3 => \N__9412\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.BANK0_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__4293\,
            in1 => \N__6243\,
            in2 => \N__4312\,
            in3 => \N__5086\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8772\,
            ce => 'H',
            sr => \N__10141\
        );

    \U712_CHIP_RAM.BANK0_RNO_2_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__5146\,
            in1 => \_gnd_net_\,
            in2 => \N__5896\,
            in3 => \N__5976\,
            lcout => \U712_CHIP_RAM.BANK0_RNOZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVLD65_1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5977\,
            in1 => \N__5891\,
            in2 => \_gnd_net_\,
            in3 => \N__5912\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_2_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7506\,
            in1 => \N__6446\,
            in2 => \N__7648\,
            in3 => \N__6298\,
            lcout => \U712_CHIP_RAM.N_357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNIGMCR2_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6447\,
            in1 => \N__5005\,
            in2 => \N__6325\,
            in3 => \N__7612\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNISBTD7_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__5145\,
            in1 => \N__7416\,
            in2 => \N__4426\,
            in3 => \N__5975\,
            lcout => \U712_CHIP_RAM.N_344\,
            ltout => \U712_CHIP_RAM.N_344_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIT2EQB_0_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__6448\,
            in1 => \N__6326\,
            in2 => \N__4423\,
            in3 => \N__6022\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI71B91_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111001010100"
        )
    port map (
            in0 => \N__6439\,
            in1 => \N__7507\,
            in2 => \N__10974\,
            in3 => \N__5004\,
            lcout => \U712_CHIP_RAM.N_217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5159\,
            in1 => \N__7440\,
            in2 => \_gnd_net_\,
            in3 => \N__5998\,
            lcout => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4420\,
            in1 => \N__4408\,
            in2 => \_gnd_net_\,
            in3 => \N__9528\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__6440\,
            in1 => \N__7508\,
            in2 => \_gnd_net_\,
            in3 => \N__6146\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_253_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110101111"
        )
    port map (
            in0 => \N__7646\,
            in1 => \N__5889\,
            in2 => \N__4393\,
            in3 => \N__10959\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011101110"
        )
    port map (
            in0 => \N__5044\,
            in1 => \N__4390\,
            in2 => \N__4444\,
            in3 => \N__9796\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8780\,
            ce => 'H',
            sr => \N__10134\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010011111110"
        )
    port map (
            in0 => \N__4450\,
            in1 => \N__4353\,
            in2 => \N__4375\,
            in3 => \N__4432\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8780\,
            ce => 'H',
            sr => \N__10134\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110100010"
        )
    port map (
            in0 => \N__4497\,
            in1 => \N__5310\,
            in2 => \N__9391\,
            in3 => \N__4957\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8780\,
            ce => 'H',
            sr => \N__10134\
        );

    \U712_CHIP_RAM.DBDIR_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__5202\,
            in1 => \N__4464\,
            in2 => \_gnd_net_\,
            in3 => \N__4486\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8780\,
            ce => 'H',
            sr => \N__10134\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5881\,
            in2 => \_gnd_net_\,
            in3 => \N__6142\,
            lcout => \U712_CHIP_RAM.N_274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_3_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7439\,
            in1 => \N__7541\,
            in2 => \N__10982\,
            in3 => \N__7661\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__6334\,
            in1 => \_gnd_net_\,
            in2 => \N__4453\,
            in3 => \N__6452\,
            lcout => \U712_CHIP_RAM.N_345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__5022\,
            in1 => \N__5045\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101101"
        )
    port map (
            in0 => \N__7662\,
            in1 => \N__10973\,
            in2 => \N__7549\,
            in3 => \N__6453\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5888\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6010\,
            lcout => \U712_CHIP_RAM.N_71_i\,
            ltout => \U712_CHIP_RAM.N_71_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111111"
        )
    port map (
            in0 => \N__5068\,
            in1 => \N__5160\,
            in2 => \N__4435\,
            in3 => \N__5021\,
            lcout => \U712_CHIP_RAM.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__4978\,
            in1 => \N__7663\,
            in2 => \N__6340\,
            in3 => \N__7545\,
            lcout => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111011111111"
        )
    port map (
            in0 => \N__6335\,
            in1 => \N__5890\,
            in2 => \N__6454\,
            in3 => \N__6151\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__4555\,
            in1 => \N__4570\,
            in2 => \N__4564\,
            in3 => \N__4561\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8785\,
            ce => 'H',
            sr => \N__10119\
        );

    \U712_REG_SM.REG_TACK_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__7734\,
            in1 => \N__5335\,
            in2 => \N__4540\,
            in3 => \N__4972\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8785\,
            ce => 'H',
            sr => \N__10119\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010101"
        )
    port map (
            in0 => \N__5302\,
            in1 => \N__4536\,
            in2 => \N__5269\,
            in3 => \N__4554\,
            lcout => \U712_CYCLE_TERM.N_340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9243\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4953\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4553\,
            in2 => \_gnd_net_\,
            in3 => \N__4535\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__9242\,
            in1 => \N__5280\,
            in2 => \N__4522\,
            in3 => \N__5263\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_239_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10176\,
            in1 => \_gnd_net_\,
            in2 => \N__4519\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.N_239_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__9244\,
            in1 => \N__5267\,
            in2 => \_gnd_net_\,
            in3 => \N__5323\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8790\,
            ce => \N__4699\,
            sr => \N__10108\
        );

    \U712_CHIP_RAM.BANK0_RNO_1_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4684\,
            in2 => \_gnd_net_\,
            in3 => \N__10483\,
            lcout => \U712_CHIP_RAM.BANK0_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__9722\,
            in1 => \N__10935\,
            in2 => \_gnd_net_\,
            in3 => \N__7530\,
            lcout => \U712_CHIP_RAM.CLK_EN_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIM0601_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__5504\,
            in1 => \N__9299\,
            in2 => \_gnd_net_\,
            in3 => \N__5474\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a2_2_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a3_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9723\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10009\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010001100"
        )
    port map (
            in0 => \N__4639\,
            in1 => \N__9300\,
            in2 => \N__4621\,
            in3 => \N__4606\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8759\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIEH9V_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5475\,
            in1 => \N__4587\,
            in2 => \_gnd_net_\,
            in3 => \N__5505\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_354_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIQ6QH5_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__7441\,
            in1 => \N__5148\,
            in2 => \N__4594\,
            in3 => \N__5991\,
            lcout => \U712_CHIP_RAM.N_414\,
            ltout => \U712_CHIP_RAM.N_414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4591\,
            in3 => \N__10179\,
            lcout => \U712_CHIP_RAM.N_414_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4588\,
            in1 => \N__9301\,
            in2 => \N__6135\,
            in3 => \N__5147\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6419\,
            in2 => \_gnd_net_\,
            in3 => \N__4723\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5869\,
            in2 => \_gnd_net_\,
            in3 => \N__4720\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6215\,
            in1 => \N__7532\,
            in2 => \_gnd_net_\,
            in3 => \N__4717\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \N__8765\,
            ce => \N__6173\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6203\,
            in1 => \N__7647\,
            in2 => \_gnd_net_\,
            in3 => \N__4714\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__8765\,
            ce => \N__6173\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6216\,
            in1 => \N__4768\,
            in2 => \_gnd_net_\,
            in3 => \N__4711\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__8765\,
            ce => \N__6173\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6204\,
            in1 => \N__4795\,
            in2 => \_gnd_net_\,
            in3 => \N__4708\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__8765\,
            ce => \N__6173\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6217\,
            in1 => \N__4807\,
            in2 => \_gnd_net_\,
            in3 => \N__4705\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__8765\,
            ce => \N__6173\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6205\,
            in1 => \N__4782\,
            in2 => \_gnd_net_\,
            in3 => \N__4702\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8765\,
            ce => \N__6173\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110111"
        )
    port map (
            in0 => \N__7533\,
            in1 => \N__6424\,
            in2 => \N__7651\,
            in3 => \N__6309\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_0_a2_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110100000001"
        )
    port map (
            in0 => \N__4849\,
            in1 => \N__5424\,
            in2 => \N__4840\,
            in3 => \N__4818\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8773\,
            ce => 'H',
            sr => \N__10135\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4806\,
            in1 => \N__4794\,
            in2 => \N__4783\,
            in3 => \N__4767\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4756\,
            in3 => \N__9266\,
            lcout => \U712_CHIP_RAM.N_230\,
            ltout => \U712_CHIP_RAM.N_230_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5368\,
            in1 => \N__7645\,
            in2 => \N__4753\,
            in3 => \N__7531\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__4750\,
            in1 => \N__5359\,
            in2 => \N__4741\,
            in3 => \N__6012\,
            lcout => \U712_CHIP_RAM.N_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAGAE4_3_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4738\,
            in1 => \N__7434\,
            in2 => \N__7650\,
            in3 => \N__6308\,
            lcout => \U712_CHIP_RAM.N_282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__4865\,
            in1 => \N__4732\,
            in2 => \_gnd_net_\,
            in3 => \N__9525\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIEMD13_3_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100000001"
        )
    port map (
            in0 => \N__5343\,
            in1 => \N__5420\,
            in2 => \N__7668\,
            in3 => \N__7438\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_113_tz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3T4K7_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__6046\,
            in1 => \N__5353\,
            in2 => \N__4726\,
            in3 => \N__4897\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3T4KZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNILMT6D_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5482\,
            in1 => \N__5397\,
            in2 => \N__4927\,
            in3 => \N__6011\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001110"
        )
    port map (
            in0 => \N__4924\,
            in1 => \N__4909\,
            in2 => \N__4918\,
            in3 => \N__7953\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__7548\,
            in1 => \N__7659\,
            in2 => \_gnd_net_\,
            in3 => \N__5344\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000110010"
        )
    port map (
            in0 => \N__4873\,
            in1 => \N__4866\,
            in2 => \N__4915\,
            in3 => \N__8136\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000110000"
        )
    port map (
            in0 => \N__5883\,
            in1 => \N__6433\,
            in2 => \N__6150\,
            in3 => \N__10976\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_284_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__6133\,
            in1 => \N__4903\,
            in2 => \N__4912\,
            in3 => \N__4896\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7652\,
            in2 => \_gnd_net_\,
            in3 => \N__7540\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRTZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITVCO3_1_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4895\,
            in2 => \N__4876\,
            in3 => \N__5884\,
            lcout => \U712_CHIP_RAM.N_271\,
            ltout => \U712_CHIP_RAM.N_271_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000110010"
        )
    port map (
            in0 => \N__5062\,
            in1 => \N__4867\,
            in2 => \N__4852\,
            in3 => \N__8072\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8781\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_2_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6432\,
            in1 => \N__5882\,
            in2 => \N__7667\,
            in3 => \N__6333\,
            lcout => \U712_CHIP_RAM.N_347\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011100110"
        )
    port map (
            in0 => \N__7546\,
            in1 => \N__6434\,
            in2 => \N__7669\,
            in3 => \N__6134\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5046\,
            in2 => \_gnd_net_\,
            in3 => \N__5023\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4965\,
            in2 => \_gnd_net_\,
            in3 => \N__4949\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__9380\,
            in1 => \N__9193\,
            in2 => \_gnd_net_\,
            in3 => \N__5309\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8784\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001000000000"
        )
    port map (
            in0 => \N__10975\,
            in1 => \N__6435\,
            in2 => \N__5895\,
            in3 => \N__9709\,
            lcout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6727\,
            in1 => \N__6898\,
            in2 => \_gnd_net_\,
            in3 => \N__6923\,
            lcout => \U712_REG_SM.N_304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__9194\,
            in1 => \N__4966\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8784\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__4933\,
            in1 => \N__9192\,
            in2 => \N__9384\,
            in3 => \N__5268\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8784\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__7759\,
            in1 => \N__11116\,
            in2 => \N__6838\,
            in3 => \N__7802\,
            lcout => \U712_REG_SM.N_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111100001000"
        )
    port map (
            in0 => \N__5329\,
            in1 => \N__5322\,
            in2 => \N__5311\,
            in3 => \N__5281\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8786\,
            ce => 'H',
            sr => \N__10109\
        );

    \U712_REG_SM.C1_SYNC_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5242\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8786\,
            ce => 'H',
            sr => \N__10109\
        );

    \U712_BYTE_ENABLE.LLBE_i_o3_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010111011"
        )
    port map (
            in0 => \N__8443\,
            in1 => \N__8506\,
            in2 => \N__8260\,
            in3 => \N__8363\,
            lcout => \U712_BYTE_ENABLE.N_242\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__11122\,
            in1 => \N__5203\,
            in2 => \_gnd_net_\,
            in3 => \N__5161\,
            lcout => \WRITE_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8756\,
            ce => \N__5101\,
            sr => \N__10139\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_2_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7608\,
            in2 => \_gnd_net_\,
            in3 => \N__7505\,
            lcout => \U712_CHIP_RAM.N_363\,
            ltout => \U712_CHIP_RAM.N_363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5573\,
            in1 => \N__6418\,
            in2 => \N__5089\,
            in3 => \N__6310\,
            lcout => \U712_CHIP_RAM.N_292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI0Q6U4_3_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9298\,
            in2 => \_gnd_net_\,
            in3 => \N__5085\,
            lcout => \U712_CHIP_RAM.N_236\,
            ltout => \U712_CHIP_RAM.N_236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIUJS3D_0_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__5575\,
            in1 => \N__5074\,
            in2 => \N__5431\,
            in3 => \N__6004\,
            lcout => \U712_CHIP_RAM.N_48_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI27TJ3_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6311\,
            in1 => \N__5574\,
            in2 => \_gnd_net_\,
            in3 => \N__6042\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__5428\,
            in1 => \_gnd_net_\,
            in2 => \N__5404\,
            in3 => \N__6005\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_i_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIGGM16_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__6003\,
            in1 => \N__5401\,
            in2 => \N__7432\,
            in3 => \N__5380\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__9297\,
            in1 => \N__5374\,
            in2 => \_gnd_net_\,
            in3 => \N__6125\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8760\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_5_1_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6100\,
            in1 => \N__6416\,
            in2 => \_gnd_net_\,
            in3 => \N__5851\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_4_1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011000010100"
        )
    port map (
            in0 => \N__7516\,
            in1 => \N__5831\,
            in2 => \N__7660\,
            in3 => \N__6101\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_252_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__9259\,
            in1 => \N__6417\,
            in2 => \N__5362\,
            in3 => \N__6324\,
            lcout => \U712_CHIP_RAM.N_286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMT791_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6415\,
            in1 => \N__5830\,
            in2 => \_gnd_net_\,
            in3 => \N__6099\,
            lcout => \U712_CHIP_RAM.N_267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7515\,
            in2 => \_gnd_net_\,
            in3 => \N__6414\,
            lcout => \U712_CHIP_RAM.N_225_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__5596\,
            in1 => \N__5590\,
            in2 => \N__5584\,
            in3 => \N__6206\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8766\,
            ce => \N__6177\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5829\,
            in2 => \_gnd_net_\,
            in3 => \N__6098\,
            lcout => \U712_CHIP_RAM.N_234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100110001"
        )
    port map (
            in0 => \N__7942\,
            in1 => \N__8065\,
            in2 => \N__9527\,
            in3 => \N__8125\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8064\,
            in1 => \N__8124\,
            in2 => \N__9526\,
            in3 => \N__7941\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__5554\,
            in1 => \N__9018\,
            in2 => \N__10750\,
            in3 => \N__9710\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8774\,
            ce => \N__8668\,
            sr => \N__10120\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIHHIB1_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__5461\,
            in1 => \N__9254\,
            in2 => \N__5515\,
            in3 => \N__6129\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5442\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8778\,
            ce => 'H',
            sr => \N__10113\
        );

    \DBR_SYNC_0_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6508\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8778\,
            ce => 'H',
            sr => \N__10113\
        );

    \U712_REG_SM.C1_SYNC_RNIS63V_1_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__6579\,
            in1 => \N__5462\,
            in2 => \N__5443\,
            in3 => \N__6549\,
            lcout => OPEN,
            ltout => \U712_REG_SM.STATE_COUNT_srsts_i_i_o2_0_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI35EO1_1_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__6770\,
            in1 => \_gnd_net_\,
            in2 => \N__5602\,
            in3 => \N__6799\,
            lcout => \U712_REG_SM.N_266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_1_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6550\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8778\,
            ce => 'H',
            sr => \N__10113\
        );

    \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__6769\,
            in1 => \N__6578\,
            in2 => \N__6555\,
            in3 => \N__6798\,
            lcout => \U712_REG_SM.N_220\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6507\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6807\,
            in1 => \N__6577\,
            in2 => \N__6551\,
            in3 => \N__6772\,
            lcout => \U712_REG_SM.N_367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000011000000"
        )
    port map (
            in0 => \N__6900\,
            in1 => \N__9190\,
            in2 => \N__6859\,
            in3 => \N__7242\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_4_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__6834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6924\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_272_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__9191\,
            in1 => \N__7818\,
            in2 => \N__5599\,
            in3 => \N__7760\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100011101"
        )
    port map (
            in0 => \N__6731\,
            in1 => \N__7705\,
            in2 => \N__7123\,
            in3 => \N__6925\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_270_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__7306\,
            in1 => \N__9189\,
            in2 => \N__5773\,
            in3 => \N__6742\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8782\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_202_i_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__5611\,
            in1 => \N__5718\,
            in2 => \N__11059\,
            in3 => \N__9731\,
            lcout => \N_202_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_188_i_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100010101"
        )
    port map (
            in0 => \N__5683\,
            in1 => \N__5746\,
            in2 => \N__9733\,
            in3 => \N__10885\,
            lcout => \N_188_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_203_i_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__10886\,
            in1 => \N__5719\,
            in2 => \N__5626\,
            in3 => \N__9732\,
            lcout => \N_203_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_186_i_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__5617\,
            in1 => \N__5682\,
            in2 => \N__11058\,
            in3 => \N__9727\,
            lcout => \N_186_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__10897\,
            in1 => \N__9255\,
            in2 => \_gnd_net_\,
            in3 => \N__11051\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_i_o3_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010001011111"
        )
    port map (
            in0 => \N__8442\,
            in1 => \N__8263\,
            in2 => \N__8507\,
            in3 => \N__8373\,
            lcout => \U712_BYTE_ENABLE.N_243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LMBE_i_o3_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111101101"
        )
    port map (
            in0 => \N__8496\,
            in1 => \N__8441\,
            in2 => \N__8374\,
            in3 => \N__8262\,
            lcout => \U712_BYTE_ENABLE.N_244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_i_o3_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100011111"
        )
    port map (
            in0 => \N__8440\,
            in1 => \N__8261\,
            in2 => \N__8364\,
            in3 => \N__8495\,
            lcout => \U712_BYTE_ENABLE.N_245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__9275\,
            in1 => \N__6492\,
            in2 => \_gnd_net_\,
            in3 => \N__7212\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10240\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DMA_LATCH_EN_0_a3_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__10893\,
            in1 => \N__11050\,
            in2 => \_gnd_net_\,
            in3 => \N__10989\,
            lcout => \DMA_LATCH_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6423\,
            in1 => \N__7363\,
            in2 => \_gnd_net_\,
            in3 => \N__6339\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_320_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5925\,
            in1 => \N__7412\,
            in2 => \N__6253\,
            in3 => \N__6006\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10177\,
            in1 => \_gnd_net_\,
            in2 => \N__6250\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__9276\,
            in1 => \N__6247\,
            in2 => \N__6229\,
            in3 => \N__6207\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8757\,
            ce => \N__6178\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_1_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5825\,
            in2 => \_gnd_net_\,
            in3 => \N__6097\,
            lcout => \U712_CHIP_RAM.N_358\,
            ltout => \U712_CHIP_RAM.N_358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIQIR12_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6041\,
            in2 => \N__6025\,
            in3 => \N__10926\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6013\,
            in1 => \N__5926\,
            in2 => \_gnd_net_\,
            in3 => \N__5852\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8761\,
            ce => \N__5779\,
            sr => \N__10121\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6697\,
            in1 => \N__6679\,
            in2 => \_gnd_net_\,
            in3 => \N__9556\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9557\,
            in1 => \N__9673\,
            in2 => \N__6661\,
            in3 => \N__9859\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6658\,
            in1 => \N__6640\,
            in2 => \_gnd_net_\,
            in3 => \N__9555\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9554\,
            in1 => \N__6619\,
            in2 => \_gnd_net_\,
            in3 => \N__6598\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__6774\,
            in1 => \N__11120\,
            in2 => \_gnd_net_\,
            in3 => \N__7803\,
            lcout => \U712_REG_SM.DS_EN_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_3_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111101110"
        )
    port map (
            in0 => \N__6899\,
            in1 => \N__6800\,
            in2 => \_gnd_net_\,
            in3 => \N__6773\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_269_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_2_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110101"
        )
    port map (
            in0 => \N__6732\,
            in1 => \N__6580\,
            in2 => \N__6559\,
            in3 => \N__6556\,
            lcout => OPEN,
            ltout => \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100011"
        )
    port map (
            in0 => \N__8576\,
            in1 => \N__6517\,
            in2 => \N__6511\,
            in3 => \N__6931\,
            lcout => \DS_ENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8775\,
            ce => 'H',
            sr => \N__10110\
        );

    \U712_REG_SM.C3_SYNC_1_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6775\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8775\,
            ce => 'H',
            sr => \N__10110\
        );

    \U712_REG_SM.C3_SYNC_0_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6960\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8775\,
            ce => 'H',
            sr => \N__10110\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__7804\,
            in1 => \N__6897\,
            in2 => \N__6736\,
            in3 => \N__7305\,
            lcout => \U712_REG_SM.N_313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6725\,
            in1 => \N__6829\,
            in2 => \_gnd_net_\,
            in3 => \N__6895\,
            lcout => \U712_REG_SM.N_374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_RNO_0_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7801\,
            in2 => \_gnd_net_\,
            in3 => \N__7758\,
            lcout => \U712_REG_SM.ASn_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7118\,
            in2 => \_gnd_net_\,
            in3 => \N__6921\,
            lcout => \U712_REG_SM.N_226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__6833\,
            in1 => \N__6896\,
            in2 => \_gnd_net_\,
            in3 => \N__6922\,
            lcout => OPEN,
            ltout => \U712_REG_SM.STATE_COUNTc_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__9188\,
            in1 => \N__6901\,
            in2 => \N__6862\,
            in3 => \N__6852\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI7UAP_1_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6808\,
            in2 => \_gnd_net_\,
            in3 => \N__6771\,
            lcout => \U712_REG_SM.N_222\,
            ltout => \U712_REG_SM.N_222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6726\,
            in2 => \N__7309\,
            in3 => \N__7304\,
            lcout => \U712_REG_SM.N_241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110111110000"
        )
    port map (
            in0 => \N__7704\,
            in1 => \N__7716\,
            in2 => \N__7231\,
            in3 => \N__7202\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8783\,
            ce => 'H',
            sr => \N__10103\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001101"
        )
    port map (
            in0 => \N__7179\,
            in1 => \N__7122\,
            in2 => \N__7147\,
            in3 => \N__9998\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8783\,
            ce => 'H',
            sr => \N__10103\
        );

    \U712_BYTE_ENABLE.N_243_i_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010110000"
        )
    port map (
            in0 => \N__8428\,
            in1 => \N__8264\,
            in2 => \N__8359\,
            in3 => \N__8508\,
            lcout => \N_243_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7966\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8752\,
            ce => 'H',
            sr => \N__10133\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8148\,
            in1 => \N__9571\,
            in2 => \N__8083\,
            in3 => \N__7962\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8754\,
            ce => \N__8660\,
            sr => \N__10125\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8915\,
            in1 => \N__9847\,
            in2 => \N__8887\,
            in3 => \N__7687\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8754\,
            ce => \N__8660\,
            sr => \N__10125\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7009\,
            in1 => \N__6994\,
            in2 => \_gnd_net_\,
            in3 => \N__9583\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__9112\,
            in1 => \N__9585\,
            in2 => \N__7690\,
            in3 => \N__9677\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__9584\,
            in1 => \N__10576\,
            in2 => \N__9708\,
            in3 => \N__7681\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_2_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__10960\,
            in1 => \N__7649\,
            in2 => \N__7547\,
            in3 => \N__7408\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8917\,
            in1 => \N__9103\,
            in2 => \N__8883\,
            in3 => \N__7357\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8755\,
            ce => \N__8644\,
            sr => \N__10112\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011110000"
        )
    port map (
            in0 => \N__9663\,
            in1 => \N__10761\,
            in2 => \N__8885\,
            in3 => \N__9552\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7336\,
            in1 => \N__9662\,
            in2 => \_gnd_net_\,
            in3 => \N__10774\,
            lcout => \U712_CHIP_RAM.N_333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10175\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7321\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__9551\,
            in1 => \N__8138\,
            in2 => \_gnd_net_\,
            in3 => \N__7955\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => \U712_CHIP_RAM.CMA_5_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110101111"
        )
    port map (
            in0 => \N__9088\,
            in1 => \N__7915\,
            in2 => \N__7312\,
            in3 => \N__9672\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8137\,
            in2 => \_gnd_net_\,
            in3 => \N__7954\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011111111"
        )
    port map (
            in0 => \N__9664\,
            in1 => \N__10762\,
            in2 => \N__7918\,
            in3 => \N__9553\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__7914\,
            in1 => \N__9665\,
            in2 => \N__9017\,
            in3 => \N__9087\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__7891\,
            in1 => \N__9707\,
            in2 => \N__10693\,
            in3 => \N__9587\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7885\,
            in2 => \N__7879\,
            in3 => \N__7876\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8763\,
            ce => \N__8645\,
            sr => \N__10104\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9586\,
            in2 => \N__7858\,
            in3 => \N__8865\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7849\,
            in2 => \N__7843\,
            in3 => \N__7840\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8763\,
            ce => \N__8645\,
            sr => \N__10104\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__7817\,
            in1 => \N__7767\,
            in2 => \N__7735\,
            in3 => \N__7717\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8768\,
            ce => 'H',
            sr => \N__10102\
        );

    \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__8595\,
            in1 => \N__8362\,
            in2 => \_gnd_net_\,
            in3 => \N__8251\,
            lcout => \N_182\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__8361\,
            in1 => \N__8252\,
            in2 => \_gnd_net_\,
            in3 => \N__8596\,
            lcout => \N_184\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_245_i_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011001000"
        )
    port map (
            in0 => \N__8424\,
            in1 => \N__8518\,
            in2 => \N__8266\,
            in3 => \N__8343\,
            lcout => \N_245_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_242_i_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101000100"
        )
    port map (
            in0 => \N__8422\,
            in1 => \N__8516\,
            in2 => \N__8265\,
            in3 => \N__8339\,
            lcout => \N_242_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_244_i_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000010010"
        )
    port map (
            in0 => \N__8517\,
            in1 => \N__8423\,
            in2 => \N__8360\,
            in3 => \N__8256\,
            lcout => \N_244_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RASn_LC_13_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8152\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8750\,
            ce => 'H',
            sr => \N__10156\
        );

    \U712_CHIP_RAM.CRCSn_LC_13_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8079\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8751\,
            ce => 'H',
            sr => \N__10152\
        );

    \U712_CHIP_RAM.CASn_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9589\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8753\,
            ce => 'H',
            sr => \N__10142\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8002\,
            in1 => \N__7984\,
            in2 => \_gnd_net_\,
            in3 => \N__9572\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9573\,
            in1 => \N__9721\,
            in2 => \N__9073\,
            in3 => \N__9781\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__9720\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9574\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\,
            ltout => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__8886\,
            in1 => \N__9835\,
            in2 => \N__9070\,
            in3 => \N__9067\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8758\,
            ce => \N__8667\,
            sr => \N__10127\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__9040\,
            in1 => \N__9703\,
            in2 => \N__9019\,
            in3 => \N__10249\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8762\,
            ce => \N__8650\,
            sr => \N__10122\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__8872\,
            in1 => \N__8908\,
            in2 => \N__9943\,
            in3 => \N__8971\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8762\,
            ce => \N__8650\,
            sr => \N__10122\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8907\,
            in1 => \N__9094\,
            in2 => \N__8884\,
            in3 => \N__9442\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8762\,
            ce => \N__8650\,
            sr => \N__10122\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__8926\,
            in1 => \N__9725\,
            in2 => \N__9588\,
            in3 => \N__10492\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__8916\,
            in1 => \N__8873\,
            in2 => \N__8818\,
            in3 => \N__9949\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8767\,
            ce => \N__8646\,
            sr => \N__10114\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9769\,
            in1 => \N__9751\,
            in2 => \_gnd_net_\,
            in3 => \N__9575\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9724\,
            in1 => \N__9576\,
            in2 => \N__9445\,
            in3 => \N__9934\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_A20_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__9432\,
            in1 => \N__10457\,
            in2 => \N__10309\,
            in3 => \N__9405\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__10111\
        );

    \pll_RNI8MQ3_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9376\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9296\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9928\,
            in1 => \N__10418\,
            in2 => \_gnd_net_\,
            in3 => \N__10723\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__10214\,
            sr => \N__10136\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10414\,
            in1 => \N__9923\,
            in2 => \_gnd_net_\,
            in3 => \N__10737\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10238\,
            ce => \N__10212\,
            sr => \N__10128\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9924\,
            in1 => \N__10415\,
            in2 => \_gnd_net_\,
            in3 => \N__9888\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10238\,
            ce => \N__10212\,
            sr => \N__10128\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9889\,
            in1 => \N__10472\,
            in2 => \_gnd_net_\,
            in3 => \N__10815\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10238\,
            ce => \N__10212\,
            sr => \N__10128\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10816\,
            in1 => \N__10563\,
            in2 => \_gnd_net_\,
            in3 => \N__10416\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10238\,
            ce => \N__10212\,
            sr => \N__10128\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__10528\,
            in1 => \_gnd_net_\,
            in2 => \N__10567\,
            in3 => \N__10473\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10238\,
            ce => \N__10212\,
            sr => \N__10128\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10799\,
            in1 => \N__10470\,
            in2 => \_gnd_net_\,
            in3 => \N__9887\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__10210\,
            sr => \N__10123\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9922\,
            in1 => \N__10410\,
            in2 => \_gnd_net_\,
            in3 => \N__9886\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__10209\,
            sr => \N__10115\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10676\,
            in1 => \N__10479\,
            in2 => \_gnd_net_\,
            in3 => \N__10738\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10239\,
            ce => \N__10217\,
            sr => \N__10140\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9826\,
            in1 => \N__10478\,
            in2 => \_gnd_net_\,
            in3 => \N__10626\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10239\,
            ce => \N__10217\,
            sr => \N__10140\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10627\,
            in1 => \N__10468\,
            in2 => \_gnd_net_\,
            in3 => \N__9825\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10215\,
            sr => \N__10137\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10527\,
            in1 => \N__10469\,
            in2 => \_gnd_net_\,
            in3 => \N__10308\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10215\,
            sr => \N__10137\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10471\,
            in1 => \N__10562\,
            in2 => \_gnd_net_\,
            in3 => \N__10814\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10215\,
            sr => \N__10137\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10612\,
            in1 => \N__10681\,
            in2 => \_gnd_net_\,
            in3 => \N__10466\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10237\,
            ce => \N__10213\,
            sr => \N__10129\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10301\,
            in1 => \N__10467\,
            in2 => \_gnd_net_\,
            in3 => \N__10515\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10237\,
            ce => \N__10213\,
            sr => \N__10129\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10677\,
            in1 => \N__10465\,
            in2 => \_gnd_net_\,
            in3 => \N__10733\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10211\,
            sr => \N__10124\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10675\,
            in1 => \N__10417\,
            in2 => \_gnd_net_\,
            in3 => \N__10625\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10218\,
            sr => \N__10143\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10553\,
            in1 => \N__10474\,
            in2 => \_gnd_net_\,
            in3 => \N__10514\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__10216\,
            sr => \N__10138\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10458\,
            in1 => \N__10318\,
            in2 => \_gnd_net_\,
            in3 => \N__10283\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10236\,
            ce => \N__10219\,
            sr => \N__10151\
        );

    \U712_BUFFERS.un1_DRDENn_0_a3_LC_24_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__11049\,
            in1 => \_gnd_net_\,
            in2 => \N__10879\,
            in3 => \N__10008\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_0_m2_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100001111"
        )
    port map (
            in0 => \N__11121\,
            in1 => \N__11048\,
            in2 => \N__11005\,
            in3 => \N__10867\,
            lcout => \N_268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

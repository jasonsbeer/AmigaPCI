// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Feb 9 2025 17:04:52

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    TT,
    A,
    CIACS1n,
    TICK50,
    RAMSPACEn,
    TICK60,
    CLKCIA,
    CIACS0n,
    CLK6,
    CLK40_IN,
    CLK28_IN,
    REGSPACEn,
    BUFENn,
    TSn,
    RESETn,
    OVL,
    TACKn,
    ROMENn,
    PORTSIZE);

    input [1:0] TT;
    input [31:1] A;
    output CIACS1n;
    output TICK50;
    output RAMSPACEn;
    output TICK60;
    output CLKCIA;
    output CIACS0n;
    input CLK6;
    input CLK40_IN;
    input CLK28_IN;
    output REGSPACEn;
    output BUFENn;
    input TSn;
    input RESETn;
    input OVL;
    inout TACKn;
    output ROMENn;
    output PORTSIZE;

    wire N__6394;
    wire N__6393;
    wire N__6392;
    wire N__6384;
    wire N__6383;
    wire N__6382;
    wire N__6373;
    wire N__6372;
    wire N__6371;
    wire N__6364;
    wire N__6363;
    wire N__6362;
    wire N__6355;
    wire N__6354;
    wire N__6353;
    wire N__6346;
    wire N__6345;
    wire N__6344;
    wire N__6337;
    wire N__6336;
    wire N__6335;
    wire N__6328;
    wire N__6327;
    wire N__6326;
    wire N__6319;
    wire N__6318;
    wire N__6317;
    wire N__6310;
    wire N__6309;
    wire N__6308;
    wire N__6301;
    wire N__6300;
    wire N__6299;
    wire N__6292;
    wire N__6291;
    wire N__6290;
    wire N__6283;
    wire N__6282;
    wire N__6281;
    wire N__6274;
    wire N__6273;
    wire N__6272;
    wire N__6265;
    wire N__6264;
    wire N__6263;
    wire N__6256;
    wire N__6255;
    wire N__6254;
    wire N__6247;
    wire N__6246;
    wire N__6245;
    wire N__6238;
    wire N__6237;
    wire N__6236;
    wire N__6229;
    wire N__6228;
    wire N__6227;
    wire N__6220;
    wire N__6219;
    wire N__6218;
    wire N__6211;
    wire N__6210;
    wire N__6209;
    wire N__6202;
    wire N__6201;
    wire N__6200;
    wire N__6193;
    wire N__6192;
    wire N__6191;
    wire N__6184;
    wire N__6183;
    wire N__6182;
    wire N__6175;
    wire N__6174;
    wire N__6173;
    wire N__6166;
    wire N__6165;
    wire N__6164;
    wire N__6157;
    wire N__6156;
    wire N__6155;
    wire N__6148;
    wire N__6147;
    wire N__6146;
    wire N__6139;
    wire N__6138;
    wire N__6137;
    wire N__6130;
    wire N__6129;
    wire N__6128;
    wire N__6121;
    wire N__6120;
    wire N__6119;
    wire N__6112;
    wire N__6111;
    wire N__6110;
    wire N__6103;
    wire N__6102;
    wire N__6101;
    wire N__6094;
    wire N__6093;
    wire N__6092;
    wire N__6085;
    wire N__6084;
    wire N__6083;
    wire N__6076;
    wire N__6075;
    wire N__6074;
    wire N__6067;
    wire N__6066;
    wire N__6065;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6036;
    wire N__6035;
    wire N__6032;
    wire N__6029;
    wire N__6024;
    wire N__6023;
    wire N__6022;
    wire N__6021;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6006;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5990;
    wire N__5987;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5977;
    wire N__5976;
    wire N__5975;
    wire N__5974;
    wire N__5973;
    wire N__5972;
    wire N__5971;
    wire N__5970;
    wire N__5969;
    wire N__5968;
    wire N__5967;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5949;
    wire N__5946;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5925;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5881;
    wire N__5878;
    wire N__5873;
    wire N__5868;
    wire N__5865;
    wire N__5864;
    wire N__5863;
    wire N__5862;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5848;
    wire N__5841;
    wire N__5840;
    wire N__5837;
    wire N__5834;
    wire N__5829;
    wire N__5826;
    wire N__5823;
    wire N__5820;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5802;
    wire N__5799;
    wire N__5796;
    wire N__5793;
    wire N__5790;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5772;
    wire N__5771;
    wire N__5770;
    wire N__5769;
    wire N__5766;
    wire N__5763;
    wire N__5758;
    wire N__5751;
    wire N__5748;
    wire N__5745;
    wire N__5742;
    wire N__5741;
    wire N__5740;
    wire N__5739;
    wire N__5738;
    wire N__5735;
    wire N__5726;
    wire N__5721;
    wire N__5720;
    wire N__5719;
    wire N__5718;
    wire N__5717;
    wire N__5716;
    wire N__5707;
    wire N__5702;
    wire N__5697;
    wire N__5696;
    wire N__5695;
    wire N__5694;
    wire N__5693;
    wire N__5690;
    wire N__5689;
    wire N__5680;
    wire N__5675;
    wire N__5670;
    wire N__5667;
    wire N__5666;
    wire N__5665;
    wire N__5664;
    wire N__5663;
    wire N__5656;
    wire N__5651;
    wire N__5646;
    wire N__5643;
    wire N__5642;
    wire N__5641;
    wire N__5640;
    wire N__5639;
    wire N__5636;
    wire N__5633;
    wire N__5630;
    wire N__5627;
    wire N__5624;
    wire N__5619;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5598;
    wire N__5593;
    wire N__5586;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5574;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5559;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5544;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5532;
    wire N__5529;
    wire N__5528;
    wire N__5527;
    wire N__5526;
    wire N__5523;
    wire N__5516;
    wire N__5511;
    wire N__5508;
    wire N__5507;
    wire N__5504;
    wire N__5503;
    wire N__5500;
    wire N__5495;
    wire N__5490;
    wire N__5487;
    wire N__5484;
    wire N__5481;
    wire N__5478;
    wire N__5475;
    wire N__5472;
    wire N__5469;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5459;
    wire N__5456;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5438;
    wire N__5433;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5409;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5397;
    wire N__5394;
    wire N__5391;
    wire N__5388;
    wire N__5387;
    wire N__5384;
    wire N__5381;
    wire N__5376;
    wire N__5373;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5355;
    wire N__5354;
    wire N__5351;
    wire N__5346;
    wire N__5343;
    wire N__5342;
    wire N__5339;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5310;
    wire N__5307;
    wire N__5304;
    wire N__5303;
    wire N__5302;
    wire N__5301;
    wire N__5300;
    wire N__5299;
    wire N__5298;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5282;
    wire N__5275;
    wire N__5268;
    wire N__5267;
    wire N__5266;
    wire N__5265;
    wire N__5264;
    wire N__5263;
    wire N__5254;
    wire N__5249;
    wire N__5244;
    wire N__5243;
    wire N__5242;
    wire N__5241;
    wire N__5240;
    wire N__5239;
    wire N__5238;
    wire N__5229;
    wire N__5222;
    wire N__5217;
    wire N__5214;
    wire N__5213;
    wire N__5208;
    wire N__5205;
    wire N__5204;
    wire N__5203;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5191;
    wire N__5184;
    wire N__5183;
    wire N__5182;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5166;
    wire N__5163;
    wire N__5160;
    wire N__5159;
    wire N__5158;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5142;
    wire N__5139;
    wire N__5136;
    wire N__5135;
    wire N__5134;
    wire N__5131;
    wire N__5126;
    wire N__5121;
    wire N__5118;
    wire N__5117;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5091;
    wire N__5090;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5075;
    wire N__5074;
    wire N__5073;
    wire N__5070;
    wire N__5065;
    wire N__5062;
    wire N__5055;
    wire N__5054;
    wire N__5051;
    wire N__5050;
    wire N__5047;
    wire N__5046;
    wire N__5041;
    wire N__5036;
    wire N__5031;
    wire N__5030;
    wire N__5029;
    wire N__5028;
    wire N__5023;
    wire N__5018;
    wire N__5013;
    wire N__5010;
    wire N__5007;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4986;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4956;
    wire N__4955;
    wire N__4954;
    wire N__4953;
    wire N__4952;
    wire N__4951;
    wire N__4950;
    wire N__4949;
    wire N__4944;
    wire N__4939;
    wire N__4930;
    wire N__4923;
    wire N__4922;
    wire N__4921;
    wire N__4920;
    wire N__4919;
    wire N__4918;
    wire N__4915;
    wire N__4914;
    wire N__4913;
    wire N__4902;
    wire N__4895;
    wire N__4890;
    wire N__4889;
    wire N__4888;
    wire N__4885;
    wire N__4884;
    wire N__4883;
    wire N__4882;
    wire N__4881;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4862;
    wire N__4855;
    wire N__4848;
    wire N__4845;
    wire N__4842;
    wire N__4839;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4827;
    wire N__4826;
    wire N__4825;
    wire N__4824;
    wire N__4823;
    wire N__4822;
    wire N__4821;
    wire N__4820;
    wire N__4819;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4761;
    wire N__4760;
    wire N__4759;
    wire N__4756;
    wire N__4753;
    wire N__4748;
    wire N__4747;
    wire N__4746;
    wire N__4741;
    wire N__4736;
    wire N__4731;
    wire N__4730;
    wire N__4729;
    wire N__4724;
    wire N__4721;
    wire N__4716;
    wire N__4715;
    wire N__4714;
    wire N__4713;
    wire N__4710;
    wire N__4709;
    wire N__4704;
    wire N__4701;
    wire N__4696;
    wire N__4689;
    wire N__4688;
    wire N__4687;
    wire N__4686;
    wire N__4685;
    wire N__4682;
    wire N__4681;
    wire N__4676;
    wire N__4667;
    wire N__4662;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4650;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4638;
    wire N__4635;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4627;
    wire N__4626;
    wire N__4621;
    wire N__4618;
    wire N__4615;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4596;
    wire N__4593;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4575;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4542;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4530;
    wire N__4527;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4485;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4473;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4461;
    wire N__4458;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4446;
    wire N__4445;
    wire N__4442;
    wire N__4439;
    wire N__4434;
    wire N__4433;
    wire N__4430;
    wire N__4429;
    wire N__4428;
    wire N__4427;
    wire N__4426;
    wire N__4425;
    wire N__4424;
    wire N__4417;
    wire N__4408;
    wire N__4405;
    wire N__4398;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4386;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4374;
    wire N__4371;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4359;
    wire N__4356;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4344;
    wire N__4343;
    wire N__4342;
    wire N__4341;
    wire N__4340;
    wire N__4337;
    wire N__4336;
    wire N__4333;
    wire N__4332;
    wire N__4331;
    wire N__4324;
    wire N__4315;
    wire N__4312;
    wire N__4305;
    wire N__4304;
    wire N__4299;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4289;
    wire N__4288;
    wire N__4285;
    wire N__4280;
    wire N__4275;
    wire N__4274;
    wire N__4269;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4251;
    wire N__4248;
    wire N__4247;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4232;
    wire N__4229;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4212;
    wire N__4209;
    wire N__4206;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4191;
    wire N__4188;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4170;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4158;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4146;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4138;
    wire N__4133;
    wire N__4130;
    wire N__4125;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4113;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4101;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4086;
    wire N__4085;
    wire N__4082;
    wire N__4081;
    wire N__4080;
    wire N__4077;
    wire N__4072;
    wire N__4069;
    wire N__4066;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4041;
    wire N__4038;
    wire N__4037;
    wire N__4034;
    wire N__4031;
    wire N__4026;
    wire N__4025;
    wire N__4024;
    wire N__4023;
    wire N__4022;
    wire N__4021;
    wire N__4020;
    wire N__4013;
    wire N__4004;
    wire N__3999;
    wire N__3996;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3984;
    wire N__3981;
    wire N__3978;
    wire N__3975;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3963;
    wire N__3960;
    wire N__3957;
    wire N__3954;
    wire N__3953;
    wire N__3950;
    wire N__3947;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3912;
    wire N__3911;
    wire N__3908;
    wire N__3905;
    wire N__3900;
    wire N__3897;
    wire N__3896;
    wire N__3895;
    wire N__3890;
    wire N__3887;
    wire N__3882;
    wire N__3881;
    wire N__3878;
    wire N__3877;
    wire N__3876;
    wire N__3873;
    wire N__3870;
    wire N__3865;
    wire N__3862;
    wire N__3855;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3843;
    wire N__3840;
    wire N__3839;
    wire N__3836;
    wire N__3833;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3821;
    wire N__3818;
    wire N__3815;
    wire N__3810;
    wire N__3807;
    wire N__3804;
    wire N__3801;
    wire N__3798;
    wire N__3795;
    wire N__3792;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3761;
    wire N__3758;
    wire N__3755;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3743;
    wire N__3738;
    wire N__3735;
    wire N__3732;
    wire N__3729;
    wire N__3726;
    wire N__3723;
    wire N__3720;
    wire N__3717;
    wire N__3714;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3696;
    wire N__3693;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3681;
    wire N__3678;
    wire N__3675;
    wire N__3672;
    wire N__3669;
    wire N__3666;
    wire N__3663;
    wire N__3660;
    wire N__3657;
    wire N__3654;
    wire N__3651;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3639;
    wire N__3638;
    wire N__3637;
    wire N__3634;
    wire N__3631;
    wire N__3628;
    wire N__3621;
    wire N__3618;
    wire N__3615;
    wire N__3612;
    wire N__3611;
    wire N__3610;
    wire N__3605;
    wire N__3602;
    wire N__3597;
    wire N__3596;
    wire N__3595;
    wire N__3592;
    wire N__3591;
    wire N__3586;
    wire N__3581;
    wire N__3576;
    wire N__3575;
    wire N__3574;
    wire N__3573;
    wire N__3572;
    wire N__3567;
    wire N__3564;
    wire N__3559;
    wire N__3552;
    wire N__3549;
    wire N__3546;
    wire N__3543;
    wire N__3542;
    wire N__3541;
    wire N__3540;
    wire N__3539;
    wire N__3538;
    wire N__3535;
    wire N__3530;
    wire N__3527;
    wire N__3522;
    wire N__3513;
    wire N__3512;
    wire N__3511;
    wire N__3510;
    wire N__3507;
    wire N__3504;
    wire N__3499;
    wire N__3492;
    wire N__3489;
    wire N__3486;
    wire N__3483;
    wire N__3480;
    wire N__3477;
    wire N__3474;
    wire N__3471;
    wire N__3468;
    wire N__3465;
    wire N__3462;
    wire N__3459;
    wire N__3456;
    wire N__3453;
    wire N__3450;
    wire N__3447;
    wire N__3444;
    wire N__3441;
    wire N__3438;
    wire N__3435;
    wire N__3432;
    wire N__3429;
    wire N__3426;
    wire N__3423;
    wire N__3422;
    wire N__3421;
    wire N__3414;
    wire N__3411;
    wire N__3408;
    wire N__3407;
    wire N__3406;
    wire N__3405;
    wire N__3398;
    wire N__3395;
    wire N__3392;
    wire N__3389;
    wire N__3388;
    wire N__3385;
    wire N__3382;
    wire N__3379;
    wire N__3378;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3362;
    wire N__3357;
    wire N__3354;
    wire N__3351;
    wire N__3348;
    wire N__3345;
    wire N__3342;
    wire N__3341;
    wire N__3338;
    wire N__3337;
    wire N__3330;
    wire N__3327;
    wire N__3324;
    wire N__3321;
    wire N__3318;
    wire N__3315;
    wire N__3312;
    wire N__3309;
    wire N__3306;
    wire N__3303;
    wire N__3300;
    wire N__3299;
    wire N__3296;
    wire N__3293;
    wire N__3290;
    wire N__3289;
    wire N__3286;
    wire N__3283;
    wire N__3280;
    wire N__3273;
    wire N__3272;
    wire N__3271;
    wire N__3270;
    wire N__3269;
    wire N__3266;
    wire N__3263;
    wire N__3262;
    wire N__3259;
    wire N__3256;
    wire N__3249;
    wire N__3246;
    wire N__3243;
    wire N__3240;
    wire N__3231;
    wire N__3228;
    wire N__3225;
    wire N__3224;
    wire N__3221;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3211;
    wire N__3208;
    wire N__3203;
    wire N__3198;
    wire N__3195;
    wire N__3192;
    wire N__3189;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3171;
    wire N__3168;
    wire N__3165;
    wire N__3164;
    wire N__3163;
    wire N__3160;
    wire N__3157;
    wire N__3154;
    wire N__3151;
    wire N__3146;
    wire N__3143;
    wire N__3140;
    wire N__3137;
    wire N__3134;
    wire N__3129;
    wire N__3126;
    wire N__3123;
    wire N__3120;
    wire N__3117;
    wire N__3114;
    wire N__3111;
    wire N__3108;
    wire N__3107;
    wire N__3104;
    wire N__3101;
    wire N__3098;
    wire N__3095;
    wire N__3090;
    wire N__3087;
    wire N__3084;
    wire N__3081;
    wire N__3078;
    wire N__3075;
    wire N__3072;
    wire N__3069;
    wire N__3066;
    wire N__3063;
    wire N__3060;
    wire N__3059;
    wire N__3058;
    wire N__3055;
    wire N__3054;
    wire N__3053;
    wire N__3052;
    wire N__3049;
    wire N__3046;
    wire N__3043;
    wire N__3040;
    wire N__3035;
    wire N__3032;
    wire N__3029;
    wire N__3028;
    wire N__3023;
    wire N__3020;
    wire N__3015;
    wire N__3012;
    wire N__3007;
    wire N__3000;
    wire N__2997;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2984;
    wire N__2981;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2966;
    wire N__2961;
    wire N__2958;
    wire N__2955;
    wire N__2952;
    wire N__2949;
    wire N__2946;
    wire N__2943;
    wire N__2942;
    wire N__2937;
    wire N__2936;
    wire N__2933;
    wire N__2930;
    wire N__2925;
    wire N__2922;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2909;
    wire N__2906;
    wire N__2905;
    wire N__2900;
    wire N__2897;
    wire N__2892;
    wire N__2889;
    wire N__2886;
    wire N__2883;
    wire N__2880;
    wire N__2877;
    wire N__2876;
    wire N__2873;
    wire N__2870;
    wire N__2869;
    wire N__2866;
    wire N__2861;
    wire N__2856;
    wire N__2853;
    wire N__2852;
    wire N__2851;
    wire N__2846;
    wire N__2843;
    wire N__2840;
    wire N__2837;
    wire N__2832;
    wire N__2829;
    wire N__2826;
    wire N__2823;
    wire N__2820;
    wire N__2817;
    wire N__2814;
    wire N__2813;
    wire N__2810;
    wire N__2805;
    wire N__2802;
    wire N__2799;
    wire N__2796;
    wire N__2793;
    wire N__2792;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2778;
    wire N__2775;
    wire N__2772;
    wire N__2769;
    wire N__2766;
    wire N__2765;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2755;
    wire N__2752;
    wire N__2747;
    wire N__2742;
    wire N__2739;
    wire N__2738;
    wire N__2735;
    wire N__2732;
    wire N__2727;
    wire N__2724;
    wire N__2721;
    wire N__2718;
    wire N__2715;
    wire N__2712;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2702;
    wire N__2701;
    wire N__2698;
    wire N__2693;
    wire N__2690;
    wire N__2687;
    wire N__2684;
    wire N__2681;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2669;
    wire N__2666;
    wire N__2663;
    wire N__2660;
    wire N__2659;
    wire N__2656;
    wire N__2653;
    wire N__2650;
    wire N__2647;
    wire N__2642;
    wire N__2637;
    wire N__2636;
    wire N__2635;
    wire N__2634;
    wire N__2631;
    wire N__2626;
    wire N__2623;
    wire N__2616;
    wire N__2613;
    wire N__2610;
    wire N__2607;
    wire N__2604;
    wire N__2601;
    wire N__2598;
    wire N__2597;
    wire N__2596;
    wire N__2591;
    wire N__2588;
    wire N__2585;
    wire N__2582;
    wire N__2577;
    wire N__2574;
    wire N__2571;
    wire N__2570;
    wire N__2565;
    wire N__2564;
    wire N__2561;
    wire N__2558;
    wire N__2553;
    wire N__2550;
    wire N__2547;
    wire N__2544;
    wire N__2543;
    wire N__2542;
    wire N__2541;
    wire N__2540;
    wire N__2539;
    wire N__2538;
    wire N__2537;
    wire N__2536;
    wire N__2535;
    wire N__2534;
    wire N__2533;
    wire N__2532;
    wire N__2531;
    wire N__2530;
    wire N__2499;
    wire CLK80_OUT;
    wire GNDG0;
    wire VCCG0;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_ ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3 ;
    wire A_c_30;
    wire A_c_29;
    wire A_c_28;
    wire \U409_CIA.g0Z0Z_2_cascade_ ;
    wire A_c_26;
    wire A_c_27;
    wire A_c_24;
    wire \U409_CIA.g0Z0Z_10 ;
    wire \U409_CIA.g0Z0Z_8_cascade_ ;
    wire A_c_16;
    wire A_c_17;
    wire A_c_25;
    wire A_c_18;
    wire \U409_CIA.g0Z0Z_11 ;
    wire A_c_19;
    wire A_c_20;
    wire A_c_21;
    wire CIA_SPACEm_3;
    wire A_c_22;
    wire CIA_SPACEm_6;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_8 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_9 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_10_cascade_ ;
    wire TT_c_1;
    wire A_c_31;
    wire TT_c_0;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_11 ;
    wire \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3 ;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn_i;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ;
    wire A_c_23;
    wire PORTSIZE_0_i;
    wire \U409_ADDRESS_DECODE.un1_REGSPACEnZ0 ;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn_i;
    wire U409_ADDRESS_DECODE_un5_RAMSPACEn;
    wire U409_ADDRESS_DECODE_Z2_SPACE;
    wire U409_ADDRESS_DECODE_HIROM;
    wire OVL_c;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ;
    wire bfn_10_8_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire bfn_10_9_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_11 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_2_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_5 ;
    wire TACKn_in;
    wire BUFENn_c;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_CIACS1n_i;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_CIACS0n_i;
    wire \U409_TICK.TICK503_8 ;
    wire \U409_TICK.TICK503_11_cascade_ ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire TICK50_c;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire bfn_11_6_0_;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire bfn_11_7_0_;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire \U409_TICK.TICK603_11 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.TICK603_8_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire TICK60_c;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.TICK603_9 ;
    wire CIA_ENABLEm;
    wire \U409_CIA.CIA_HOLDZ0 ;
    wire \U409_CIA.g0Z0Z_14 ;
    wire \U409_CIA.g0Z0Z_13 ;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ;
    wire ROMENn_c;
    wire \INVU409_TRANSFER_ACK.ROMENnC_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire CONSTANT_ONE_NET;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire CLK6_c_g;
    wire bfn_12_9_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a2_2 ;
    wire \U409_CIA.N_20_cascade_ ;
    wire \U409_CIA.CLKCIAZ0_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CLKCIA6_0_a2_1 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.N_9_cascade_ ;
    wire \U409_CIA.CLKCIA8_0_a2_0 ;
    wire \U409_CIA.VMAZ0 ;
    wire CLK28_IN_c_g;
    wire CLKCIA_c;
    wire \INVU409_TRANSFER_ACK.LASTCLK_0C_net ;
    wire \U409_TRANSFER_ACK.i6_mux_0_cascade_ ;
    wire \U409_TRANSFER_ACK.N_132_cascade_ ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_4 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_4_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \U409_TRANSFER_ACK.m9_am_cascade_ ;
    wire \U409_TRANSFER_ACK.m9_bm ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_1C_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER15Z0Z_1 ;
    wire TSn_c;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_14 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ;
    wire CLK40_IN_c;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_132 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ;
    wire RESETn_c_i;
    wire \U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ;
    wire \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ;
    wire TACK_OUTn;
    wire \INVU409_TRANSFER_ACK.TACK_OUTnC_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire RESETn_c;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6 ;
    wire \INVU409_TRANSFER_ACK.TACK_EN_iC_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ;
    wire TACK_EN_i;
    wire N_359_i;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__5376),
            .RESETB(N__4596),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6392),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__6394),
            .DIN(N__6393),
            .DOUT(N__6392),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__6394),
            .PADOUT(N__6393),
            .PADIN(N__6392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6382),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__6384),
            .DIN(N__6383),
            .DOUT(N__6382),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__6384),
            .PADOUT(N__6383),
            .PADIN(N__6382),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__6373),
            .DIN(N__6372),
            .DOUT(N__6371),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__6373),
            .PADOUT(N__6372),
            .PADIN(N__6371),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKCIA_obuf_iopad (
            .OE(N__6364),
            .DIN(N__6363),
            .DOUT(N__6362),
            .PACKAGEPIN(CLKCIA));
    defparam CLKCIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKCIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKCIA_obuf_preio (
            .PADOEN(N__6364),
            .PADOUT(N__6363),
            .PADIN(N__6362),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5169),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__6355),
            .DIN(N__6354),
            .DOUT(N__6353),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__6355),
            .PADOUT(N__6354),
            .PADIN(N__6353),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__6346),
            .DIN(N__6345),
            .DOUT(N__6344),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__6346),
            .PADOUT(N__6345),
            .PADIN(N__6344),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS1n_obuf_iopad (
            .OE(N__6337),
            .DIN(N__6336),
            .DOUT(N__6335),
            .PACKAGEPIN(CIACS1n));
    defparam CIACS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS1n_obuf_preio (
            .PADOEN(N__6337),
            .PADOUT(N__6336),
            .PADIN(N__6335),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3720),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_obuf_iopad (
            .OE(N__6328),
            .DIN(N__6327),
            .DOUT(N__6326),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGSPACEn_obuf_preio (
            .PADOEN(N__6328),
            .PADOUT(N__6327),
            .PADIN(N__6326),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3090),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__6319),
            .DIN(N__6318),
            .DOUT(N__6317),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__6319),
            .PADOUT(N__6318),
            .PADIN(N__6317),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__6310),
            .DIN(N__6309),
            .DOUT(N__6308),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__6310),
            .PADOUT(N__6309),
            .PADIN(N__6308),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_obuf_iopad (
            .OE(N__6301),
            .DIN(N__6300),
            .DOUT(N__6299),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMSPACEn_obuf_preio (
            .PADOEN(N__6301),
            .PADOUT(N__6300),
            .PADIN(N__6299),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2961),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_iobuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__6292),
            .DIN(N__6291),
            .DOUT(N__6290),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__6292),
            .PADOUT(N__6291),
            .PADIN(N__6290),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5811),
            .DIN0(TACKn_in),
            .DOUT0(N__6045),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__6283),
            .DIN(N__6282),
            .DOUT(N__6281),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__6283),
            .PADOUT(N__6282),
            .PADIN(N__6281),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ROMENn_obuf_iopad (
            .OE(N__6274),
            .DIN(N__6273),
            .DOUT(N__6272),
            .PACKAGEPIN(ROMENn));
    defparam ROMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ROMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ROMENn_obuf_preio (
            .PADOEN(N__6274),
            .PADOUT(N__6273),
            .PADIN(N__6272),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4782),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__6265),
            .DIN(N__6264),
            .DOUT(N__6263),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__6265),
            .PADOUT(N__6264),
            .PADIN(N__6263),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__6256),
            .DIN(N__6255),
            .DOUT(N__6254),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__6256),
            .PADOUT(N__6255),
            .PADIN(N__6254),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__6247),
            .DIN(N__6246),
            .DOUT(N__6245),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__6247),
            .PADOUT(N__6246),
            .PADIN(N__6245),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3771),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__6238),
            .DIN(N__6237),
            .DOUT(N__6236),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__6238),
            .PADOUT(N__6237),
            .PADIN(N__6236),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2997),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__6229),
            .DIN(N__6228),
            .DOUT(N__6227),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__6229),
            .PADOUT(N__6228),
            .PADIN(N__6227),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__6220),
            .DIN(N__6219),
            .DOUT(N__6218),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__6220),
            .PADOUT(N__6219),
            .PADIN(N__6218),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__6211),
            .DIN(N__6210),
            .DOUT(N__6209),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__6211),
            .PADOUT(N__6210),
            .PADIN(N__6209),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__6202),
            .DIN(N__6201),
            .DOUT(N__6200),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__6202),
            .PADOUT(N__6201),
            .PADIN(N__6200),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__6193),
            .DIN(N__6192),
            .DOUT(N__6191),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__6193),
            .PADOUT(N__6192),
            .PADIN(N__6191),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__6184),
            .DIN(N__6183),
            .DOUT(N__6182),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__6184),
            .PADOUT(N__6183),
            .PADIN(N__6182),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__6175),
            .DIN(N__6174),
            .DOUT(N__6173),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__6175),
            .PADOUT(N__6174),
            .PADIN(N__6173),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__6166),
            .DIN(N__6165),
            .DOUT(N__6164),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__6166),
            .PADOUT(N__6165),
            .PADIN(N__6164),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__6157),
            .DIN(N__6156),
            .DOUT(N__6155),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__6157),
            .PADOUT(N__6156),
            .PADIN(N__6155),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS0n_obuf_iopad (
            .OE(N__6148),
            .DIN(N__6147),
            .DOUT(N__6146),
            .PACKAGEPIN(CIACS0n));
    defparam CIACS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS0n_obuf_preio (
            .PADOEN(N__6148),
            .PADOUT(N__6147),
            .PADIN(N__6146),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3681),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__6139),
            .DIN(N__6138),
            .DOUT(N__6137),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__6139),
            .PADOUT(N__6138),
            .PADIN(N__6137),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3918),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__6130),
            .DIN(N__6129),
            .DOUT(N__6128),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__6130),
            .PADOUT(N__6129),
            .PADIN(N__6128),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__6121),
            .DIN(N__6120),
            .DOUT(N__6119),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__6121),
            .PADOUT(N__6120),
            .PADIN(N__6119),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__6112),
            .DIN(N__6111),
            .DOUT(N__6110),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__6112),
            .PADOUT(N__6111),
            .PADIN(N__6110),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__6103),
            .DIN(N__6102),
            .DOUT(N__6101),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__6103),
            .PADOUT(N__6102),
            .PADIN(N__6101),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__6094),
            .DIN(N__6093),
            .DOUT(N__6092),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__6094),
            .PADOUT(N__6093),
            .PADIN(N__6092),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__6085),
            .DIN(N__6084),
            .DOUT(N__6083),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__6085),
            .PADOUT(N__6084),
            .PADIN(N__6083),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4512),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__6076),
            .DIN(N__6075),
            .DOUT(N__6074),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__6076),
            .PADOUT(N__6075),
            .PADIN(N__6074),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__6067),
            .DIN(N__6066),
            .DOUT(N__6065),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__6067),
            .PADOUT(N__6066),
            .PADIN(N__6065),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__1404 (
            .O(N__6048),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ));
    IoInMux I__1403 (
            .O(N__6045),
            .I(N__6042));
    LocalMux I__1402 (
            .O(N__6042),
            .I(N__6039));
    Span12Mux_s1_v I__1401 (
            .O(N__6039),
            .I(N__6036));
    Span12Mux_v I__1400 (
            .O(N__6036),
            .I(N__6032));
    InMux I__1399 (
            .O(N__6035),
            .I(N__6029));
    Odrv12 I__1398 (
            .O(N__6032),
            .I(TACK_OUTn));
    LocalMux I__1397 (
            .O(N__6029),
            .I(TACK_OUTn));
    InMux I__1396 (
            .O(N__6024),
            .I(N__6017));
    InMux I__1395 (
            .O(N__6023),
            .I(N__6014));
    InMux I__1394 (
            .O(N__6022),
            .I(N__6011));
    InMux I__1393 (
            .O(N__6021),
            .I(N__6006));
    InMux I__1392 (
            .O(N__6020),
            .I(N__6006));
    LocalMux I__1391 (
            .O(N__6017),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__1390 (
            .O(N__6014),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__1389 (
            .O(N__6011),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__1388 (
            .O(N__6006),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    InMux I__1387 (
            .O(N__5997),
            .I(N__5994));
    LocalMux I__1386 (
            .O(N__5994),
            .I(N__5991));
    Span4Mux_v I__1385 (
            .O(N__5991),
            .I(N__5987));
    InMux I__1384 (
            .O(N__5990),
            .I(N__5984));
    Span4Mux_h I__1383 (
            .O(N__5987),
            .I(N__5981));
    LocalMux I__1382 (
            .O(N__5984),
            .I(N__5978));
    Span4Mux_h I__1381 (
            .O(N__5981),
            .I(N__5962));
    Span4Mux_v I__1380 (
            .O(N__5978),
            .I(N__5962));
    InMux I__1379 (
            .O(N__5977),
            .I(N__5959));
    InMux I__1378 (
            .O(N__5976),
            .I(N__5956));
    InMux I__1377 (
            .O(N__5975),
            .I(N__5949));
    InMux I__1376 (
            .O(N__5974),
            .I(N__5949));
    InMux I__1375 (
            .O(N__5973),
            .I(N__5949));
    InMux I__1374 (
            .O(N__5972),
            .I(N__5946));
    InMux I__1373 (
            .O(N__5971),
            .I(N__5941));
    InMux I__1372 (
            .O(N__5970),
            .I(N__5941));
    InMux I__1371 (
            .O(N__5969),
            .I(N__5938));
    InMux I__1370 (
            .O(N__5968),
            .I(N__5935));
    InMux I__1369 (
            .O(N__5967),
            .I(N__5932));
    Span4Mux_h I__1368 (
            .O(N__5962),
            .I(N__5925));
    LocalMux I__1367 (
            .O(N__5959),
            .I(N__5925));
    LocalMux I__1366 (
            .O(N__5956),
            .I(N__5925));
    LocalMux I__1365 (
            .O(N__5949),
            .I(N__5918));
    LocalMux I__1364 (
            .O(N__5946),
            .I(N__5918));
    LocalMux I__1363 (
            .O(N__5941),
            .I(N__5918));
    LocalMux I__1362 (
            .O(N__5938),
            .I(N__5915));
    LocalMux I__1361 (
            .O(N__5935),
            .I(N__5912));
    LocalMux I__1360 (
            .O(N__5932),
            .I(N__5909));
    Span4Mux_v I__1359 (
            .O(N__5925),
            .I(N__5906));
    Span4Mux_v I__1358 (
            .O(N__5918),
            .I(N__5901));
    Span4Mux_v I__1357 (
            .O(N__5915),
            .I(N__5901));
    Span12Mux_h I__1356 (
            .O(N__5912),
            .I(N__5898));
    Span12Mux_h I__1355 (
            .O(N__5909),
            .I(N__5895));
    Sp12to4 I__1354 (
            .O(N__5906),
            .I(N__5890));
    Sp12to4 I__1353 (
            .O(N__5901),
            .I(N__5890));
    Span12Mux_v I__1352 (
            .O(N__5898),
            .I(N__5887));
    Span12Mux_v I__1351 (
            .O(N__5895),
            .I(N__5884));
    Span12Mux_h I__1350 (
            .O(N__5890),
            .I(N__5881));
    Span12Mux_h I__1349 (
            .O(N__5887),
            .I(N__5878));
    Span12Mux_h I__1348 (
            .O(N__5884),
            .I(N__5873));
    Span12Mux_v I__1347 (
            .O(N__5881),
            .I(N__5873));
    Odrv12 I__1346 (
            .O(N__5878),
            .I(RESETn_c));
    Odrv12 I__1345 (
            .O(N__5873),
            .I(RESETn_c));
    CascadeMux I__1344 (
            .O(N__5868),
            .I(N__5865));
    InMux I__1343 (
            .O(N__5865),
            .I(N__5858));
    InMux I__1342 (
            .O(N__5864),
            .I(N__5855));
    InMux I__1341 (
            .O(N__5863),
            .I(N__5848));
    InMux I__1340 (
            .O(N__5862),
            .I(N__5848));
    InMux I__1339 (
            .O(N__5861),
            .I(N__5848));
    LocalMux I__1338 (
            .O(N__5858),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__1337 (
            .O(N__5855),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__1336 (
            .O(N__5848),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    InMux I__1335 (
            .O(N__5841),
            .I(N__5837));
    InMux I__1334 (
            .O(N__5840),
            .I(N__5834));
    LocalMux I__1333 (
            .O(N__5837),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    LocalMux I__1332 (
            .O(N__5834),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    CEMux I__1331 (
            .O(N__5829),
            .I(N__5826));
    LocalMux I__1330 (
            .O(N__5826),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ));
    InMux I__1329 (
            .O(N__5823),
            .I(N__5820));
    LocalMux I__1328 (
            .O(N__5820),
            .I(N__5817));
    Span4Mux_v I__1327 (
            .O(N__5817),
            .I(N__5814));
    Odrv4 I__1326 (
            .O(N__5814),
            .I(TACK_EN_i));
    IoInMux I__1325 (
            .O(N__5811),
            .I(N__5808));
    LocalMux I__1324 (
            .O(N__5808),
            .I(N__5805));
    IoSpan4Mux I__1323 (
            .O(N__5805),
            .I(N__5802));
    Span4Mux_s3_v I__1322 (
            .O(N__5802),
            .I(N__5799));
    Span4Mux_v I__1321 (
            .O(N__5799),
            .I(N__5796));
    Span4Mux_v I__1320 (
            .O(N__5796),
            .I(N__5793));
    Odrv4 I__1319 (
            .O(N__5793),
            .I(N_359_i));
    CascadeMux I__1318 (
            .O(N__5790),
            .I(N__5786));
    CascadeMux I__1317 (
            .O(N__5789),
            .I(N__5783));
    InMux I__1316 (
            .O(N__5786),
            .I(N__5780));
    InMux I__1315 (
            .O(N__5783),
            .I(N__5777));
    LocalMux I__1314 (
            .O(N__5780),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ));
    LocalMux I__1313 (
            .O(N__5777),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ));
    InMux I__1312 (
            .O(N__5772),
            .I(N__5766));
    InMux I__1311 (
            .O(N__5771),
            .I(N__5763));
    InMux I__1310 (
            .O(N__5770),
            .I(N__5758));
    InMux I__1309 (
            .O(N__5769),
            .I(N__5758));
    LocalMux I__1308 (
            .O(N__5766),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1307 (
            .O(N__5763),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1306 (
            .O(N__5758),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    CascadeMux I__1305 (
            .O(N__5751),
            .I(N__5748));
    InMux I__1304 (
            .O(N__5748),
            .I(N__5745));
    LocalMux I__1303 (
            .O(N__5745),
            .I(\U409_TRANSFER_ACK.N_132 ));
    InMux I__1302 (
            .O(N__5742),
            .I(N__5735));
    InMux I__1301 (
            .O(N__5741),
            .I(N__5726));
    InMux I__1300 (
            .O(N__5740),
            .I(N__5726));
    InMux I__1299 (
            .O(N__5739),
            .I(N__5726));
    InMux I__1298 (
            .O(N__5738),
            .I(N__5726));
    LocalMux I__1297 (
            .O(N__5735),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__1296 (
            .O(N__5726),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    InMux I__1295 (
            .O(N__5721),
            .I(N__5707));
    InMux I__1294 (
            .O(N__5720),
            .I(N__5707));
    InMux I__1293 (
            .O(N__5719),
            .I(N__5707));
    InMux I__1292 (
            .O(N__5718),
            .I(N__5707));
    InMux I__1291 (
            .O(N__5717),
            .I(N__5702));
    InMux I__1290 (
            .O(N__5716),
            .I(N__5702));
    LocalMux I__1289 (
            .O(N__5707),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1288 (
            .O(N__5702),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    CascadeMux I__1287 (
            .O(N__5697),
            .I(N__5690));
    InMux I__1286 (
            .O(N__5696),
            .I(N__5680));
    InMux I__1285 (
            .O(N__5695),
            .I(N__5680));
    InMux I__1284 (
            .O(N__5694),
            .I(N__5680));
    InMux I__1283 (
            .O(N__5693),
            .I(N__5680));
    InMux I__1282 (
            .O(N__5690),
            .I(N__5675));
    InMux I__1281 (
            .O(N__5689),
            .I(N__5675));
    LocalMux I__1280 (
            .O(N__5680),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1279 (
            .O(N__5675),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    CascadeMux I__1278 (
            .O(N__5670),
            .I(N__5667));
    InMux I__1277 (
            .O(N__5667),
            .I(N__5656));
    InMux I__1276 (
            .O(N__5666),
            .I(N__5656));
    InMux I__1275 (
            .O(N__5665),
            .I(N__5656));
    InMux I__1274 (
            .O(N__5664),
            .I(N__5651));
    InMux I__1273 (
            .O(N__5663),
            .I(N__5651));
    LocalMux I__1272 (
            .O(N__5656),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1271 (
            .O(N__5651),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    SRMux I__1270 (
            .O(N__5646),
            .I(N__5643));
    LocalMux I__1269 (
            .O(N__5643),
            .I(N__5636));
    SRMux I__1268 (
            .O(N__5642),
            .I(N__5633));
    SRMux I__1267 (
            .O(N__5641),
            .I(N__5630));
    SRMux I__1266 (
            .O(N__5640),
            .I(N__5627));
    SRMux I__1265 (
            .O(N__5639),
            .I(N__5624));
    Span4Mux_v I__1264 (
            .O(N__5636),
            .I(N__5619));
    LocalMux I__1263 (
            .O(N__5633),
            .I(N__5619));
    LocalMux I__1262 (
            .O(N__5630),
            .I(N__5615));
    LocalMux I__1261 (
            .O(N__5627),
            .I(N__5612));
    LocalMux I__1260 (
            .O(N__5624),
            .I(N__5607));
    Sp12to4 I__1259 (
            .O(N__5619),
            .I(N__5607));
    SRMux I__1258 (
            .O(N__5618),
            .I(N__5604));
    Span4Mux_h I__1257 (
            .O(N__5615),
            .I(N__5601));
    Span4Mux_h I__1256 (
            .O(N__5612),
            .I(N__5598));
    Span12Mux_h I__1255 (
            .O(N__5607),
            .I(N__5593));
    LocalMux I__1254 (
            .O(N__5604),
            .I(N__5593));
    Odrv4 I__1253 (
            .O(N__5601),
            .I(RESETn_c_i));
    Odrv4 I__1252 (
            .O(N__5598),
            .I(RESETn_c_i));
    Odrv12 I__1251 (
            .O(N__5593),
            .I(RESETn_c_i));
    InMux I__1250 (
            .O(N__5586),
            .I(N__5582));
    InMux I__1249 (
            .O(N__5585),
            .I(N__5579));
    LocalMux I__1248 (
            .O(N__5582),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    LocalMux I__1247 (
            .O(N__5579),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    InMux I__1246 (
            .O(N__5574),
            .I(N__5570));
    InMux I__1245 (
            .O(N__5573),
            .I(N__5567));
    LocalMux I__1244 (
            .O(N__5570),
            .I(N__5564));
    LocalMux I__1243 (
            .O(N__5567),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    Odrv4 I__1242 (
            .O(N__5564),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    CascadeMux I__1241 (
            .O(N__5559),
            .I(N__5555));
    InMux I__1240 (
            .O(N__5558),
            .I(N__5552));
    InMux I__1239 (
            .O(N__5555),
            .I(N__5549));
    LocalMux I__1238 (
            .O(N__5552),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__1237 (
            .O(N__5549),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__1236 (
            .O(N__5544),
            .I(N__5540));
    InMux I__1235 (
            .O(N__5543),
            .I(N__5537));
    LocalMux I__1234 (
            .O(N__5540),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__1233 (
            .O(N__5537),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    CascadeMux I__1232 (
            .O(N__5532),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ));
    InMux I__1231 (
            .O(N__5529),
            .I(N__5523));
    InMux I__1230 (
            .O(N__5528),
            .I(N__5516));
    InMux I__1229 (
            .O(N__5527),
            .I(N__5516));
    InMux I__1228 (
            .O(N__5526),
            .I(N__5516));
    LocalMux I__1227 (
            .O(N__5523),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__1226 (
            .O(N__5516),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    CascadeMux I__1225 (
            .O(N__5511),
            .I(\U409_TRANSFER_ACK.N_4_cascade_ ));
    CascadeMux I__1224 (
            .O(N__5508),
            .I(N__5504));
    InMux I__1223 (
            .O(N__5507),
            .I(N__5500));
    InMux I__1222 (
            .O(N__5504),
            .I(N__5495));
    InMux I__1221 (
            .O(N__5503),
            .I(N__5495));
    LocalMux I__1220 (
            .O(N__5500),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    LocalMux I__1219 (
            .O(N__5495),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    CascadeMux I__1218 (
            .O(N__5490),
            .I(\U409_TRANSFER_ACK.m9_am_cascade_ ));
    InMux I__1217 (
            .O(N__5487),
            .I(N__5484));
    LocalMux I__1216 (
            .O(N__5484),
            .I(\U409_TRANSFER_ACK.m9_bm ));
    InMux I__1215 (
            .O(N__5481),
            .I(N__5478));
    LocalMux I__1214 (
            .O(N__5478),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ));
    InMux I__1213 (
            .O(N__5475),
            .I(N__5472));
    LocalMux I__1212 (
            .O(N__5472),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ));
    InMux I__1211 (
            .O(N__5469),
            .I(N__5466));
    LocalMux I__1210 (
            .O(N__5466),
            .I(N__5463));
    Odrv12 I__1209 (
            .O(N__5463),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER15Z0Z_1 ));
    InMux I__1208 (
            .O(N__5460),
            .I(N__5456));
    InMux I__1207 (
            .O(N__5459),
            .I(N__5452));
    LocalMux I__1206 (
            .O(N__5456),
            .I(N__5449));
    InMux I__1205 (
            .O(N__5455),
            .I(N__5446));
    LocalMux I__1204 (
            .O(N__5452),
            .I(N__5443));
    Span4Mux_h I__1203 (
            .O(N__5449),
            .I(N__5438));
    LocalMux I__1202 (
            .O(N__5446),
            .I(N__5438));
    Span4Mux_h I__1201 (
            .O(N__5443),
            .I(N__5433));
    Span4Mux_h I__1200 (
            .O(N__5438),
            .I(N__5433));
    Span4Mux_h I__1199 (
            .O(N__5433),
            .I(N__5429));
    InMux I__1198 (
            .O(N__5432),
            .I(N__5426));
    Sp12to4 I__1197 (
            .O(N__5429),
            .I(N__5423));
    LocalMux I__1196 (
            .O(N__5426),
            .I(N__5420));
    Span12Mux_v I__1195 (
            .O(N__5423),
            .I(N__5417));
    Sp12to4 I__1194 (
            .O(N__5420),
            .I(N__5414));
    Odrv12 I__1193 (
            .O(N__5417),
            .I(TSn_c));
    Odrv12 I__1192 (
            .O(N__5414),
            .I(TSn_c));
    InMux I__1191 (
            .O(N__5409),
            .I(N__5405));
    InMux I__1190 (
            .O(N__5408),
            .I(N__5402));
    LocalMux I__1189 (
            .O(N__5405),
            .I(N__5397));
    LocalMux I__1188 (
            .O(N__5402),
            .I(N__5397));
    Span4Mux_v I__1187 (
            .O(N__5397),
            .I(N__5394));
    Sp12to4 I__1186 (
            .O(N__5394),
            .I(N__5391));
    Odrv12 I__1185 (
            .O(N__5391),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_14 ));
    InMux I__1184 (
            .O(N__5388),
            .I(N__5384));
    InMux I__1183 (
            .O(N__5387),
            .I(N__5381));
    LocalMux I__1182 (
            .O(N__5384),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    LocalMux I__1181 (
            .O(N__5381),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    IoInMux I__1180 (
            .O(N__5376),
            .I(N__5373));
    LocalMux I__1179 (
            .O(N__5373),
            .I(N__5369));
    CascadeMux I__1178 (
            .O(N__5372),
            .I(N__5366));
    IoSpan4Mux I__1177 (
            .O(N__5369),
            .I(N__5362));
    InMux I__1176 (
            .O(N__5366),
            .I(N__5359));
    InMux I__1175 (
            .O(N__5365),
            .I(N__5356));
    Span4Mux_s0_v I__1174 (
            .O(N__5362),
            .I(N__5351));
    LocalMux I__1173 (
            .O(N__5359),
            .I(N__5346));
    LocalMux I__1172 (
            .O(N__5356),
            .I(N__5346));
    CascadeMux I__1171 (
            .O(N__5355),
            .I(N__5343));
    CascadeMux I__1170 (
            .O(N__5354),
            .I(N__5339));
    Sp12to4 I__1169 (
            .O(N__5351),
            .I(N__5335));
    Span4Mux_h I__1168 (
            .O(N__5346),
            .I(N__5332));
    InMux I__1167 (
            .O(N__5343),
            .I(N__5327));
    InMux I__1166 (
            .O(N__5342),
            .I(N__5327));
    InMux I__1165 (
            .O(N__5339),
            .I(N__5324));
    InMux I__1164 (
            .O(N__5338),
            .I(N__5321));
    Span12Mux_v I__1163 (
            .O(N__5335),
            .I(N__5310));
    Sp12to4 I__1162 (
            .O(N__5332),
            .I(N__5310));
    LocalMux I__1161 (
            .O(N__5327),
            .I(N__5310));
    LocalMux I__1160 (
            .O(N__5324),
            .I(N__5310));
    LocalMux I__1159 (
            .O(N__5321),
            .I(N__5310));
    Span12Mux_v I__1158 (
            .O(N__5310),
            .I(N__5307));
    Odrv12 I__1157 (
            .O(N__5307),
            .I(CLK40_IN_c));
    CascadeMux I__1156 (
            .O(N__5304),
            .I(N__5294));
    InMux I__1155 (
            .O(N__5303),
            .I(N__5291));
    InMux I__1154 (
            .O(N__5302),
            .I(N__5282));
    InMux I__1153 (
            .O(N__5301),
            .I(N__5282));
    InMux I__1152 (
            .O(N__5300),
            .I(N__5282));
    InMux I__1151 (
            .O(N__5299),
            .I(N__5282));
    InMux I__1150 (
            .O(N__5298),
            .I(N__5275));
    InMux I__1149 (
            .O(N__5297),
            .I(N__5275));
    InMux I__1148 (
            .O(N__5294),
            .I(N__5275));
    LocalMux I__1147 (
            .O(N__5291),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1146 (
            .O(N__5282),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1145 (
            .O(N__5275),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    InMux I__1144 (
            .O(N__5268),
            .I(N__5254));
    InMux I__1143 (
            .O(N__5267),
            .I(N__5254));
    InMux I__1142 (
            .O(N__5266),
            .I(N__5254));
    InMux I__1141 (
            .O(N__5265),
            .I(N__5254));
    InMux I__1140 (
            .O(N__5264),
            .I(N__5249));
    InMux I__1139 (
            .O(N__5263),
            .I(N__5249));
    LocalMux I__1138 (
            .O(N__5254),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1137 (
            .O(N__5249),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    InMux I__1136 (
            .O(N__5244),
            .I(N__5229));
    InMux I__1135 (
            .O(N__5243),
            .I(N__5229));
    InMux I__1134 (
            .O(N__5242),
            .I(N__5229));
    InMux I__1133 (
            .O(N__5241),
            .I(N__5229));
    InMux I__1132 (
            .O(N__5240),
            .I(N__5222));
    InMux I__1131 (
            .O(N__5239),
            .I(N__5222));
    InMux I__1130 (
            .O(N__5238),
            .I(N__5222));
    LocalMux I__1129 (
            .O(N__5229),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1128 (
            .O(N__5222),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    CascadeMux I__1127 (
            .O(N__5217),
            .I(\U409_CIA.N_9_cascade_ ));
    InMux I__1126 (
            .O(N__5214),
            .I(N__5208));
    InMux I__1125 (
            .O(N__5213),
            .I(N__5208));
    LocalMux I__1124 (
            .O(N__5208),
            .I(\U409_CIA.CLKCIA8_0_a2_0 ));
    InMux I__1123 (
            .O(N__5205),
            .I(N__5199));
    InMux I__1122 (
            .O(N__5204),
            .I(N__5196));
    InMux I__1121 (
            .O(N__5203),
            .I(N__5191));
    InMux I__1120 (
            .O(N__5202),
            .I(N__5191));
    LocalMux I__1119 (
            .O(N__5199),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__1118 (
            .O(N__5196),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__1117 (
            .O(N__5191),
            .I(\U409_CIA.VMAZ0 ));
    ClkMux I__1116 (
            .O(N__5184),
            .I(N__5175));
    ClkMux I__1115 (
            .O(N__5183),
            .I(N__5175));
    ClkMux I__1114 (
            .O(N__5182),
            .I(N__5175));
    GlobalMux I__1113 (
            .O(N__5175),
            .I(N__5172));
    gio2CtrlBuf I__1112 (
            .O(N__5172),
            .I(CLK28_IN_c_g));
    IoInMux I__1111 (
            .O(N__5169),
            .I(N__5166));
    LocalMux I__1110 (
            .O(N__5166),
            .I(N__5163));
    Span12Mux_s4_v I__1109 (
            .O(N__5163),
            .I(N__5160));
    Span12Mux_v I__1108 (
            .O(N__5160),
            .I(N__5155));
    InMux I__1107 (
            .O(N__5159),
            .I(N__5152));
    InMux I__1106 (
            .O(N__5158),
            .I(N__5149));
    Odrv12 I__1105 (
            .O(N__5155),
            .I(CLKCIA_c));
    LocalMux I__1104 (
            .O(N__5152),
            .I(CLKCIA_c));
    LocalMux I__1103 (
            .O(N__5149),
            .I(CLKCIA_c));
    CascadeMux I__1102 (
            .O(N__5142),
            .I(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ));
    CascadeMux I__1101 (
            .O(N__5139),
            .I(\U409_TRANSFER_ACK.N_132_cascade_ ));
    InMux I__1100 (
            .O(N__5136),
            .I(N__5131));
    InMux I__1099 (
            .O(N__5135),
            .I(N__5126));
    InMux I__1098 (
            .O(N__5134),
            .I(N__5126));
    LocalMux I__1097 (
            .O(N__5131),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__1096 (
            .O(N__5126),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    CascadeMux I__1095 (
            .O(N__5121),
            .I(N__5118));
    InMux I__1094 (
            .O(N__5118),
            .I(N__5112));
    InMux I__1093 (
            .O(N__5117),
            .I(N__5112));
    LocalMux I__1092 (
            .O(N__5112),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    InMux I__1091 (
            .O(N__5109),
            .I(N__5106));
    LocalMux I__1090 (
            .O(N__5106),
            .I(\U409_TRANSFER_ACK.N_4 ));
    CascadeMux I__1089 (
            .O(N__5103),
            .I(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ));
    InMux I__1088 (
            .O(N__5100),
            .I(N__5097));
    LocalMux I__1087 (
            .O(N__5097),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ));
    CascadeMux I__1086 (
            .O(N__5094),
            .I(N__5091));
    InMux I__1085 (
            .O(N__5091),
            .I(N__5085));
    InMux I__1084 (
            .O(N__5090),
            .I(N__5085));
    LocalMux I__1083 (
            .O(N__5085),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ));
    CascadeMux I__1082 (
            .O(N__5082),
            .I(\U409_CIA.N_20_cascade_ ));
    CascadeMux I__1081 (
            .O(N__5079),
            .I(\U409_CIA.CLKCIAZ0_cascade_ ));
    InMux I__1080 (
            .O(N__5076),
            .I(N__5070));
    InMux I__1079 (
            .O(N__5075),
            .I(N__5065));
    InMux I__1078 (
            .O(N__5074),
            .I(N__5065));
    InMux I__1077 (
            .O(N__5073),
            .I(N__5062));
    LocalMux I__1076 (
            .O(N__5070),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1075 (
            .O(N__5065),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1074 (
            .O(N__5062),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    CascadeMux I__1073 (
            .O(N__5055),
            .I(N__5051));
    CascadeMux I__1072 (
            .O(N__5054),
            .I(N__5047));
    InMux I__1071 (
            .O(N__5051),
            .I(N__5041));
    InMux I__1070 (
            .O(N__5050),
            .I(N__5041));
    InMux I__1069 (
            .O(N__5047),
            .I(N__5036));
    InMux I__1068 (
            .O(N__5046),
            .I(N__5036));
    LocalMux I__1067 (
            .O(N__5041),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1066 (
            .O(N__5036),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    InMux I__1065 (
            .O(N__5031),
            .I(N__5023));
    InMux I__1064 (
            .O(N__5030),
            .I(N__5023));
    InMux I__1063 (
            .O(N__5029),
            .I(N__5018));
    InMux I__1062 (
            .O(N__5028),
            .I(N__5018));
    LocalMux I__1061 (
            .O(N__5023),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1060 (
            .O(N__5018),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    InMux I__1059 (
            .O(N__5013),
            .I(N__5010));
    LocalMux I__1058 (
            .O(N__5010),
            .I(\U409_CIA.CLKCIA6_0_a2_1 ));
    InMux I__1057 (
            .O(N__5007),
            .I(N__5003));
    InMux I__1056 (
            .O(N__5006),
            .I(N__5000));
    LocalMux I__1055 (
            .O(N__5003),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__1054 (
            .O(N__5000),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    CascadeMux I__1053 (
            .O(N__4995),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    InMux I__1052 (
            .O(N__4992),
            .I(N__4989));
    LocalMux I__1051 (
            .O(N__4989),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__1050 (
            .O(N__4986),
            .I(N__4982));
    InMux I__1049 (
            .O(N__4985),
            .I(N__4979));
    LocalMux I__1048 (
            .O(N__4982),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__1047 (
            .O(N__4979),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__1046 (
            .O(N__4974),
            .I(N__4971));
    LocalMux I__1045 (
            .O(N__4971),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__1044 (
            .O(N__4968),
            .I(N__4964));
    InMux I__1043 (
            .O(N__4967),
            .I(N__4961));
    LocalMux I__1042 (
            .O(N__4964),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__1041 (
            .O(N__4961),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    InMux I__1040 (
            .O(N__4956),
            .I(N__4944));
    InMux I__1039 (
            .O(N__4955),
            .I(N__4944));
    InMux I__1038 (
            .O(N__4954),
            .I(N__4939));
    InMux I__1037 (
            .O(N__4953),
            .I(N__4939));
    InMux I__1036 (
            .O(N__4952),
            .I(N__4930));
    InMux I__1035 (
            .O(N__4951),
            .I(N__4930));
    InMux I__1034 (
            .O(N__4950),
            .I(N__4930));
    InMux I__1033 (
            .O(N__4949),
            .I(N__4930));
    LocalMux I__1032 (
            .O(N__4944),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__1031 (
            .O(N__4939),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__1030 (
            .O(N__4930),
            .I(\U409_TICK.TICK503_10 ));
    CascadeMux I__1029 (
            .O(N__4923),
            .I(N__4915));
    InMux I__1028 (
            .O(N__4922),
            .I(N__4902));
    InMux I__1027 (
            .O(N__4921),
            .I(N__4902));
    InMux I__1026 (
            .O(N__4920),
            .I(N__4902));
    InMux I__1025 (
            .O(N__4919),
            .I(N__4902));
    InMux I__1024 (
            .O(N__4918),
            .I(N__4902));
    InMux I__1023 (
            .O(N__4915),
            .I(N__4895));
    InMux I__1022 (
            .O(N__4914),
            .I(N__4895));
    InMux I__1021 (
            .O(N__4913),
            .I(N__4895));
    LocalMux I__1020 (
            .O(N__4902),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__1019 (
            .O(N__4895),
            .I(\U409_TICK.TICK503_14 ));
    CascadeMux I__1018 (
            .O(N__4890),
            .I(N__4885));
    CascadeMux I__1017 (
            .O(N__4889),
            .I(N__4877));
    CascadeMux I__1016 (
            .O(N__4888),
            .I(N__4874));
    InMux I__1015 (
            .O(N__4885),
            .I(N__4871));
    InMux I__1014 (
            .O(N__4884),
            .I(N__4862));
    InMux I__1013 (
            .O(N__4883),
            .I(N__4862));
    InMux I__1012 (
            .O(N__4882),
            .I(N__4862));
    InMux I__1011 (
            .O(N__4881),
            .I(N__4862));
    InMux I__1010 (
            .O(N__4880),
            .I(N__4855));
    InMux I__1009 (
            .O(N__4877),
            .I(N__4855));
    InMux I__1008 (
            .O(N__4874),
            .I(N__4855));
    LocalMux I__1007 (
            .O(N__4871),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1006 (
            .O(N__4862),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1005 (
            .O(N__4855),
            .I(\U409_TICK.TICK503_9 ));
    InMux I__1004 (
            .O(N__4848),
            .I(N__4845));
    LocalMux I__1003 (
            .O(N__4845),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    CascadeMux I__1002 (
            .O(N__4842),
            .I(N__4839));
    InMux I__1001 (
            .O(N__4839),
            .I(N__4835));
    InMux I__1000 (
            .O(N__4838),
            .I(N__4832));
    LocalMux I__999 (
            .O(N__4835),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__998 (
            .O(N__4832),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    ClkMux I__997 (
            .O(N__4827),
            .I(N__4800));
    ClkMux I__996 (
            .O(N__4826),
            .I(N__4800));
    ClkMux I__995 (
            .O(N__4825),
            .I(N__4800));
    ClkMux I__994 (
            .O(N__4824),
            .I(N__4800));
    ClkMux I__993 (
            .O(N__4823),
            .I(N__4800));
    ClkMux I__992 (
            .O(N__4822),
            .I(N__4800));
    ClkMux I__991 (
            .O(N__4821),
            .I(N__4800));
    ClkMux I__990 (
            .O(N__4820),
            .I(N__4800));
    ClkMux I__989 (
            .O(N__4819),
            .I(N__4800));
    GlobalMux I__988 (
            .O(N__4800),
            .I(N__4797));
    gio2CtrlBuf I__987 (
            .O(N__4797),
            .I(CLK6_c_g));
    InMux I__986 (
            .O(N__4794),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__985 (
            .O(N__4791),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__984 (
            .O(N__4788),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__983 (
            .O(N__4785),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    IoInMux I__982 (
            .O(N__4782),
            .I(N__4779));
    LocalMux I__981 (
            .O(N__4779),
            .I(N__4776));
    Span12Mux_s1_v I__980 (
            .O(N__4776),
            .I(N__4773));
    Span12Mux_v I__979 (
            .O(N__4773),
            .I(N__4769));
    InMux I__978 (
            .O(N__4772),
            .I(N__4766));
    Odrv12 I__977 (
            .O(N__4769),
            .I(ROMENn_c));
    LocalMux I__976 (
            .O(N__4766),
            .I(ROMENn_c));
    CascadeMux I__975 (
            .O(N__4761),
            .I(N__4756));
    InMux I__974 (
            .O(N__4760),
            .I(N__4753));
    InMux I__973 (
            .O(N__4759),
            .I(N__4748));
    InMux I__972 (
            .O(N__4756),
            .I(N__4748));
    LocalMux I__971 (
            .O(N__4753),
            .I(N__4741));
    LocalMux I__970 (
            .O(N__4748),
            .I(N__4741));
    InMux I__969 (
            .O(N__4747),
            .I(N__4736));
    InMux I__968 (
            .O(N__4746),
            .I(N__4736));
    Odrv4 I__967 (
            .O(N__4741),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__966 (
            .O(N__4736),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    InMux I__965 (
            .O(N__4731),
            .I(N__4724));
    InMux I__964 (
            .O(N__4730),
            .I(N__4724));
    InMux I__963 (
            .O(N__4729),
            .I(N__4721));
    LocalMux I__962 (
            .O(N__4724),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    LocalMux I__961 (
            .O(N__4721),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    CascadeMux I__960 (
            .O(N__4716),
            .I(N__4710));
    InMux I__959 (
            .O(N__4715),
            .I(N__4704));
    InMux I__958 (
            .O(N__4714),
            .I(N__4704));
    InMux I__957 (
            .O(N__4713),
            .I(N__4701));
    InMux I__956 (
            .O(N__4710),
            .I(N__4696));
    InMux I__955 (
            .O(N__4709),
            .I(N__4696));
    LocalMux I__954 (
            .O(N__4704),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__953 (
            .O(N__4701),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__952 (
            .O(N__4696),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    CascadeMux I__951 (
            .O(N__4689),
            .I(N__4682));
    InMux I__950 (
            .O(N__4688),
            .I(N__4676));
    InMux I__949 (
            .O(N__4687),
            .I(N__4676));
    InMux I__948 (
            .O(N__4686),
            .I(N__4667));
    InMux I__947 (
            .O(N__4685),
            .I(N__4667));
    InMux I__946 (
            .O(N__4682),
            .I(N__4667));
    InMux I__945 (
            .O(N__4681),
            .I(N__4667));
    LocalMux I__944 (
            .O(N__4676),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__943 (
            .O(N__4667),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    InMux I__942 (
            .O(N__4662),
            .I(N__4658));
    InMux I__941 (
            .O(N__4661),
            .I(N__4655));
    LocalMux I__940 (
            .O(N__4658),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    LocalMux I__939 (
            .O(N__4655),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    InMux I__938 (
            .O(N__4650),
            .I(N__4646));
    InMux I__937 (
            .O(N__4649),
            .I(N__4643));
    LocalMux I__936 (
            .O(N__4646),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    LocalMux I__935 (
            .O(N__4643),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    SRMux I__934 (
            .O(N__4638),
            .I(N__4635));
    LocalMux I__933 (
            .O(N__4635),
            .I(N__4631));
    SRMux I__932 (
            .O(N__4634),
            .I(N__4628));
    Span4Mux_v I__931 (
            .O(N__4631),
            .I(N__4621));
    LocalMux I__930 (
            .O(N__4628),
            .I(N__4621));
    SRMux I__929 (
            .O(N__4627),
            .I(N__4618));
    SRMux I__928 (
            .O(N__4626),
            .I(N__4615));
    Span4Mux_h I__927 (
            .O(N__4621),
            .I(N__4610));
    LocalMux I__926 (
            .O(N__4618),
            .I(N__4610));
    LocalMux I__925 (
            .O(N__4615),
            .I(N__4607));
    Span4Mux_h I__924 (
            .O(N__4610),
            .I(N__4604));
    Span4Mux_v I__923 (
            .O(N__4607),
            .I(N__4601));
    Odrv4 I__922 (
            .O(N__4604),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv4 I__921 (
            .O(N__4601),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    IoInMux I__920 (
            .O(N__4596),
            .I(N__4593));
    LocalMux I__919 (
            .O(N__4593),
            .I(N__4590));
    Span4Mux_s2_v I__918 (
            .O(N__4590),
            .I(N__4587));
    Span4Mux_v I__917 (
            .O(N__4587),
            .I(N__4584));
    Odrv4 I__916 (
            .O(N__4584),
            .I(CONSTANT_ONE_NET));
    InMux I__915 (
            .O(N__4581),
            .I(N__4578));
    LocalMux I__914 (
            .O(N__4578),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__913 (
            .O(N__4575),
            .I(N__4571));
    InMux I__912 (
            .O(N__4574),
            .I(N__4568));
    LocalMux I__911 (
            .O(N__4571),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__910 (
            .O(N__4568),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    CascadeMux I__909 (
            .O(N__4563),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    InMux I__908 (
            .O(N__4560),
            .I(N__4557));
    LocalMux I__907 (
            .O(N__4557),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__906 (
            .O(N__4554),
            .I(N__4550));
    InMux I__905 (
            .O(N__4553),
            .I(N__4547));
    LocalMux I__904 (
            .O(N__4550),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__903 (
            .O(N__4547),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__902 (
            .O(N__4542),
            .I(N__4538));
    InMux I__901 (
            .O(N__4541),
            .I(N__4535));
    LocalMux I__900 (
            .O(N__4538),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__899 (
            .O(N__4535),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    CascadeMux I__898 (
            .O(N__4530),
            .I(N__4527));
    InMux I__897 (
            .O(N__4527),
            .I(N__4523));
    InMux I__896 (
            .O(N__4526),
            .I(N__4520));
    LocalMux I__895 (
            .O(N__4523),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__894 (
            .O(N__4520),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    CascadeMux I__893 (
            .O(N__4515),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    IoInMux I__892 (
            .O(N__4512),
            .I(N__4509));
    LocalMux I__891 (
            .O(N__4509),
            .I(N__4506));
    Span4Mux_s2_v I__890 (
            .O(N__4506),
            .I(N__4503));
    Sp12to4 I__889 (
            .O(N__4503),
            .I(N__4500));
    Span12Mux_h I__888 (
            .O(N__4500),
            .I(N__4497));
    Span12Mux_v I__887 (
            .O(N__4497),
            .I(N__4493));
    InMux I__886 (
            .O(N__4496),
            .I(N__4490));
    Odrv12 I__885 (
            .O(N__4493),
            .I(TICK60_c));
    LocalMux I__884 (
            .O(N__4490),
            .I(TICK60_c));
    InMux I__883 (
            .O(N__4485),
            .I(N__4481));
    InMux I__882 (
            .O(N__4484),
            .I(N__4478));
    LocalMux I__881 (
            .O(N__4481),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__880 (
            .O(N__4478),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    InMux I__879 (
            .O(N__4473),
            .I(N__4469));
    InMux I__878 (
            .O(N__4472),
            .I(N__4466));
    LocalMux I__877 (
            .O(N__4469),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__876 (
            .O(N__4466),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    CascadeMux I__875 (
            .O(N__4461),
            .I(N__4458));
    InMux I__874 (
            .O(N__4458),
            .I(N__4454));
    InMux I__873 (
            .O(N__4457),
            .I(N__4451));
    LocalMux I__872 (
            .O(N__4454),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__871 (
            .O(N__4451),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__870 (
            .O(N__4446),
            .I(N__4442));
    InMux I__869 (
            .O(N__4445),
            .I(N__4439));
    LocalMux I__868 (
            .O(N__4442),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__867 (
            .O(N__4439),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    CascadeMux I__866 (
            .O(N__4434),
            .I(N__4430));
    InMux I__865 (
            .O(N__4433),
            .I(N__4417));
    InMux I__864 (
            .O(N__4430),
            .I(N__4417));
    InMux I__863 (
            .O(N__4429),
            .I(N__4417));
    InMux I__862 (
            .O(N__4428),
            .I(N__4408));
    InMux I__861 (
            .O(N__4427),
            .I(N__4408));
    InMux I__860 (
            .O(N__4426),
            .I(N__4408));
    InMux I__859 (
            .O(N__4425),
            .I(N__4408));
    InMux I__858 (
            .O(N__4424),
            .I(N__4405));
    LocalMux I__857 (
            .O(N__4417),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__856 (
            .O(N__4408),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__855 (
            .O(N__4405),
            .I(\U409_TICK.TICK603_10 ));
    InMux I__854 (
            .O(N__4398),
            .I(N__4394));
    InMux I__853 (
            .O(N__4397),
            .I(N__4391));
    LocalMux I__852 (
            .O(N__4394),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__851 (
            .O(N__4391),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    InMux I__850 (
            .O(N__4386),
            .I(N__4382));
    InMux I__849 (
            .O(N__4385),
            .I(N__4379));
    LocalMux I__848 (
            .O(N__4382),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__847 (
            .O(N__4379),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    CascadeMux I__846 (
            .O(N__4374),
            .I(N__4371));
    InMux I__845 (
            .O(N__4371),
            .I(N__4367));
    InMux I__844 (
            .O(N__4370),
            .I(N__4364));
    LocalMux I__843 (
            .O(N__4367),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__842 (
            .O(N__4364),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    InMux I__841 (
            .O(N__4359),
            .I(N__4356));
    LocalMux I__840 (
            .O(N__4356),
            .I(N__4352));
    InMux I__839 (
            .O(N__4355),
            .I(N__4349));
    Odrv4 I__838 (
            .O(N__4352),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__837 (
            .O(N__4349),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    CascadeMux I__836 (
            .O(N__4344),
            .I(N__4337));
    CascadeMux I__835 (
            .O(N__4343),
            .I(N__4333));
    InMux I__834 (
            .O(N__4342),
            .I(N__4324));
    InMux I__833 (
            .O(N__4341),
            .I(N__4324));
    InMux I__832 (
            .O(N__4340),
            .I(N__4324));
    InMux I__831 (
            .O(N__4337),
            .I(N__4315));
    InMux I__830 (
            .O(N__4336),
            .I(N__4315));
    InMux I__829 (
            .O(N__4333),
            .I(N__4315));
    InMux I__828 (
            .O(N__4332),
            .I(N__4315));
    InMux I__827 (
            .O(N__4331),
            .I(N__4312));
    LocalMux I__826 (
            .O(N__4324),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__825 (
            .O(N__4315),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__824 (
            .O(N__4312),
            .I(\U409_TICK.TICK603_9 ));
    InMux I__823 (
            .O(N__4305),
            .I(N__4299));
    InMux I__822 (
            .O(N__4304),
            .I(N__4299));
    LocalMux I__821 (
            .O(N__4299),
            .I(N__4296));
    Span4Mux_v I__820 (
            .O(N__4296),
            .I(N__4293));
    Odrv4 I__819 (
            .O(N__4293),
            .I(CIA_ENABLEm));
    InMux I__818 (
            .O(N__4290),
            .I(N__4285));
    InMux I__817 (
            .O(N__4289),
            .I(N__4280));
    InMux I__816 (
            .O(N__4288),
            .I(N__4280));
    LocalMux I__815 (
            .O(N__4285),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    LocalMux I__814 (
            .O(N__4280),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    InMux I__813 (
            .O(N__4275),
            .I(N__4269));
    InMux I__812 (
            .O(N__4274),
            .I(N__4269));
    LocalMux I__811 (
            .O(N__4269),
            .I(N__4265));
    InMux I__810 (
            .O(N__4268),
            .I(N__4262));
    Span4Mux_v I__809 (
            .O(N__4265),
            .I(N__4259));
    LocalMux I__808 (
            .O(N__4262),
            .I(N__4256));
    Sp12to4 I__807 (
            .O(N__4259),
            .I(N__4251));
    Span12Mux_h I__806 (
            .O(N__4256),
            .I(N__4251));
    Odrv12 I__805 (
            .O(N__4251),
            .I(\U409_CIA.g0Z0Z_14 ));
    CascadeMux I__804 (
            .O(N__4248),
            .I(N__4243));
    CascadeMux I__803 (
            .O(N__4247),
            .I(N__4240));
    CascadeMux I__802 (
            .O(N__4246),
            .I(N__4237));
    InMux I__801 (
            .O(N__4243),
            .I(N__4232));
    InMux I__800 (
            .O(N__4240),
            .I(N__4232));
    InMux I__799 (
            .O(N__4237),
            .I(N__4229));
    LocalMux I__798 (
            .O(N__4232),
            .I(N__4224));
    LocalMux I__797 (
            .O(N__4229),
            .I(N__4224));
    Span4Mux_v I__796 (
            .O(N__4224),
            .I(N__4221));
    Sp12to4 I__795 (
            .O(N__4221),
            .I(N__4218));
    Span12Mux_h I__794 (
            .O(N__4218),
            .I(N__4215));
    Odrv12 I__793 (
            .O(N__4215),
            .I(\U409_CIA.g0Z0Z_13 ));
    InMux I__792 (
            .O(N__4212),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    CascadeMux I__791 (
            .O(N__4209),
            .I(N__4206));
    InMux I__790 (
            .O(N__4206),
            .I(N__4202));
    InMux I__789 (
            .O(N__4205),
            .I(N__4199));
    LocalMux I__788 (
            .O(N__4202),
            .I(N__4196));
    LocalMux I__787 (
            .O(N__4199),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    Odrv4 I__786 (
            .O(N__4196),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    InMux I__785 (
            .O(N__4191),
            .I(N__4188));
    LocalMux I__784 (
            .O(N__4188),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__783 (
            .O(N__4185),
            .I(N__4182));
    LocalMux I__782 (
            .O(N__4182),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    CascadeMux I__781 (
            .O(N__4179),
            .I(N__4176));
    InMux I__780 (
            .O(N__4176),
            .I(N__4173));
    LocalMux I__779 (
            .O(N__4173),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__778 (
            .O(N__4170),
            .I(N__4166));
    InMux I__777 (
            .O(N__4169),
            .I(N__4163));
    LocalMux I__776 (
            .O(N__4166),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__775 (
            .O(N__4163),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__774 (
            .O(N__4158),
            .I(N__4154));
    InMux I__773 (
            .O(N__4157),
            .I(N__4151));
    LocalMux I__772 (
            .O(N__4154),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__771 (
            .O(N__4151),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    CascadeMux I__770 (
            .O(N__4146),
            .I(N__4142));
    CascadeMux I__769 (
            .O(N__4145),
            .I(N__4139));
    InMux I__768 (
            .O(N__4142),
            .I(N__4133));
    InMux I__767 (
            .O(N__4139),
            .I(N__4133));
    InMux I__766 (
            .O(N__4138),
            .I(N__4130));
    LocalMux I__765 (
            .O(N__4133),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__764 (
            .O(N__4130),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    InMux I__763 (
            .O(N__4125),
            .I(N__4121));
    InMux I__762 (
            .O(N__4124),
            .I(N__4118));
    LocalMux I__761 (
            .O(N__4121),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__760 (
            .O(N__4118),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    InMux I__759 (
            .O(N__4113),
            .I(N__4109));
    InMux I__758 (
            .O(N__4112),
            .I(N__4106));
    LocalMux I__757 (
            .O(N__4109),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__756 (
            .O(N__4106),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    CascadeMux I__755 (
            .O(N__4101),
            .I(N__4097));
    InMux I__754 (
            .O(N__4100),
            .I(N__4094));
    InMux I__753 (
            .O(N__4097),
            .I(N__4091));
    LocalMux I__752 (
            .O(N__4094),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__751 (
            .O(N__4091),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    CascadeMux I__750 (
            .O(N__4086),
            .I(N__4082));
    CascadeMux I__749 (
            .O(N__4085),
            .I(N__4077));
    InMux I__748 (
            .O(N__4082),
            .I(N__4072));
    InMux I__747 (
            .O(N__4081),
            .I(N__4072));
    InMux I__746 (
            .O(N__4080),
            .I(N__4069));
    InMux I__745 (
            .O(N__4077),
            .I(N__4066));
    LocalMux I__744 (
            .O(N__4072),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__743 (
            .O(N__4069),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__742 (
            .O(N__4066),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__741 (
            .O(N__4059),
            .I(N__4056));
    LocalMux I__740 (
            .O(N__4056),
            .I(\U409_TICK.TICK603_11 ));
    InMux I__739 (
            .O(N__4053),
            .I(N__4049));
    InMux I__738 (
            .O(N__4052),
            .I(N__4046));
    LocalMux I__737 (
            .O(N__4049),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__736 (
            .O(N__4046),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    CascadeMux I__735 (
            .O(N__4041),
            .I(\U409_TICK.TICK603_8_cascade_ ));
    InMux I__734 (
            .O(N__4038),
            .I(N__4034));
    InMux I__733 (
            .O(N__4037),
            .I(N__4031));
    LocalMux I__732 (
            .O(N__4034),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__731 (
            .O(N__4031),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    InMux I__730 (
            .O(N__4026),
            .I(N__4013));
    InMux I__729 (
            .O(N__4025),
            .I(N__4013));
    InMux I__728 (
            .O(N__4024),
            .I(N__4013));
    InMux I__727 (
            .O(N__4023),
            .I(N__4004));
    InMux I__726 (
            .O(N__4022),
            .I(N__4004));
    InMux I__725 (
            .O(N__4021),
            .I(N__4004));
    InMux I__724 (
            .O(N__4020),
            .I(N__4004));
    LocalMux I__723 (
            .O(N__4013),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__722 (
            .O(N__4004),
            .I(\U409_TICK.TICK603_14 ));
    InMux I__721 (
            .O(N__3999),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__720 (
            .O(N__3996),
            .I(N__3992));
    InMux I__719 (
            .O(N__3995),
            .I(N__3989));
    LocalMux I__718 (
            .O(N__3992),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__717 (
            .O(N__3989),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__716 (
            .O(N__3984),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__715 (
            .O(N__3981),
            .I(bfn_11_7_0_));
    InMux I__714 (
            .O(N__3978),
            .I(N__3975));
    LocalMux I__713 (
            .O(N__3975),
            .I(N__3971));
    InMux I__712 (
            .O(N__3974),
            .I(N__3968));
    Odrv4 I__711 (
            .O(N__3971),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__710 (
            .O(N__3968),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    InMux I__709 (
            .O(N__3963),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__708 (
            .O(N__3960),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__707 (
            .O(N__3957),
            .I(N__3954));
    LocalMux I__706 (
            .O(N__3954),
            .I(N__3950));
    InMux I__705 (
            .O(N__3953),
            .I(N__3947));
    Odrv4 I__704 (
            .O(N__3950),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__703 (
            .O(N__3947),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    InMux I__702 (
            .O(N__3942),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__701 (
            .O(N__3939),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__700 (
            .O(N__3936),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__699 (
            .O(N__3933),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__698 (
            .O(N__3930),
            .I(N__3927));
    LocalMux I__697 (
            .O(N__3927),
            .I(\U409_TICK.TICK503_8 ));
    CascadeMux I__696 (
            .O(N__3924),
            .I(\U409_TICK.TICK503_11_cascade_ ));
    CascadeMux I__695 (
            .O(N__3921),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    IoInMux I__694 (
            .O(N__3918),
            .I(N__3915));
    LocalMux I__693 (
            .O(N__3915),
            .I(N__3912));
    Span12Mux_s10_v I__692 (
            .O(N__3912),
            .I(N__3908));
    InMux I__691 (
            .O(N__3911),
            .I(N__3905));
    Odrv12 I__690 (
            .O(N__3908),
            .I(TICK50_c));
    LocalMux I__689 (
            .O(N__3905),
            .I(TICK50_c));
    CascadeMux I__688 (
            .O(N__3900),
            .I(N__3897));
    InMux I__687 (
            .O(N__3897),
            .I(N__3890));
    InMux I__686 (
            .O(N__3896),
            .I(N__3890));
    InMux I__685 (
            .O(N__3895),
            .I(N__3887));
    LocalMux I__684 (
            .O(N__3890),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__683 (
            .O(N__3887),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    CascadeMux I__682 (
            .O(N__3882),
            .I(N__3878));
    CascadeMux I__681 (
            .O(N__3881),
            .I(N__3873));
    InMux I__680 (
            .O(N__3878),
            .I(N__3870));
    InMux I__679 (
            .O(N__3877),
            .I(N__3865));
    InMux I__678 (
            .O(N__3876),
            .I(N__3865));
    InMux I__677 (
            .O(N__3873),
            .I(N__3862));
    LocalMux I__676 (
            .O(N__3870),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__675 (
            .O(N__3865),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__674 (
            .O(N__3862),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__673 (
            .O(N__3855),
            .I(N__3851));
    InMux I__672 (
            .O(N__3854),
            .I(N__3848));
    LocalMux I__671 (
            .O(N__3851),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__670 (
            .O(N__3848),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__669 (
            .O(N__3843),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__668 (
            .O(N__3840),
            .I(N__3836));
    InMux I__667 (
            .O(N__3839),
            .I(N__3833));
    LocalMux I__666 (
            .O(N__3836),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__665 (
            .O(N__3833),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__664 (
            .O(N__3828),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    InMux I__663 (
            .O(N__3825),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__662 (
            .O(N__3822),
            .I(N__3818));
    InMux I__661 (
            .O(N__3821),
            .I(N__3815));
    LocalMux I__660 (
            .O(N__3818),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__659 (
            .O(N__3815),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__658 (
            .O(N__3810),
            .I(N__3807));
    LocalMux I__657 (
            .O(N__3807),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__656 (
            .O(N__3804),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    CascadeMux I__655 (
            .O(N__3801),
            .I(N__3798));
    InMux I__654 (
            .O(N__3798),
            .I(N__3795));
    LocalMux I__653 (
            .O(N__3795),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__652 (
            .O(N__3792),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__651 (
            .O(N__3789),
            .I(N__3786));
    LocalMux I__650 (
            .O(N__3786),
            .I(N__3783));
    Span4Mux_v I__649 (
            .O(N__3783),
            .I(N__3780));
    Sp12to4 I__648 (
            .O(N__3780),
            .I(N__3777));
    Span12Mux_h I__647 (
            .O(N__3777),
            .I(N__3774));
    Odrv12 I__646 (
            .O(N__3774),
            .I(TACKn_in));
    IoInMux I__645 (
            .O(N__3771),
            .I(N__3768));
    LocalMux I__644 (
            .O(N__3768),
            .I(N__3765));
    Span4Mux_s1_v I__643 (
            .O(N__3765),
            .I(N__3762));
    Sp12to4 I__642 (
            .O(N__3762),
            .I(N__3758));
    InMux I__641 (
            .O(N__3761),
            .I(N__3755));
    Span12Mux_s11_h I__640 (
            .O(N__3758),
            .I(N__3752));
    LocalMux I__639 (
            .O(N__3755),
            .I(N__3749));
    Span12Mux_v I__638 (
            .O(N__3752),
            .I(N__3746));
    Span4Mux_v I__637 (
            .O(N__3749),
            .I(N__3743));
    Odrv12 I__636 (
            .O(N__3746),
            .I(BUFENn_c));
    Odrv4 I__635 (
            .O(N__3743),
            .I(BUFENn_c));
    InMux I__634 (
            .O(N__3738),
            .I(N__3735));
    LocalMux I__633 (
            .O(N__3735),
            .I(N__3732));
    Span4Mux_v I__632 (
            .O(N__3732),
            .I(N__3729));
    Sp12to4 I__631 (
            .O(N__3729),
            .I(N__3726));
    Span12Mux_h I__630 (
            .O(N__3726),
            .I(N__3723));
    Odrv12 I__629 (
            .O(N__3723),
            .I(A_c_13));
    IoInMux I__628 (
            .O(N__3720),
            .I(N__3717));
    LocalMux I__627 (
            .O(N__3717),
            .I(N__3714));
    Span4Mux_s1_h I__626 (
            .O(N__3714),
            .I(N__3711));
    Sp12to4 I__625 (
            .O(N__3711),
            .I(N__3708));
    Span12Mux_s9_v I__624 (
            .O(N__3708),
            .I(N__3705));
    Span12Mux_h I__623 (
            .O(N__3705),
            .I(N__3702));
    Odrv12 I__622 (
            .O(N__3702),
            .I(U409_ADDRESS_DECODE_un1_CIACS1n_i));
    InMux I__621 (
            .O(N__3699),
            .I(N__3696));
    LocalMux I__620 (
            .O(N__3696),
            .I(N__3693));
    Span4Mux_v I__619 (
            .O(N__3693),
            .I(N__3690));
    Sp12to4 I__618 (
            .O(N__3690),
            .I(N__3687));
    Span12Mux_h I__617 (
            .O(N__3687),
            .I(N__3684));
    Odrv12 I__616 (
            .O(N__3684),
            .I(A_c_12));
    IoInMux I__615 (
            .O(N__3681),
            .I(N__3678));
    LocalMux I__614 (
            .O(N__3678),
            .I(N__3675));
    IoSpan4Mux I__613 (
            .O(N__3675),
            .I(N__3672));
    Span4Mux_s3_h I__612 (
            .O(N__3672),
            .I(N__3669));
    Sp12to4 I__611 (
            .O(N__3669),
            .I(N__3666));
    Span12Mux_h I__610 (
            .O(N__3666),
            .I(N__3663));
    Odrv12 I__609 (
            .O(N__3663),
            .I(U409_ADDRESS_DECODE_un1_CIACS0n_i));
    CascadeMux I__608 (
            .O(N__3660),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    CascadeMux I__607 (
            .O(N__3657),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ));
    CascadeMux I__606 (
            .O(N__3654),
            .I(N__3651));
    InMux I__605 (
            .O(N__3651),
            .I(N__3647));
    InMux I__604 (
            .O(N__3650),
            .I(N__3644));
    LocalMux I__603 (
            .O(N__3647),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5 ));
    LocalMux I__602 (
            .O(N__3644),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5 ));
    InMux I__601 (
            .O(N__3639),
            .I(N__3634));
    InMux I__600 (
            .O(N__3638),
            .I(N__3631));
    InMux I__599 (
            .O(N__3637),
            .I(N__3628));
    LocalMux I__598 (
            .O(N__3634),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__597 (
            .O(N__3631),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__596 (
            .O(N__3628),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    CascadeMux I__595 (
            .O(N__3621),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_ ));
    InMux I__594 (
            .O(N__3618),
            .I(N__3615));
    LocalMux I__593 (
            .O(N__3615),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_11 ));
    InMux I__592 (
            .O(N__3612),
            .I(N__3605));
    InMux I__591 (
            .O(N__3611),
            .I(N__3605));
    InMux I__590 (
            .O(N__3610),
            .I(N__3602));
    LocalMux I__589 (
            .O(N__3605),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__588 (
            .O(N__3602),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    CascadeMux I__587 (
            .O(N__3597),
            .I(N__3592));
    InMux I__586 (
            .O(N__3596),
            .I(N__3586));
    InMux I__585 (
            .O(N__3595),
            .I(N__3586));
    InMux I__584 (
            .O(N__3592),
            .I(N__3581));
    InMux I__583 (
            .O(N__3591),
            .I(N__3581));
    LocalMux I__582 (
            .O(N__3586),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__581 (
            .O(N__3581),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    InMux I__580 (
            .O(N__3576),
            .I(N__3567));
    InMux I__579 (
            .O(N__3575),
            .I(N__3567));
    InMux I__578 (
            .O(N__3574),
            .I(N__3564));
    InMux I__577 (
            .O(N__3573),
            .I(N__3559));
    InMux I__576 (
            .O(N__3572),
            .I(N__3559));
    LocalMux I__575 (
            .O(N__3567),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__574 (
            .O(N__3564),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__573 (
            .O(N__3559),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    CascadeMux I__572 (
            .O(N__3552),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_2_cascade_ ));
    InMux I__571 (
            .O(N__3549),
            .I(N__3546));
    LocalMux I__570 (
            .O(N__3546),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1 ));
    InMux I__569 (
            .O(N__3543),
            .I(N__3535));
    InMux I__568 (
            .O(N__3542),
            .I(N__3530));
    InMux I__567 (
            .O(N__3541),
            .I(N__3530));
    InMux I__566 (
            .O(N__3540),
            .I(N__3527));
    InMux I__565 (
            .O(N__3539),
            .I(N__3522));
    InMux I__564 (
            .O(N__3538),
            .I(N__3522));
    LocalMux I__563 (
            .O(N__3535),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__562 (
            .O(N__3530),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__561 (
            .O(N__3527),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__560 (
            .O(N__3522),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    InMux I__559 (
            .O(N__3513),
            .I(N__3507));
    InMux I__558 (
            .O(N__3512),
            .I(N__3504));
    InMux I__557 (
            .O(N__3511),
            .I(N__3499));
    InMux I__556 (
            .O(N__3510),
            .I(N__3499));
    LocalMux I__555 (
            .O(N__3507),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__554 (
            .O(N__3504),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__553 (
            .O(N__3499),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    InMux I__552 (
            .O(N__3492),
            .I(N__3489));
    LocalMux I__551 (
            .O(N__3489),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_5 ));
    InMux I__550 (
            .O(N__3486),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__549 (
            .O(N__3483),
            .I(N__3480));
    LocalMux I__548 (
            .O(N__3480),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    CascadeMux I__547 (
            .O(N__3477),
            .I(N__3474));
    InMux I__546 (
            .O(N__3474),
            .I(N__3471));
    LocalMux I__545 (
            .O(N__3471),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    CascadeMux I__544 (
            .O(N__3468),
            .I(N__3465));
    InMux I__543 (
            .O(N__3465),
            .I(N__3462));
    LocalMux I__542 (
            .O(N__3462),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    CascadeMux I__541 (
            .O(N__3459),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_ ));
    CascadeMux I__540 (
            .O(N__3456),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_cascade_ ));
    InMux I__539 (
            .O(N__3453),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__538 (
            .O(N__3450),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__537 (
            .O(N__3447),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__536 (
            .O(N__3444),
            .I(bfn_10_9_0_));
    InMux I__535 (
            .O(N__3441),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__534 (
            .O(N__3438),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__533 (
            .O(N__3435),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__532 (
            .O(N__3432),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__531 (
            .O(N__3429),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__530 (
            .O(N__3426),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__529 (
            .O(N__3423),
            .I(N__3414));
    InMux I__528 (
            .O(N__3422),
            .I(N__3414));
    InMux I__527 (
            .O(N__3421),
            .I(N__3414));
    LocalMux I__526 (
            .O(N__3414),
            .I(N__3411));
    Odrv12 I__525 (
            .O(N__3411),
            .I(U409_ADDRESS_DECODE_un5_RAMSPACEn));
    InMux I__524 (
            .O(N__3408),
            .I(N__3398));
    InMux I__523 (
            .O(N__3407),
            .I(N__3398));
    InMux I__522 (
            .O(N__3406),
            .I(N__3398));
    InMux I__521 (
            .O(N__3405),
            .I(N__3395));
    LocalMux I__520 (
            .O(N__3398),
            .I(N__3392));
    LocalMux I__519 (
            .O(N__3395),
            .I(N__3389));
    Span4Mux_v I__518 (
            .O(N__3392),
            .I(N__3385));
    Span4Mux_v I__517 (
            .O(N__3389),
            .I(N__3382));
    InMux I__516 (
            .O(N__3388),
            .I(N__3379));
    Sp12to4 I__515 (
            .O(N__3385),
            .I(N__3371));
    Sp12to4 I__514 (
            .O(N__3382),
            .I(N__3371));
    LocalMux I__513 (
            .O(N__3379),
            .I(N__3371));
    CascadeMux I__512 (
            .O(N__3378),
            .I(N__3368));
    Span12Mux_h I__511 (
            .O(N__3371),
            .I(N__3365));
    InMux I__510 (
            .O(N__3368),
            .I(N__3362));
    Odrv12 I__509 (
            .O(N__3365),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    LocalMux I__508 (
            .O(N__3362),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    CascadeMux I__507 (
            .O(N__3357),
            .I(N__3354));
    InMux I__506 (
            .O(N__3354),
            .I(N__3351));
    LocalMux I__505 (
            .O(N__3351),
            .I(N__3348));
    Span4Mux_h I__504 (
            .O(N__3348),
            .I(N__3345));
    Odrv4 I__503 (
            .O(N__3345),
            .I(U409_ADDRESS_DECODE_HIROM));
    CascadeMux I__502 (
            .O(N__3342),
            .I(N__3338));
    InMux I__501 (
            .O(N__3341),
            .I(N__3330));
    InMux I__500 (
            .O(N__3338),
            .I(N__3330));
    InMux I__499 (
            .O(N__3337),
            .I(N__3330));
    LocalMux I__498 (
            .O(N__3330),
            .I(N__3327));
    Span4Mux_v I__497 (
            .O(N__3327),
            .I(N__3324));
    Sp12to4 I__496 (
            .O(N__3324),
            .I(N__3321));
    Span12Mux_h I__495 (
            .O(N__3321),
            .I(N__3318));
    Span12Mux_v I__494 (
            .O(N__3318),
            .I(N__3315));
    Odrv12 I__493 (
            .O(N__3315),
            .I(OVL_c));
    InMux I__492 (
            .O(N__3312),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__491 (
            .O(N__3309),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__490 (
            .O(N__3306),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__489 (
            .O(N__3303),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    CascadeMux I__488 (
            .O(N__3300),
            .I(N__3296));
    InMux I__487 (
            .O(N__3299),
            .I(N__3293));
    InMux I__486 (
            .O(N__3296),
            .I(N__3290));
    LocalMux I__485 (
            .O(N__3293),
            .I(N__3286));
    LocalMux I__484 (
            .O(N__3290),
            .I(N__3283));
    InMux I__483 (
            .O(N__3289),
            .I(N__3280));
    Odrv4 I__482 (
            .O(N__3286),
            .I(CIA_SPACEm_3));
    Odrv4 I__481 (
            .O(N__3283),
            .I(CIA_SPACEm_3));
    LocalMux I__480 (
            .O(N__3280),
            .I(CIA_SPACEm_3));
    CascadeMux I__479 (
            .O(N__3273),
            .I(N__3266));
    CascadeMux I__478 (
            .O(N__3272),
            .I(N__3263));
    CascadeMux I__477 (
            .O(N__3271),
            .I(N__3259));
    InMux I__476 (
            .O(N__3270),
            .I(N__3256));
    InMux I__475 (
            .O(N__3269),
            .I(N__3249));
    InMux I__474 (
            .O(N__3266),
            .I(N__3249));
    InMux I__473 (
            .O(N__3263),
            .I(N__3249));
    InMux I__472 (
            .O(N__3262),
            .I(N__3246));
    InMux I__471 (
            .O(N__3259),
            .I(N__3243));
    LocalMux I__470 (
            .O(N__3256),
            .I(N__3240));
    LocalMux I__469 (
            .O(N__3249),
            .I(N__3231));
    LocalMux I__468 (
            .O(N__3246),
            .I(N__3231));
    LocalMux I__467 (
            .O(N__3243),
            .I(N__3231));
    Sp12to4 I__466 (
            .O(N__3240),
            .I(N__3231));
    Span12Mux_v I__465 (
            .O(N__3231),
            .I(N__3228));
    Odrv12 I__464 (
            .O(N__3228),
            .I(A_c_22));
    InMux I__463 (
            .O(N__3225),
            .I(N__3221));
    InMux I__462 (
            .O(N__3224),
            .I(N__3217));
    LocalMux I__461 (
            .O(N__3221),
            .I(N__3214));
    InMux I__460 (
            .O(N__3220),
            .I(N__3211));
    LocalMux I__459 (
            .O(N__3217),
            .I(N__3208));
    Span4Mux_v I__458 (
            .O(N__3214),
            .I(N__3203));
    LocalMux I__457 (
            .O(N__3211),
            .I(N__3203));
    Odrv12 I__456 (
            .O(N__3208),
            .I(CIA_SPACEm_6));
    Odrv4 I__455 (
            .O(N__3203),
            .I(CIA_SPACEm_6));
    InMux I__454 (
            .O(N__3198),
            .I(N__3195));
    LocalMux I__453 (
            .O(N__3195),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_8 ));
    InMux I__452 (
            .O(N__3192),
            .I(N__3189));
    LocalMux I__451 (
            .O(N__3189),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_9 ));
    CascadeMux I__450 (
            .O(N__3186),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_10_cascade_ ));
    InMux I__449 (
            .O(N__3183),
            .I(N__3180));
    LocalMux I__448 (
            .O(N__3180),
            .I(N__3177));
    Span4Mux_h I__447 (
            .O(N__3177),
            .I(N__3174));
    Sp12to4 I__446 (
            .O(N__3174),
            .I(N__3171));
    Odrv12 I__445 (
            .O(N__3171),
            .I(TT_c_1));
    CascadeMux I__444 (
            .O(N__3168),
            .I(N__3165));
    InMux I__443 (
            .O(N__3165),
            .I(N__3160));
    InMux I__442 (
            .O(N__3164),
            .I(N__3157));
    InMux I__441 (
            .O(N__3163),
            .I(N__3154));
    LocalMux I__440 (
            .O(N__3160),
            .I(N__3151));
    LocalMux I__439 (
            .O(N__3157),
            .I(N__3146));
    LocalMux I__438 (
            .O(N__3154),
            .I(N__3146));
    Span4Mux_v I__437 (
            .O(N__3151),
            .I(N__3143));
    Span4Mux_v I__436 (
            .O(N__3146),
            .I(N__3140));
    Sp12to4 I__435 (
            .O(N__3143),
            .I(N__3137));
    Span4Mux_h I__434 (
            .O(N__3140),
            .I(N__3134));
    Odrv12 I__433 (
            .O(N__3137),
            .I(A_c_31));
    Odrv4 I__432 (
            .O(N__3134),
            .I(A_c_31));
    InMux I__431 (
            .O(N__3129),
            .I(N__3126));
    LocalMux I__430 (
            .O(N__3126),
            .I(N__3123));
    Span12Mux_h I__429 (
            .O(N__3123),
            .I(N__3120));
    Odrv12 I__428 (
            .O(N__3120),
            .I(TT_c_0));
    InMux I__427 (
            .O(N__3117),
            .I(N__3114));
    LocalMux I__426 (
            .O(N__3114),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_11 ));
    InMux I__425 (
            .O(N__3111),
            .I(N__3108));
    LocalMux I__424 (
            .O(N__3108),
            .I(N__3104));
    InMux I__423 (
            .O(N__3107),
            .I(N__3101));
    Span4Mux_v I__422 (
            .O(N__3104),
            .I(N__3098));
    LocalMux I__421 (
            .O(N__3101),
            .I(N__3095));
    Odrv4 I__420 (
            .O(N__3098),
            .I(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3 ));
    Odrv12 I__419 (
            .O(N__3095),
            .I(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3 ));
    IoInMux I__418 (
            .O(N__3090),
            .I(N__3087));
    LocalMux I__417 (
            .O(N__3087),
            .I(N__3084));
    Span4Mux_s0_v I__416 (
            .O(N__3084),
            .I(N__3081));
    Sp12to4 I__415 (
            .O(N__3081),
            .I(N__3078));
    Span12Mux_s11_h I__414 (
            .O(N__3078),
            .I(N__3075));
    Span12Mux_v I__413 (
            .O(N__3075),
            .I(N__3072));
    Odrv12 I__412 (
            .O(N__3072),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn_i));
    InMux I__411 (
            .O(N__3069),
            .I(N__3066));
    LocalMux I__410 (
            .O(N__3066),
            .I(N__3063));
    Odrv12 I__409 (
            .O(N__3063),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ));
    InMux I__408 (
            .O(N__3060),
            .I(N__3055));
    InMux I__407 (
            .O(N__3059),
            .I(N__3049));
    InMux I__406 (
            .O(N__3058),
            .I(N__3046));
    LocalMux I__405 (
            .O(N__3055),
            .I(N__3043));
    InMux I__404 (
            .O(N__3054),
            .I(N__3040));
    InMux I__403 (
            .O(N__3053),
            .I(N__3035));
    InMux I__402 (
            .O(N__3052),
            .I(N__3035));
    LocalMux I__401 (
            .O(N__3049),
            .I(N__3032));
    LocalMux I__400 (
            .O(N__3046),
            .I(N__3029));
    Span4Mux_v I__399 (
            .O(N__3043),
            .I(N__3023));
    LocalMux I__398 (
            .O(N__3040),
            .I(N__3023));
    LocalMux I__397 (
            .O(N__3035),
            .I(N__3020));
    Span4Mux_v I__396 (
            .O(N__3032),
            .I(N__3015));
    Span4Mux_v I__395 (
            .O(N__3029),
            .I(N__3015));
    InMux I__394 (
            .O(N__3028),
            .I(N__3012));
    Span4Mux_v I__393 (
            .O(N__3023),
            .I(N__3007));
    Span4Mux_v I__392 (
            .O(N__3020),
            .I(N__3007));
    Sp12to4 I__391 (
            .O(N__3015),
            .I(N__3000));
    LocalMux I__390 (
            .O(N__3012),
            .I(N__3000));
    Sp12to4 I__389 (
            .O(N__3007),
            .I(N__3000));
    Odrv12 I__388 (
            .O(N__3000),
            .I(A_c_23));
    IoInMux I__387 (
            .O(N__2997),
            .I(N__2994));
    LocalMux I__386 (
            .O(N__2994),
            .I(N__2991));
    Span12Mux_s11_v I__385 (
            .O(N__2991),
            .I(N__2988));
    Odrv12 I__384 (
            .O(N__2988),
            .I(PORTSIZE_0_i));
    CascadeMux I__383 (
            .O(N__2985),
            .I(N__2981));
    CascadeMux I__382 (
            .O(N__2984),
            .I(N__2978));
    InMux I__381 (
            .O(N__2981),
            .I(N__2975));
    InMux I__380 (
            .O(N__2978),
            .I(N__2972));
    LocalMux I__379 (
            .O(N__2975),
            .I(N__2969));
    LocalMux I__378 (
            .O(N__2972),
            .I(N__2966));
    Odrv12 I__377 (
            .O(N__2969),
            .I(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0 ));
    Odrv4 I__376 (
            .O(N__2966),
            .I(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0 ));
    IoInMux I__375 (
            .O(N__2961),
            .I(N__2958));
    LocalMux I__374 (
            .O(N__2958),
            .I(N__2955));
    IoSpan4Mux I__373 (
            .O(N__2955),
            .I(N__2952));
    Sp12to4 I__372 (
            .O(N__2952),
            .I(N__2949));
    Span12Mux_s7_v I__371 (
            .O(N__2949),
            .I(N__2946));
    Odrv12 I__370 (
            .O(N__2946),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn_i));
    InMux I__369 (
            .O(N__2943),
            .I(N__2937));
    InMux I__368 (
            .O(N__2942),
            .I(N__2937));
    LocalMux I__367 (
            .O(N__2937),
            .I(N__2933));
    InMux I__366 (
            .O(N__2936),
            .I(N__2930));
    Span4Mux_h I__365 (
            .O(N__2933),
            .I(N__2925));
    LocalMux I__364 (
            .O(N__2930),
            .I(N__2925));
    Span4Mux_v I__363 (
            .O(N__2925),
            .I(N__2922));
    Span4Mux_v I__362 (
            .O(N__2922),
            .I(N__2919));
    Span4Mux_h I__361 (
            .O(N__2919),
            .I(N__2916));
    Odrv4 I__360 (
            .O(N__2916),
            .I(A_c_28));
    CascadeMux I__359 (
            .O(N__2913),
            .I(\U409_CIA.g0Z0Z_2_cascade_ ));
    CascadeMux I__358 (
            .O(N__2910),
            .I(N__2906));
    InMux I__357 (
            .O(N__2909),
            .I(N__2900));
    InMux I__356 (
            .O(N__2906),
            .I(N__2900));
    InMux I__355 (
            .O(N__2905),
            .I(N__2897));
    LocalMux I__354 (
            .O(N__2900),
            .I(N__2892));
    LocalMux I__353 (
            .O(N__2897),
            .I(N__2892));
    Span4Mux_v I__352 (
            .O(N__2892),
            .I(N__2889));
    Span4Mux_v I__351 (
            .O(N__2889),
            .I(N__2886));
    Sp12to4 I__350 (
            .O(N__2886),
            .I(N__2883));
    Odrv12 I__349 (
            .O(N__2883),
            .I(A_c_26));
    InMux I__348 (
            .O(N__2880),
            .I(N__2877));
    LocalMux I__347 (
            .O(N__2877),
            .I(N__2873));
    CascadeMux I__346 (
            .O(N__2876),
            .I(N__2870));
    Span4Mux_v I__345 (
            .O(N__2873),
            .I(N__2866));
    InMux I__344 (
            .O(N__2870),
            .I(N__2861));
    InMux I__343 (
            .O(N__2869),
            .I(N__2861));
    Sp12to4 I__342 (
            .O(N__2866),
            .I(N__2856));
    LocalMux I__341 (
            .O(N__2861),
            .I(N__2856));
    Odrv12 I__340 (
            .O(N__2856),
            .I(A_c_27));
    InMux I__339 (
            .O(N__2853),
            .I(N__2846));
    InMux I__338 (
            .O(N__2852),
            .I(N__2846));
    CascadeMux I__337 (
            .O(N__2851),
            .I(N__2843));
    LocalMux I__336 (
            .O(N__2846),
            .I(N__2840));
    InMux I__335 (
            .O(N__2843),
            .I(N__2837));
    Span4Mux_v I__334 (
            .O(N__2840),
            .I(N__2832));
    LocalMux I__333 (
            .O(N__2837),
            .I(N__2832));
    Span4Mux_h I__332 (
            .O(N__2832),
            .I(N__2829));
    Span4Mux_v I__331 (
            .O(N__2829),
            .I(N__2826));
    Odrv4 I__330 (
            .O(N__2826),
            .I(A_c_24));
    InMux I__329 (
            .O(N__2823),
            .I(N__2820));
    LocalMux I__328 (
            .O(N__2820),
            .I(\U409_CIA.g0Z0Z_10 ));
    CascadeMux I__327 (
            .O(N__2817),
            .I(\U409_CIA.g0Z0Z_8_cascade_ ));
    CascadeMux I__326 (
            .O(N__2814),
            .I(N__2810));
    InMux I__325 (
            .O(N__2813),
            .I(N__2805));
    InMux I__324 (
            .O(N__2810),
            .I(N__2805));
    LocalMux I__323 (
            .O(N__2805),
            .I(N__2802));
    Span12Mux_s7_h I__322 (
            .O(N__2802),
            .I(N__2799));
    Span12Mux_v I__321 (
            .O(N__2799),
            .I(N__2796));
    Odrv12 I__320 (
            .O(N__2796),
            .I(A_c_16));
    InMux I__319 (
            .O(N__2793),
            .I(N__2787));
    InMux I__318 (
            .O(N__2792),
            .I(N__2787));
    LocalMux I__317 (
            .O(N__2787),
            .I(N__2784));
    Span4Mux_v I__316 (
            .O(N__2784),
            .I(N__2781));
    Sp12to4 I__315 (
            .O(N__2781),
            .I(N__2778));
    Span12Mux_v I__314 (
            .O(N__2778),
            .I(N__2775));
    Odrv12 I__313 (
            .O(N__2775),
            .I(A_c_17));
    InMux I__312 (
            .O(N__2772),
            .I(N__2769));
    LocalMux I__311 (
            .O(N__2769),
            .I(N__2766));
    Span4Mux_h I__310 (
            .O(N__2766),
            .I(N__2761));
    InMux I__309 (
            .O(N__2765),
            .I(N__2758));
    InMux I__308 (
            .O(N__2764),
            .I(N__2755));
    Span4Mux_v I__307 (
            .O(N__2761),
            .I(N__2752));
    LocalMux I__306 (
            .O(N__2758),
            .I(N__2747));
    LocalMux I__305 (
            .O(N__2755),
            .I(N__2747));
    Odrv4 I__304 (
            .O(N__2752),
            .I(A_c_25));
    Odrv12 I__303 (
            .O(N__2747),
            .I(A_c_25));
    CascadeMux I__302 (
            .O(N__2742),
            .I(N__2739));
    InMux I__301 (
            .O(N__2739),
            .I(N__2735));
    InMux I__300 (
            .O(N__2738),
            .I(N__2732));
    LocalMux I__299 (
            .O(N__2735),
            .I(N__2727));
    LocalMux I__298 (
            .O(N__2732),
            .I(N__2727));
    Span4Mux_v I__297 (
            .O(N__2727),
            .I(N__2724));
    Sp12to4 I__296 (
            .O(N__2724),
            .I(N__2721));
    Span12Mux_h I__295 (
            .O(N__2721),
            .I(N__2718));
    Span12Mux_v I__294 (
            .O(N__2718),
            .I(N__2715));
    Odrv12 I__293 (
            .O(N__2715),
            .I(A_c_18));
    InMux I__292 (
            .O(N__2712),
            .I(N__2709));
    LocalMux I__291 (
            .O(N__2709),
            .I(\U409_CIA.g0Z0Z_11 ));
    InMux I__290 (
            .O(N__2706),
            .I(N__2703));
    LocalMux I__289 (
            .O(N__2703),
            .I(N__2698));
    InMux I__288 (
            .O(N__2702),
            .I(N__2693));
    InMux I__287 (
            .O(N__2701),
            .I(N__2693));
    Span4Mux_h I__286 (
            .O(N__2698),
            .I(N__2690));
    LocalMux I__285 (
            .O(N__2693),
            .I(N__2687));
    Span4Mux_v I__284 (
            .O(N__2690),
            .I(N__2684));
    Span4Mux_h I__283 (
            .O(N__2687),
            .I(N__2681));
    Sp12to4 I__282 (
            .O(N__2684),
            .I(N__2676));
    Sp12to4 I__281 (
            .O(N__2681),
            .I(N__2676));
    Span12Mux_v I__280 (
            .O(N__2676),
            .I(N__2673));
    Odrv12 I__279 (
            .O(N__2673),
            .I(A_c_19));
    InMux I__278 (
            .O(N__2670),
            .I(N__2666));
    InMux I__277 (
            .O(N__2669),
            .I(N__2663));
    LocalMux I__276 (
            .O(N__2666),
            .I(N__2660));
    LocalMux I__275 (
            .O(N__2663),
            .I(N__2656));
    Span4Mux_v I__274 (
            .O(N__2660),
            .I(N__2653));
    InMux I__273 (
            .O(N__2659),
            .I(N__2650));
    Span12Mux_v I__272 (
            .O(N__2656),
            .I(N__2647));
    Sp12to4 I__271 (
            .O(N__2653),
            .I(N__2642));
    LocalMux I__270 (
            .O(N__2650),
            .I(N__2642));
    Odrv12 I__269 (
            .O(N__2647),
            .I(A_c_20));
    Odrv12 I__268 (
            .O(N__2642),
            .I(A_c_20));
    InMux I__267 (
            .O(N__2637),
            .I(N__2631));
    InMux I__266 (
            .O(N__2636),
            .I(N__2626));
    InMux I__265 (
            .O(N__2635),
            .I(N__2626));
    InMux I__264 (
            .O(N__2634),
            .I(N__2623));
    LocalMux I__263 (
            .O(N__2631),
            .I(N__2616));
    LocalMux I__262 (
            .O(N__2626),
            .I(N__2616));
    LocalMux I__261 (
            .O(N__2623),
            .I(N__2616));
    Span4Mux_v I__260 (
            .O(N__2616),
            .I(N__2613));
    Span4Mux_h I__259 (
            .O(N__2613),
            .I(N__2610));
    Odrv4 I__258 (
            .O(N__2610),
            .I(A_c_21));
    CascadeMux I__257 (
            .O(N__2607),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_ ));
    InMux I__256 (
            .O(N__2604),
            .I(N__2601));
    LocalMux I__255 (
            .O(N__2601),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3 ));
    InMux I__254 (
            .O(N__2598),
            .I(N__2591));
    InMux I__253 (
            .O(N__2597),
            .I(N__2591));
    InMux I__252 (
            .O(N__2596),
            .I(N__2588));
    LocalMux I__251 (
            .O(N__2591),
            .I(N__2585));
    LocalMux I__250 (
            .O(N__2588),
            .I(N__2582));
    Span4Mux_v I__249 (
            .O(N__2585),
            .I(N__2577));
    Span4Mux_v I__248 (
            .O(N__2582),
            .I(N__2577));
    Sp12to4 I__247 (
            .O(N__2577),
            .I(N__2574));
    Odrv12 I__246 (
            .O(N__2574),
            .I(A_c_30));
    InMux I__245 (
            .O(N__2571),
            .I(N__2565));
    InMux I__244 (
            .O(N__2570),
            .I(N__2565));
    LocalMux I__243 (
            .O(N__2565),
            .I(N__2561));
    InMux I__242 (
            .O(N__2564),
            .I(N__2558));
    Span4Mux_v I__241 (
            .O(N__2561),
            .I(N__2553));
    LocalMux I__240 (
            .O(N__2558),
            .I(N__2553));
    Span4Mux_h I__239 (
            .O(N__2553),
            .I(N__2550));
    Span4Mux_v I__238 (
            .O(N__2550),
            .I(N__2547));
    Odrv4 I__237 (
            .O(N__2547),
            .I(A_c_29));
    ClkMux I__236 (
            .O(N__2544),
            .I(N__2499));
    ClkMux I__235 (
            .O(N__2543),
            .I(N__2499));
    ClkMux I__234 (
            .O(N__2542),
            .I(N__2499));
    ClkMux I__233 (
            .O(N__2541),
            .I(N__2499));
    ClkMux I__232 (
            .O(N__2540),
            .I(N__2499));
    ClkMux I__231 (
            .O(N__2539),
            .I(N__2499));
    ClkMux I__230 (
            .O(N__2538),
            .I(N__2499));
    ClkMux I__229 (
            .O(N__2537),
            .I(N__2499));
    ClkMux I__228 (
            .O(N__2536),
            .I(N__2499));
    ClkMux I__227 (
            .O(N__2535),
            .I(N__2499));
    ClkMux I__226 (
            .O(N__2534),
            .I(N__2499));
    ClkMux I__225 (
            .O(N__2533),
            .I(N__2499));
    ClkMux I__224 (
            .O(N__2532),
            .I(N__2499));
    ClkMux I__223 (
            .O(N__2531),
            .I(N__2499));
    ClkMux I__222 (
            .O(N__2530),
            .I(N__2499));
    GlobalMux I__221 (
            .O(N__2499),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.TACK_EN_iC  (
            .O(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .I(N__2543));
    INV \INVU409_TRANSFER_ACK.TACK_OUTnC  (
            .O(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .I(N__2541));
    INV \INVU409_TRANSFER_ACK.TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .I(N__2540));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .I(N__2537));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net ),
            .I(N__2535));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .I(N__2533));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .I(N__2531));
    INV \INVU409_TRANSFER_ACK.LASTCLK_0C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .I(N__2530));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .I(N__2539));
    INV \INVU409_TRANSFER_ACK.ROMENnC  (
            .O(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .I(N__2536));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .I(N__2534));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .I(N__2532));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .I(N__2538));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .I(N__2544));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .I(N__2542));
    defparam IN_MUX_bfv_10_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_8_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.HIROM_0_LC_1_13_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.HIROM_0_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.HIROM_0_LC_1_13_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.HIROM_0_LC_1_13_5  (
            .in0(N__2634),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2670),
            .lcout(CIA_SPACEm_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_9_LC_1_16_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_9_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_9_LC_1_16_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_9_LC_1_16_0  (
            .in0(N__2853),
            .in1(N__2765),
            .in2(N__3300),
            .in3(N__2909),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_1  (
            .in0(N__2869),
            .in1(N__2852),
            .in2(N__2910),
            .in3(N__2764),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_16_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_16_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_16_2  (
            .in0(N__2570),
            .in1(N__2604),
            .in2(N__2607),
            .in3(N__2942),
            .lcout(U409_ADDRESS_DECODE_Z2_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_8_LC_1_16_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_8_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_8_LC_1_16_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_8_LC_1_16_3  (
            .in0(N__2943),
            .in1(N__2598),
            .in2(N__2876),
            .in3(N__2571),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_16_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_16_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_16_5  (
            .in0(N__3164),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2597),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_2_LC_1_17_2 .C_ON=1'b0;
    defparam \U409_CIA.g0_2_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_2_LC_1_17_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_CIA.g0_2_LC_1_17_2  (
            .in0(N__2596),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2564),
            .lcout(),
            .ltout(\U409_CIA.g0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_13_LC_1_17_3 .C_ON=1'b0;
    defparam \U409_CIA.g0_13_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_13_LC_1_17_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_CIA.g0_13_LC_1_17_3  (
            .in0(N__3270),
            .in1(N__2936),
            .in2(N__2913),
            .in3(N__2823),
            .lcout(\U409_CIA.g0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_10_LC_1_17_6 .C_ON=1'b0;
    defparam \U409_CIA.g0_10_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_10_LC_1_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.g0_10_LC_1_17_6  (
            .in0(N__2905),
            .in1(N__2880),
            .in2(N__2851),
            .in3(N__3163),
            .lcout(\U409_CIA.g0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_8_LC_2_11_0 .C_ON=1'b0;
    defparam \U409_CIA.g0_8_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_8_LC_2_11_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_CIA.g0_8_LC_2_11_0  (
            .in0(N__3060),
            .in1(N__2793),
            .in2(_gnd_net_),
            .in3(N__5967),
            .lcout(),
            .ltout(\U409_CIA.g0Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_14_LC_2_11_1 .C_ON=1'b0;
    defparam \U409_CIA.g0_14_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_14_LC_2_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.g0_14_LC_2_11_1  (
            .in0(N__2712),
            .in1(N__2813),
            .in2(N__2817),
            .in3(N__2702),
            .lcout(\U409_CIA.g0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_2_11_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_2_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_2_11_4  (
            .in0(N__2701),
            .in1(N__2738),
            .in2(N__2814),
            .in3(N__2792),
            .lcout(CIA_SPACEm_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_11_LC_2_12_5 .C_ON=1'b0;
    defparam \U409_CIA.g0_11_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_11_LC_2_12_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_CIA.g0_11_LC_2_12_5  (
            .in0(N__2659),
            .in1(N__2772),
            .in2(N__2742),
            .in3(N__2637),
            .lcout(\U409_CIA.g0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un5_RAMSPACEn_LC_2_13_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un5_RAMSPACEn_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un5_RAMSPACEn_LC_2_13_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_ADDRESS_DECODE.un5_RAMSPACEn_LC_2_13_0  (
            .in0(N__3269),
            .in1(N__2636),
            .in2(_gnd_net_),
            .in3(N__3053),
            .lcout(U409_ADDRESS_DECODE_un5_RAMSPACEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.HIROM_LC_2_13_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.HIROM_LC_2_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.HIROM_LC_2_13_2  (
            .in0(N__3289),
            .in1(N__3052),
            .in2(N__3272),
            .in3(N__2706),
            .lcout(U409_ADDRESS_DECODE_HIROM),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_3_LC_2_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_3_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_3_LC_2_13_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_3_LC_2_13_4  (
            .in0(N__2669),
            .in1(N__3220),
            .in2(N__3273),
            .in3(N__2635),
            .lcout(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_2_15_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_2_15_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_2_15_1  (
            .in0(N__3224),
            .in1(N__3262),
            .in2(N__3378),
            .in3(N__3299),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_10_LC_2_16_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_10_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_10_LC_2_16_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_10_LC_2_16_4  (
            .in0(N__3054),
            .in1(N__5997),
            .in2(N__3271),
            .in3(N__3225),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_14_LC_2_16_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_14_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_14_LC_2_16_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_14_LC_2_16_5  (
            .in0(N__3198),
            .in1(N__3192),
            .in2(N__3186),
            .in3(N__3117),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_11_LC_3_17_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_11_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_11_LC_3_17_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_11_LC_3_17_2  (
            .in0(N__3183),
            .in1(N__5432),
            .in2(N__3168),
            .in3(N__3129),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_13_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_13_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_13_6  (
            .in0(N__3405),
            .in1(N__3059),
            .in2(_gnd_net_),
            .in3(N__3107),
            .lcout(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_14_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_14_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_14_5  (
            .in0(N__3028),
            .in1(N__3388),
            .in2(_gnd_net_),
            .in3(N__3111),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_6_15_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_6_15_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_6_15_6  (
            .in0(N__3069),
            .in1(N__3058),
            .in2(N__2984),
            .in3(N__5968),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_9_13_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_9_13_0 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_9_13_0  (
            .in0(N__3421),
            .in1(N__3406),
            .in2(N__2985),
            .in3(N__3337),
            .lcout(BUFENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_13_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_13_1 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_13_1  (
            .in0(N__3407),
            .in1(_gnd_net_),
            .in2(N__3342),
            .in3(N__3422),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_1_LC_9_13_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_1_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_1_LC_9_13_2 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_1_LC_9_13_2  (
            .in0(N__3423),
            .in1(N__3408),
            .in2(N__3357),
            .in3(N__3341),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER15Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_13_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_13_5 .LUT_INIT=16'b0000000001110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_13_5  (
            .in0(N__5455),
            .in1(N__4662),
            .in2(N__5372),
            .in3(N__3543),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__4638));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_14_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_14_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_14_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_14_2  (
            .in0(N__3650),
            .in1(N__3512),
            .in2(_gnd_net_),
            .in3(N__4713),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__4627));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_8_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__4138),
            .in2(N__4085),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_8_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_10_8_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_10_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(N__4157),
            .in2(_gnd_net_),
            .in3(N__3312),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__4824),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_10_8_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_10_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_10_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(N__4037),
            .in2(_gnd_net_),
            .in3(N__3309),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__4824),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_10_8_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_10_8_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4101),
            .in3(N__3306),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_10_8_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_10_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_10_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_10_8_4  (
            .in0(_gnd_net_),
            .in1(N__4112),
            .in2(_gnd_net_),
            .in3(N__3303),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__4824),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_10_8_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_10_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(N__4355),
            .in2(_gnd_net_),
            .in3(N__3453),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_10_8_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_10_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_10_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_10_8_6  (
            .in0(_gnd_net_),
            .in1(N__4457),
            .in2(_gnd_net_),
            .in3(N__3450),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__4824),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_10_8_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_10_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_10_8_7  (
            .in0(_gnd_net_),
            .in1(N__4385),
            .in2(_gnd_net_),
            .in3(N__3447),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_10_9_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_10_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__4370),
            .in2(_gnd_net_),
            .in3(N__3444),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_10_9_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_10_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__4484),
            .in2(_gnd_net_),
            .in3(N__3441),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__4826),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_10_9_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_10_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_10_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__4052),
            .in2(_gnd_net_),
            .in3(N__3438),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__4826),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_10_9_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_10_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__4169),
            .in2(_gnd_net_),
            .in3(N__3435),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__4826),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_10_9_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_10_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_10_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__4472),
            .in2(_gnd_net_),
            .in3(N__3432),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__4826),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_10_9_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_10_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__4397),
            .in2(_gnd_net_),
            .in3(N__3429),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_10_9_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_10_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__4445),
            .in2(_gnd_net_),
            .in3(N__3426),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_10_9_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_10_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_10_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__4125),
            .in2(_gnd_net_),
            .in3(N__3486),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4826),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_10_10_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_10_10_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_10_10_1  (
            .in0(N__4025),
            .in1(N__4341),
            .in2(N__4434),
            .in3(N__3483),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4827),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_10_10_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_10_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_10_10_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_10_10_2  (
            .in0(N__4342),
            .in1(N__4026),
            .in2(N__3477),
            .in3(N__4433),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4827),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_10_10_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_10_10_4 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_10_10_4  (
            .in0(N__4340),
            .in1(N__4024),
            .in2(N__3468),
            .in3(N__4429),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4827),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_13_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_13_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_13_0 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_13_0  (
            .in0(N__3575),
            .in1(N__3542),
            .in2(_gnd_net_),
            .in3(N__4714),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__4626));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_13_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_13_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_13_1 .LUT_INIT=16'b0111100001111000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_13_1  (
            .in0(N__3541),
            .in1(N__3576),
            .in2(N__3597),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__4626));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_13_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_13_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__3574),
            .in2(_gnd_net_),
            .in3(N__3591),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_13_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_13_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_10_13_3  (
            .in0(N__3638),
            .in1(N__3611),
            .in2(N__3459),
            .in3(N__3492),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_2_LC_10_13_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_2_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_2_LC_10_13_4 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_2_LC_10_13_4  (
            .in0(N__5365),
            .in1(N__5459),
            .in2(N__3456),
            .in3(N__4649),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_13_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_13_5 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(N__3618),
            .in2(N__3660),
            .in3(N__3612),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__4626));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_13_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_13_6 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_13_6  (
            .in0(N__3639),
            .in1(N__3513),
            .in2(N__3654),
            .in3(N__4715),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__4626));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_14_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_14_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_14_1  (
            .in0(N__3572),
            .in1(N__3596),
            .in2(_gnd_net_),
            .in3(N__3539),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U842_4_LC_10_14_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U842_4_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U842_4_LC_10_14_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U842_4_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__4759),
            .in2(N__3657),
            .in3(N__4685),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIH6AR_6_LC_10_14_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIH6AR_6_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIH6AR_6_LC_10_14_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIH6AR_6_LC_10_14_3  (
            .in0(N__3637),
            .in1(N__3510),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_7_LC_10_14_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_7_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_7_LC_10_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_7_LC_10_14_4  (
            .in0(N__4747),
            .in1(N__4686),
            .in2(N__3621),
            .in3(N__4729),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_7_LC_10_14_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_7_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_7_LC_10_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_7_LC_10_14_5  (
            .in0(N__4681),
            .in1(N__3538),
            .in2(N__4761),
            .in3(N__3610),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_2_LC_10_14_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_2_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_2_LC_10_14_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_2_LC_10_14_6  (
            .in0(N__3595),
            .in1(N__3573),
            .in2(N__3552),
            .in3(N__3549),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_5_LC_10_14_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_5_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_5_LC_10_14_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_5_LC_10_14_7  (
            .in0(N__3540),
            .in1(N__3511),
            .in2(N__4689),
            .in3(N__4746),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_16_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_16_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_16_5  (
            .in0(N__5990),
            .in1(N__3789),
            .in2(_gnd_net_),
            .in3(N__3761),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_4_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_4_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_4_4  (
            .in0(N__4305),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3738),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS1n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_11_4_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_11_4_7 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_11_4_7  (
            .in0(N__3699),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4304),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS0n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_11_5_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_11_5_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_11_5_0  (
            .in0(N__3877),
            .in1(_gnd_net_),
            .in2(N__3900),
            .in3(_gnd_net_),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4819),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_11_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_11_5_1 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_11_5_1  (
            .in0(N__4881),
            .in1(N__4914),
            .in2(N__3882),
            .in3(N__4953),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4819),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_11_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_11_5_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_11_5_2  (
            .in0(N__4913),
            .in1(N__4956),
            .in2(N__3801),
            .in3(N__4883),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4819),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_11_5_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_11_5_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_11_5_3  (
            .in0(N__3822),
            .in1(N__3840),
            .in2(_gnd_net_),
            .in3(N__3876),
            .lcout(\U409_TICK.TICK503_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_11_5_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_11_5_4 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_11_5_4  (
            .in0(N__3810),
            .in1(N__4955),
            .in2(N__4923),
            .in3(N__4884),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4819),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_5_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_5_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_5_5  (
            .in0(N__3996),
            .in1(N__3855),
            .in2(N__4209),
            .in3(N__3896),
            .lcout(),
            .ltout(\U409_TICK.TICK503_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_11_5_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_11_5_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_11_5_6  (
            .in0(N__3930),
            .in1(N__3957),
            .in2(N__3924),
            .in3(N__3978),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_11_5_7 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_11_5_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK50_LC_11_5_7  (
            .in0(N__4882),
            .in1(N__3911),
            .in2(N__3921),
            .in3(N__4954),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4819),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_11_6_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_11_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__3895),
            .in2(N__3881),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_11_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_11_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__3854),
            .in2(_gnd_net_),
            .in3(N__3843),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__4821),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_11_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_11_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__3839),
            .in2(_gnd_net_),
            .in3(N__3828),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__4821),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_11_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_11_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__5006),
            .in2(_gnd_net_),
            .in3(N__3825),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__4821),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_11_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_11_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(N__3821),
            .in2(_gnd_net_),
            .in3(N__3804),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_11_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_11_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__4574),
            .in2(_gnd_net_),
            .in3(N__3792),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_11_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_11_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(N__4526),
            .in2(_gnd_net_),
            .in3(N__3999),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__4821),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_11_6_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_11_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(N__3995),
            .in2(_gnd_net_),
            .in3(N__3984),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__4821),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_11_7_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_11_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__4838),
            .in2(_gnd_net_),
            .in3(N__3981),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_11_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_11_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__3974),
            .in2(_gnd_net_),
            .in3(N__3963),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__4822),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_11_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_11_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__4553),
            .in2(_gnd_net_),
            .in3(N__3960),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_11_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_11_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__3953),
            .in2(_gnd_net_),
            .in3(N__3942),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__4822),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_11_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_11_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__4985),
            .in2(_gnd_net_),
            .in3(N__3939),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_11_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_11_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__4967),
            .in2(_gnd_net_),
            .in3(N__3936),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_11_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_11_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__4541),
            .in2(_gnd_net_),
            .in3(N__3933),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_11_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_11_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__4205),
            .in2(_gnd_net_),
            .in3(N__4212),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4822),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_11_8_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_11_8_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_11_8_1  (
            .in0(N__4021),
            .in1(N__4426),
            .in2(N__4343),
            .in3(N__4191),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4823),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_11_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_11_8_2 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_11_8_2  (
            .in0(N__4425),
            .in1(N__4020),
            .in2(N__4086),
            .in3(N__4332),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4823),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_11_8_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_11_8_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_11_8_3  (
            .in0(N__4023),
            .in1(N__4428),
            .in2(N__4344),
            .in3(N__4185),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4823),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_11_8_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_11_8_4 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_11_8_4  (
            .in0(N__4427),
            .in1(N__4022),
            .in2(N__4179),
            .in3(N__4336),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4823),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_11_8_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_11_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4146),
            .in3(N__4081),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4823),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_11_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_11_8_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_11_8_7  (
            .in0(N__4170),
            .in1(N__4158),
            .in2(N__4145),
            .in3(N__4124),
            .lcout(\U409_TICK.TICK603_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_11_9_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_11_9_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_11_9_2  (
            .in0(N__4113),
            .in1(N__4100),
            .in2(_gnd_net_),
            .in3(N__4080),
            .lcout(),
            .ltout(\U409_TICK.TICK603_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_11_9_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_11_9_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_11_9_3  (
            .in0(N__4059),
            .in1(N__4053),
            .in2(N__4041),
            .in3(N__4038),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_11_9_4 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_11_9_4 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \U409_TICK.TICK60_LC_11_9_4  (
            .in0(N__4496),
            .in1(N__4424),
            .in2(N__4515),
            .in3(N__4331),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4825),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_11_9_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_11_9_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_11_9_6  (
            .in0(N__4485),
            .in1(N__4473),
            .in2(N__4461),
            .in3(N__4446),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_11_9_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_11_9_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_11_9_7  (
            .in0(N__4398),
            .in1(N__4386),
            .in2(N__4374),
            .in3(N__4359),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_11_10_2 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_11_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5303),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5183),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_HOLD_LC_11_10_3 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_HOLD_LC_11_10_3 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U409_CIA.CIA_HOLD_LC_11_10_3  (
            .in0(N__4274),
            .in1(N__5202),
            .in2(N__4247),
            .in3(N__4288),
            .lcout(\U409_CIA.CIA_HOLDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5183),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_11_10_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_11_10_7 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_11_10_7  (
            .in0(N__4275),
            .in1(N__5203),
            .in2(N__4248),
            .in3(N__4289),
            .lcout(CIA_ENABLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_11_2 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_11_2  (
            .in0(N__4290),
            .in1(N__4268),
            .in2(N__4246),
            .in3(N__5205),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__5639));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_12_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5529),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .ce(),
            .sr(N__5640));
    defparam \U409_TRANSFER_ACK.ROMENn_LC_11_13_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_11_13_3 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_11_13_3 .LUT_INIT=16'b1100101011101110;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_LC_11_13_3  (
            .in0(N__4772),
            .in1(N__5475),
            .in2(N__5789),
            .in3(N__5481),
            .lcout(ROMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .ce(),
            .sr(N__5641));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_14_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_14_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_14_1 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_14_1  (
            .in0(N__4687),
            .in1(N__4731),
            .in2(N__4716),
            .in3(N__4760),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .ce(),
            .sr(N__4634));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_14_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_14_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_14_4 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_14_4  (
            .in0(N__4730),
            .in1(N__4688),
            .in2(_gnd_net_),
            .in3(N__4709),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .ce(),
            .sr(N__4634));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_14_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_14_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_14_7 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_14_7  (
            .in0(N__5573),
            .in1(N__4661),
            .in2(_gnd_net_),
            .in3(N__4650),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .ce(),
            .sr(N__4634));
    defparam CONSTANT_ONE_LUT4_LC_12_1_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_12_6_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_12_6_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_12_6_0  (
            .in0(N__4920),
            .in1(N__4951),
            .in2(N__4890),
            .in3(N__4581),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4820),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_12_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_12_6_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_12_6_1  (
            .in0(N__4554),
            .in1(N__4575),
            .in2(N__4842),
            .in3(N__4986),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_12_6_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_12_6_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_12_6_2  (
            .in0(N__4918),
            .in1(N__4949),
            .in2(N__4563),
            .in3(N__4560),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4820),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_12_6_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_12_6_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_12_6_3  (
            .in0(N__4968),
            .in1(N__4542),
            .in2(N__4530),
            .in3(N__5007),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_12_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_12_6_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_12_6_4  (
            .in0(N__4919),
            .in1(N__4880),
            .in2(N__4995),
            .in3(N__4992),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4820),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_12_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_12_6_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_12_6_5  (
            .in0(N__4950),
            .in1(N__4921),
            .in2(N__4888),
            .in3(N__4974),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4820),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_12_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_12_6_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_12_6_7  (
            .in0(N__4952),
            .in1(N__4922),
            .in2(N__4889),
            .in3(N__4848),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4820),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__5263),
            .in2(N__5304),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__5028),
            .in2(_gnd_net_),
            .in3(N__4794),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__5184),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__5238),
            .in2(_gnd_net_),
            .in3(N__4791),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__5074),
            .in2(_gnd_net_),
            .in3(N__4788),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__5184),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__5050),
            .in2(_gnd_net_),
            .in3(N__4785),
            .lcout(),
            .ltout(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_12_9_5  (
            .in0(N__5240),
            .in1(N__5090),
            .in2(N__5103),
            .in3(N__5297),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5184),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_6 .LUT_INIT=16'b0011001101001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_12_9_6  (
            .in0(N__5298),
            .in1(N__5100),
            .in2(N__5094),
            .in3(N__5239),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5184),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_12_9_7  (
            .in0(N__5264),
            .in1(N__5075),
            .in2(N__5055),
            .in3(N__5029),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_12_10_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_12_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__5302),
            .in2(_gnd_net_),
            .in3(N__5267),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5182),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_12_10_1 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_12_10_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_12_10_1  (
            .in0(N__5046),
            .in1(N__5073),
            .in2(_gnd_net_),
            .in3(N__5030),
            .lcout(\U409_CIA.CLKCIA8_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_2_LC_12_10_2 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_12_10_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_CIA.CLKCIA_RNO_2_LC_12_10_2  (
            .in0(N__5241),
            .in1(N__5299),
            .in2(_gnd_net_),
            .in3(N__5265),
            .lcout(),
            .ltout(\U409_CIA.N_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_0_LC_12_10_3 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_12_10_3 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \U409_CIA.CLKCIA_RNO_0_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__5158),
            .in2(N__5082),
            .in3(N__5213),
            .lcout(),
            .ltout(\U409_CIA.CLKCIAZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_LC_12_10_4 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLKCIA_LC_12_10_4 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \U409_CIA.CLKCIA_LC_12_10_4  (
            .in0(N__5013),
            .in1(N__5301),
            .in2(N__5079),
            .in3(N__5268),
            .lcout(CLKCIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5182),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_1_LC_12_10_5 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_12_10_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CLKCIA_RNO_1_LC_12_10_5  (
            .in0(N__5076),
            .in1(N__5243),
            .in2(N__5054),
            .in3(N__5031),
            .lcout(\U409_CIA.CLKCIA6_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_12_10_6 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_12_10_6 .LUT_INIT=16'b0100010000100010;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_12_10_6  (
            .in0(N__5242),
            .in1(N__5300),
            .in2(_gnd_net_),
            .in3(N__5266),
            .lcout(),
            .ltout(\U409_CIA.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_12_10_7 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_12_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_12_10_7 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \U409_CIA.VMA_LC_12_10_7  (
            .in0(N__5204),
            .in1(N__5244),
            .in2(N__5217),
            .in3(N__5214),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5182),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_12_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_12_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5159),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__5642));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_12_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_12_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5136),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__5642));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_12_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_12_12_0 .LUT_INIT=16'b0000010100110011;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_12_12_0  (
            .in0(N__5528),
            .in1(N__5109),
            .in2(N__5508),
            .in3(N__5739),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_12_1 .LUT_INIT=16'b0000110010001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_12_1  (
            .in0(N__5740),
            .in1(N__5971),
            .in2(N__5142),
            .in3(N__5772),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_12_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_12_12_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_12_12_2  (
            .in0(N__5135),
            .in1(N__5338),
            .in2(N__5121),
            .in3(N__5738),
            .lcout(\U409_TRANSFER_ACK.N_132 ),
            .ltout(\U409_TRANSFER_ACK.N_132_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_12_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_12_12_3 .LUT_INIT=16'b0000010100100111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_12_12_3  (
            .in0(N__5770),
            .in1(N__5503),
            .in2(N__5139),
            .in3(N__5526),
            .lcout(\U409_TRANSFER_ACK.m9_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_12_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_12_12_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__5134),
            .in2(_gnd_net_),
            .in3(N__5117),
            .lcout(\U409_TRANSFER_ACK.N_4 ),
            .ltout(\U409_TRANSFER_ACK.N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_12_12_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_12_12_6 .LUT_INIT=16'b1101000111110011;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_12_12_6  (
            .in0(N__5527),
            .in1(N__5769),
            .in2(N__5511),
            .in3(N__5507),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.m9_am_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_12_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_12_7 .LUT_INIT=16'b0000010010001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_12_7  (
            .in0(N__5741),
            .in1(N__5970),
            .in2(N__5490),
            .in3(N__5487),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_13_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_13_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_13_2  (
            .in0(N__5663),
            .in1(N__5689),
            .in2(_gnd_net_),
            .in3(N__5716),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_13_5 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_13_5  (
            .in0(N__5717),
            .in1(_gnd_net_),
            .in2(N__5697),
            .in3(N__5664),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_12_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_12_13_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_12_13_6  (
            .in0(N__5469),
            .in1(N__5460),
            .in2(N__5355),
            .in3(N__5972),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_13_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_13_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_13_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_13_7  (
            .in0(N__5409),
            .in1(N__5387),
            .in2(_gnd_net_),
            .in3(N__5342),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_14_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_14_1 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_14_1  (
            .in0(N__5408),
            .in1(N__5388),
            .in2(N__5354),
            .in3(N__5586),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net ),
            .ce(),
            .sr(N__5646));
    defparam RESETn_ibuf_RNIM9SF_LC_13_12_3.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_13_12_3.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_13_12_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_13_12_3 (
            .in0(N__5969),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_13_13_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_13_13_0 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_13_13_0  (
            .in0(N__5696),
            .in1(N__5665),
            .in2(N__5790),
            .in3(N__5718),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5618));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_13_13_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_13_13_3 .LUT_INIT=16'b0101010000001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_13_13_3  (
            .in0(N__5771),
            .in1(N__5544),
            .in2(N__5751),
            .in3(N__5742),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5618));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_13_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_13_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_13_5  (
            .in0(N__5719),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5693),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5618));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_13_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_13_13_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_13_13_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_13_13_6  (
            .in0(N__5694),
            .in1(N__5666),
            .in2(_gnd_net_),
            .in3(N__5720),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5618));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_13_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_13_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_13_7 .LUT_INIT=16'b1011111100100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_13_7  (
            .in0(N__5721),
            .in1(N__5695),
            .in2(N__5670),
            .in3(N__5558),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5618));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_13_14_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_13_14_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_13_14_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_13_14_1  (
            .in0(N__5862),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5974),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_13_14_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_13_14_2 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_13_14_2  (
            .in0(N__5975),
            .in1(N__6022),
            .in2(_gnd_net_),
            .in3(N__5861),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_13_14_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_13_14_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_13_14_4  (
            .in0(N__5585),
            .in1(N__5574),
            .in2(N__5559),
            .in3(N__5543),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER6 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_13_14_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_13_14_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_13_14_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_13_14_5  (
            .in0(N__5863),
            .in1(N__5973),
            .in2(N__5532),
            .in3(N__6023),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_14_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_14_13_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_14_13_5  (
            .in0(N__6020),
            .in1(N__5864),
            .in2(_gnd_net_),
            .in3(N__5840),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_14_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_14_13_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_14_13_6 .LUT_INIT=16'b0100111001001100;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_14_13_6  (
            .in0(N__5976),
            .in1(N__6035),
            .in2(N__6048),
            .in3(N__6021),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_14_14_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_14_14_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_14_14_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_LC_14_14_2  (
            .in0(N__6024),
            .in1(N__5977),
            .in2(N__5868),
            .in3(N__5841),
            .lcout(TACK_EN_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .ce(N__5829),
            .sr(_gnd_net_));
    defparam TACKn_iobuf_RNO_LC_18_15_6.C_ON=1'b0;
    defparam TACKn_iobuf_RNO_LC_18_15_6.SEQ_MODE=4'b0000;
    defparam TACKn_iobuf_RNO_LC_18_15_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_iobuf_RNO_LC_18_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5823),
            .lcout(N_359_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 13 2025 09:32:57

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U111_TOP" view "INTERFACE"

module U111_TOP (
    D_LM_AMIGA,
    D_UM_AMIGA,
    D_LL_AMIGA,
    D_UU_AMIGA,
    D_LL_040,
    D_UU_040,
    D_LM_040,
    D_UM_040,
    A_AMIGA,
    A_040,
    SIZ,
    TBIn,
    TEAn,
    TSn,
    RESETn,
    CLKRAMA,
    PORTSIZE,
    DMAAn,
    TEA_CPUn,
    LBENn,
    CLK40B,
    TBI_CPUn,
    TAn,
    CPUBGn,
    BUFENn,
    RnW,
    CLK80_CPU,
    BUFDIR,
    TCI_CPUn,
    TS_CPUn,
    CLKRAMB,
    CLK40A,
    TCIn,
    CLK40C,
    CLK40_IN,
    BBn,
    TACKn,
    BGn);

    inout [7:0] D_LM_AMIGA;
    inout [7:0] D_UM_AMIGA;
    inout [7:0] D_LL_AMIGA;
    inout [7:0] D_UU_AMIGA;
    inout [7:0] D_LL_040;
    inout [7:0] D_UU_040;
    inout [7:0] D_LM_040;
    inout [7:0] D_UM_040;
    output [1:0] A_AMIGA;
    input [1:0] A_040;
    input [1:0] SIZ;
    input TBIn;
    input TEAn;
    inout TSn;
    input RESETn;
    output CLKRAMA;
    input PORTSIZE;
    output DMAAn;
    output TEA_CPUn;
    input LBENn;
    output CLK40B;
    output TBI_CPUn;
    inout TAn;
    output CPUBGn;
    output BUFENn;
    input RnW;
    output CLK80_CPU;
    output BUFDIR;
    output TCI_CPUn;
    inout TS_CPUn;
    output CLKRAMB;
    output CLK40A;
    input TCIn;
    output CLK40C;
    input CLK40_IN;
    input BBn;
    inout TACKn;
    input BGn;

    wire N__9464;
    wire N__9448;
    wire N__9447;
    wire N__9446;
    wire N__9439;
    wire N__9438;
    wire N__9437;
    wire N__9430;
    wire N__9429;
    wire N__9428;
    wire N__9421;
    wire N__9420;
    wire N__9419;
    wire N__9412;
    wire N__9411;
    wire N__9410;
    wire N__9403;
    wire N__9402;
    wire N__9401;
    wire N__9394;
    wire N__9393;
    wire N__9392;
    wire N__9385;
    wire N__9384;
    wire N__9383;
    wire N__9376;
    wire N__9375;
    wire N__9374;
    wire N__9367;
    wire N__9366;
    wire N__9365;
    wire N__9358;
    wire N__9357;
    wire N__9356;
    wire N__9349;
    wire N__9348;
    wire N__9347;
    wire N__9340;
    wire N__9339;
    wire N__9338;
    wire N__9331;
    wire N__9330;
    wire N__9329;
    wire N__9322;
    wire N__9321;
    wire N__9320;
    wire N__9313;
    wire N__9312;
    wire N__9311;
    wire N__9304;
    wire N__9303;
    wire N__9302;
    wire N__9295;
    wire N__9294;
    wire N__9293;
    wire N__9286;
    wire N__9285;
    wire N__9284;
    wire N__9277;
    wire N__9276;
    wire N__9275;
    wire N__9268;
    wire N__9267;
    wire N__9266;
    wire N__9259;
    wire N__9258;
    wire N__9257;
    wire N__9250;
    wire N__9249;
    wire N__9248;
    wire N__9241;
    wire N__9240;
    wire N__9239;
    wire N__9232;
    wire N__9231;
    wire N__9230;
    wire N__9223;
    wire N__9222;
    wire N__9221;
    wire N__9214;
    wire N__9213;
    wire N__9212;
    wire N__9205;
    wire N__9204;
    wire N__9203;
    wire N__9196;
    wire N__9195;
    wire N__9194;
    wire N__9187;
    wire N__9186;
    wire N__9185;
    wire N__9178;
    wire N__9177;
    wire N__9176;
    wire N__9169;
    wire N__9168;
    wire N__9167;
    wire N__9160;
    wire N__9159;
    wire N__9158;
    wire N__9151;
    wire N__9150;
    wire N__9149;
    wire N__9142;
    wire N__9141;
    wire N__9140;
    wire N__9133;
    wire N__9132;
    wire N__9131;
    wire N__9124;
    wire N__9123;
    wire N__9122;
    wire N__9115;
    wire N__9114;
    wire N__9113;
    wire N__9106;
    wire N__9105;
    wire N__9104;
    wire N__9097;
    wire N__9096;
    wire N__9095;
    wire N__9088;
    wire N__9087;
    wire N__9086;
    wire N__9079;
    wire N__9078;
    wire N__9077;
    wire N__9070;
    wire N__9069;
    wire N__9068;
    wire N__9061;
    wire N__9060;
    wire N__9059;
    wire N__9052;
    wire N__9051;
    wire N__9050;
    wire N__9043;
    wire N__9042;
    wire N__9041;
    wire N__9034;
    wire N__9033;
    wire N__9032;
    wire N__9025;
    wire N__9024;
    wire N__9023;
    wire N__9016;
    wire N__9015;
    wire N__9014;
    wire N__9007;
    wire N__9006;
    wire N__9005;
    wire N__8998;
    wire N__8997;
    wire N__8996;
    wire N__8989;
    wire N__8988;
    wire N__8987;
    wire N__8980;
    wire N__8979;
    wire N__8978;
    wire N__8971;
    wire N__8970;
    wire N__8969;
    wire N__8962;
    wire N__8961;
    wire N__8960;
    wire N__8953;
    wire N__8952;
    wire N__8951;
    wire N__8944;
    wire N__8943;
    wire N__8942;
    wire N__8935;
    wire N__8934;
    wire N__8933;
    wire N__8926;
    wire N__8925;
    wire N__8924;
    wire N__8917;
    wire N__8916;
    wire N__8915;
    wire N__8908;
    wire N__8907;
    wire N__8906;
    wire N__8899;
    wire N__8898;
    wire N__8897;
    wire N__8890;
    wire N__8889;
    wire N__8888;
    wire N__8881;
    wire N__8880;
    wire N__8879;
    wire N__8872;
    wire N__8871;
    wire N__8870;
    wire N__8863;
    wire N__8862;
    wire N__8861;
    wire N__8854;
    wire N__8853;
    wire N__8852;
    wire N__8845;
    wire N__8844;
    wire N__8843;
    wire N__8836;
    wire N__8835;
    wire N__8834;
    wire N__8827;
    wire N__8826;
    wire N__8825;
    wire N__8818;
    wire N__8817;
    wire N__8816;
    wire N__8809;
    wire N__8808;
    wire N__8807;
    wire N__8800;
    wire N__8799;
    wire N__8798;
    wire N__8791;
    wire N__8790;
    wire N__8789;
    wire N__8782;
    wire N__8781;
    wire N__8780;
    wire N__8773;
    wire N__8772;
    wire N__8771;
    wire N__8764;
    wire N__8763;
    wire N__8762;
    wire N__8755;
    wire N__8754;
    wire N__8753;
    wire N__8746;
    wire N__8745;
    wire N__8744;
    wire N__8737;
    wire N__8736;
    wire N__8735;
    wire N__8728;
    wire N__8727;
    wire N__8726;
    wire N__8719;
    wire N__8718;
    wire N__8717;
    wire N__8710;
    wire N__8709;
    wire N__8708;
    wire N__8701;
    wire N__8700;
    wire N__8699;
    wire N__8692;
    wire N__8691;
    wire N__8690;
    wire N__8683;
    wire N__8682;
    wire N__8681;
    wire N__8674;
    wire N__8673;
    wire N__8672;
    wire N__8665;
    wire N__8664;
    wire N__8663;
    wire N__8656;
    wire N__8655;
    wire N__8654;
    wire N__8647;
    wire N__8646;
    wire N__8645;
    wire N__8638;
    wire N__8637;
    wire N__8636;
    wire N__8629;
    wire N__8628;
    wire N__8627;
    wire N__8620;
    wire N__8619;
    wire N__8618;
    wire N__8611;
    wire N__8610;
    wire N__8609;
    wire N__8602;
    wire N__8601;
    wire N__8600;
    wire N__8593;
    wire N__8592;
    wire N__8591;
    wire N__8574;
    wire N__8571;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8544;
    wire N__8541;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8523;
    wire N__8520;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8466;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8452;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8436;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8426;
    wire N__8425;
    wire N__8424;
    wire N__8423;
    wire N__8422;
    wire N__8421;
    wire N__8416;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8404;
    wire N__8403;
    wire N__8402;
    wire N__8401;
    wire N__8398;
    wire N__8397;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8385;
    wire N__8382;
    wire N__8375;
    wire N__8372;
    wire N__8369;
    wire N__8366;
    wire N__8365;
    wire N__8364;
    wire N__8363;
    wire N__8360;
    wire N__8351;
    wire N__8346;
    wire N__8343;
    wire N__8338;
    wire N__8337;
    wire N__8334;
    wire N__8331;
    wire N__8328;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8304;
    wire N__8301;
    wire N__8298;
    wire N__8295;
    wire N__8292;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8238;
    wire N__8235;
    wire N__8232;
    wire N__8229;
    wire N__8226;
    wire N__8223;
    wire N__8220;
    wire N__8217;
    wire N__8214;
    wire N__8211;
    wire N__8208;
    wire N__8205;
    wire N__8202;
    wire N__8199;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8171;
    wire N__8168;
    wire N__8165;
    wire N__8160;
    wire N__8157;
    wire N__8154;
    wire N__8151;
    wire N__8148;
    wire N__8145;
    wire N__8142;
    wire N__8139;
    wire N__8136;
    wire N__8133;
    wire N__8132;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8097;
    wire N__8094;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8082;
    wire N__8079;
    wire N__8076;
    wire N__8073;
    wire N__8070;
    wire N__8067;
    wire N__8064;
    wire N__8061;
    wire N__8058;
    wire N__8055;
    wire N__8052;
    wire N__8049;
    wire N__8048;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8013;
    wire N__8010;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7977;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7922;
    wire N__7921;
    wire N__7920;
    wire N__7919;
    wire N__7918;
    wire N__7917;
    wire N__7910;
    wire N__7909;
    wire N__7904;
    wire N__7903;
    wire N__7902;
    wire N__7901;
    wire N__7898;
    wire N__7897;
    wire N__7896;
    wire N__7895;
    wire N__7894;
    wire N__7893;
    wire N__7890;
    wire N__7887;
    wire N__7884;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7872;
    wire N__7871;
    wire N__7868;
    wire N__7861;
    wire N__7856;
    wire N__7853;
    wire N__7852;
    wire N__7851;
    wire N__7850;
    wire N__7847;
    wire N__7844;
    wire N__7841;
    wire N__7840;
    wire N__7839;
    wire N__7834;
    wire N__7831;
    wire N__7828;
    wire N__7825;
    wire N__7822;
    wire N__7819;
    wire N__7818;
    wire N__7817;
    wire N__7814;
    wire N__7809;
    wire N__7808;
    wire N__7807;
    wire N__7806;
    wire N__7805;
    wire N__7802;
    wire N__7795;
    wire N__7790;
    wire N__7787;
    wire N__7782;
    wire N__7777;
    wire N__7774;
    wire N__7769;
    wire N__7764;
    wire N__7757;
    wire N__7754;
    wire N__7753;
    wire N__7752;
    wire N__7751;
    wire N__7750;
    wire N__7747;
    wire N__7742;
    wire N__7737;
    wire N__7730;
    wire N__7723;
    wire N__7716;
    wire N__7713;
    wire N__7698;
    wire N__7695;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7659;
    wire N__7656;
    wire N__7653;
    wire N__7650;
    wire N__7647;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7635;
    wire N__7632;
    wire N__7629;
    wire N__7626;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7602;
    wire N__7601;
    wire N__7598;
    wire N__7595;
    wire N__7590;
    wire N__7587;
    wire N__7586;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7570;
    wire N__7567;
    wire N__7564;
    wire N__7561;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7542;
    wire N__7539;
    wire N__7536;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7494;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7476;
    wire N__7473;
    wire N__7470;
    wire N__7467;
    wire N__7464;
    wire N__7461;
    wire N__7458;
    wire N__7455;
    wire N__7452;
    wire N__7449;
    wire N__7446;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7438;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7424;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7409;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7399;
    wire N__7396;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7384;
    wire N__7381;
    wire N__7374;
    wire N__7371;
    wire N__7368;
    wire N__7365;
    wire N__7362;
    wire N__7359;
    wire N__7356;
    wire N__7353;
    wire N__7350;
    wire N__7347;
    wire N__7344;
    wire N__7341;
    wire N__7338;
    wire N__7335;
    wire N__7332;
    wire N__7329;
    wire N__7326;
    wire N__7323;
    wire N__7320;
    wire N__7319;
    wire N__7318;
    wire N__7315;
    wire N__7312;
    wire N__7309;
    wire N__7302;
    wire N__7301;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7278;
    wire N__7275;
    wire N__7272;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7259;
    wire N__7258;
    wire N__7257;
    wire N__7256;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7242;
    wire N__7239;
    wire N__7236;
    wire N__7231;
    wire N__7230;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7210;
    wire N__7207;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7191;
    wire N__7190;
    wire N__7189;
    wire N__7188;
    wire N__7185;
    wire N__7178;
    wire N__7177;
    wire N__7176;
    wire N__7175;
    wire N__7174;
    wire N__7173;
    wire N__7172;
    wire N__7171;
    wire N__7170;
    wire N__7169;
    wire N__7168;
    wire N__7167;
    wire N__7164;
    wire N__7161;
    wire N__7148;
    wire N__7141;
    wire N__7140;
    wire N__7139;
    wire N__7138;
    wire N__7137;
    wire N__7134;
    wire N__7131;
    wire N__7128;
    wire N__7125;
    wire N__7122;
    wire N__7119;
    wire N__7112;
    wire N__7109;
    wire N__7092;
    wire N__7089;
    wire N__7088;
    wire N__7087;
    wire N__7084;
    wire N__7081;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7068;
    wire N__7067;
    wire N__7064;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7047;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7035;
    wire N__7032;
    wire N__7029;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7011;
    wire N__7010;
    wire N__7009;
    wire N__7006;
    wire N__7005;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6997;
    wire N__6996;
    wire N__6995;
    wire N__6994;
    wire N__6991;
    wire N__6988;
    wire N__6985;
    wire N__6980;
    wire N__6977;
    wire N__6974;
    wire N__6973;
    wire N__6972;
    wire N__6971;
    wire N__6970;
    wire N__6969;
    wire N__6966;
    wire N__6963;
    wire N__6962;
    wire N__6961;
    wire N__6960;
    wire N__6953;
    wire N__6946;
    wire N__6943;
    wire N__6940;
    wire N__6937;
    wire N__6936;
    wire N__6933;
    wire N__6932;
    wire N__6931;
    wire N__6928;
    wire N__6927;
    wire N__6926;
    wire N__6925;
    wire N__6924;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6909;
    wire N__6908;
    wire N__6897;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6885;
    wire N__6882;
    wire N__6879;
    wire N__6876;
    wire N__6873;
    wire N__6870;
    wire N__6861;
    wire N__6860;
    wire N__6859;
    wire N__6856;
    wire N__6853;
    wire N__6852;
    wire N__6851;
    wire N__6850;
    wire N__6849;
    wire N__6844;
    wire N__6837;
    wire N__6826;
    wire N__6823;
    wire N__6820;
    wire N__6817;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6800;
    wire N__6797;
    wire N__6792;
    wire N__6789;
    wire N__6784;
    wire N__6781;
    wire N__6778;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6759;
    wire N__6756;
    wire N__6753;
    wire N__6750;
    wire N__6745;
    wire N__6742;
    wire N__6739;
    wire N__6734;
    wire N__6727;
    wire N__6720;
    wire N__6717;
    wire N__6714;
    wire N__6713;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6694;
    wire N__6689;
    wire N__6686;
    wire N__6681;
    wire N__6678;
    wire N__6675;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6663;
    wire N__6660;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6648;
    wire N__6645;
    wire N__6642;
    wire N__6641;
    wire N__6636;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6628;
    wire N__6627;
    wire N__6626;
    wire N__6621;
    wire N__6618;
    wire N__6613;
    wire N__6606;
    wire N__6605;
    wire N__6604;
    wire N__6603;
    wire N__6602;
    wire N__6601;
    wire N__6600;
    wire N__6597;
    wire N__6596;
    wire N__6595;
    wire N__6594;
    wire N__6593;
    wire N__6592;
    wire N__6591;
    wire N__6590;
    wire N__6589;
    wire N__6588;
    wire N__6585;
    wire N__6580;
    wire N__6577;
    wire N__6572;
    wire N__6569;
    wire N__6556;
    wire N__6549;
    wire N__6534;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6498;
    wire N__6497;
    wire N__6494;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6480;
    wire N__6477;
    wire N__6474;
    wire N__6471;
    wire N__6468;
    wire N__6465;
    wire N__6464;
    wire N__6463;
    wire N__6462;
    wire N__6459;
    wire N__6458;
    wire N__6457;
    wire N__6454;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6441;
    wire N__6438;
    wire N__6433;
    wire N__6430;
    wire N__6417;
    wire N__6414;
    wire N__6413;
    wire N__6410;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6390;
    wire N__6387;
    wire N__6386;
    wire N__6385;
    wire N__6384;
    wire N__6383;
    wire N__6382;
    wire N__6381;
    wire N__6380;
    wire N__6379;
    wire N__6378;
    wire N__6377;
    wire N__6376;
    wire N__6375;
    wire N__6374;
    wire N__6371;
    wire N__6342;
    wire N__6339;
    wire N__6338;
    wire N__6337;
    wire N__6336;
    wire N__6335;
    wire N__6334;
    wire N__6333;
    wire N__6332;
    wire N__6331;
    wire N__6312;
    wire N__6309;
    wire N__6306;
    wire N__6303;
    wire N__6300;
    wire N__6299;
    wire N__6296;
    wire N__6293;
    wire N__6292;
    wire N__6289;
    wire N__6286;
    wire N__6283;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6264;
    wire N__6261;
    wire N__6258;
    wire N__6255;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6243;
    wire N__6240;
    wire N__6237;
    wire N__6234;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6216;
    wire N__6215;
    wire N__6212;
    wire N__6209;
    wire N__6204;
    wire N__6201;
    wire N__6200;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6183;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6171;
    wire N__6168;
    wire N__6165;
    wire N__6162;
    wire N__6159;
    wire N__6156;
    wire N__6153;
    wire N__6150;
    wire N__6147;
    wire N__6144;
    wire N__6141;
    wire N__6138;
    wire N__6137;
    wire N__6134;
    wire N__6131;
    wire N__6130;
    wire N__6127;
    wire N__6124;
    wire N__6121;
    wire N__6118;
    wire N__6115;
    wire N__6112;
    wire N__6105;
    wire N__6102;
    wire N__6099;
    wire N__6096;
    wire N__6093;
    wire N__6090;
    wire N__6087;
    wire N__6084;
    wire N__6081;
    wire N__6080;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6053;
    wire N__6050;
    wire N__6047;
    wire N__6044;
    wire N__6041;
    wire N__6036;
    wire N__6033;
    wire N__6030;
    wire N__6027;
    wire N__6026;
    wire N__6023;
    wire N__6020;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5999;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5964;
    wire N__5961;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5943;
    wire N__5940;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5922;
    wire N__5919;
    wire N__5916;
    wire N__5913;
    wire N__5910;
    wire N__5907;
    wire N__5904;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5886;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5874;
    wire N__5871;
    wire N__5868;
    wire N__5865;
    wire N__5862;
    wire N__5859;
    wire N__5856;
    wire N__5853;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5829;
    wire N__5826;
    wire N__5823;
    wire N__5820;
    wire N__5817;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5802;
    wire N__5801;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5784;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5772;
    wire N__5769;
    wire N__5768;
    wire N__5765;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5754;
    wire N__5751;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5711;
    wire N__5708;
    wire N__5703;
    wire N__5700;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5688;
    wire N__5685;
    wire N__5682;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5668;
    wire N__5663;
    wire N__5660;
    wire N__5655;
    wire N__5652;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5634;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5622;
    wire N__5619;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5611;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5592;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5577;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5565;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5527;
    wire N__5522;
    wire N__5519;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5490;
    wire N__5487;
    wire N__5484;
    wire N__5481;
    wire N__5478;
    wire N__5475;
    wire N__5472;
    wire N__5469;
    wire N__5466;
    wire N__5463;
    wire N__5462;
    wire N__5459;
    wire N__5456;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5444;
    wire N__5441;
    wire N__5440;
    wire N__5437;
    wire N__5434;
    wire N__5431;
    wire N__5428;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5412;
    wire N__5409;
    wire N__5406;
    wire N__5403;
    wire N__5400;
    wire N__5397;
    wire N__5394;
    wire N__5391;
    wire N__5388;
    wire N__5385;
    wire N__5384;
    wire N__5383;
    wire N__5382;
    wire N__5381;
    wire N__5380;
    wire N__5377;
    wire N__5370;
    wire N__5367;
    wire N__5364;
    wire N__5361;
    wire N__5358;
    wire N__5355;
    wire N__5352;
    wire N__5351;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5339;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5323;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5307;
    wire N__5304;
    wire N__5301;
    wire N__5298;
    wire N__5295;
    wire N__5292;
    wire N__5289;
    wire N__5286;
    wire N__5283;
    wire N__5280;
    wire N__5277;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5205;
    wire N__5202;
    wire N__5199;
    wire N__5198;
    wire N__5195;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5154;
    wire N__5151;
    wire N__5148;
    wire N__5145;
    wire N__5142;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5130;
    wire N__5127;
    wire N__5124;
    wire N__5123;
    wire N__5122;
    wire N__5121;
    wire N__5116;
    wire N__5115;
    wire N__5114;
    wire N__5109;
    wire N__5106;
    wire N__5101;
    wire N__5094;
    wire N__5093;
    wire N__5090;
    wire N__5089;
    wire N__5088;
    wire N__5087;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5046;
    wire N__5045;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5035;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4977;
    wire N__4974;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4960;
    wire N__4957;
    wire N__4954;
    wire N__4951;
    wire N__4948;
    wire N__4943;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4931;
    wire N__4930;
    wire N__4929;
    wire N__4926;
    wire N__4923;
    wire N__4920;
    wire N__4919;
    wire N__4918;
    wire N__4917;
    wire N__4916;
    wire N__4915;
    wire N__4914;
    wire N__4911;
    wire N__4910;
    wire N__4909;
    wire N__4902;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4892;
    wire N__4891;
    wire N__4890;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4879;
    wire N__4878;
    wire N__4877;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4866;
    wire N__4865;
    wire N__4864;
    wire N__4863;
    wire N__4854;
    wire N__4851;
    wire N__4848;
    wire N__4845;
    wire N__4842;
    wire N__4841;
    wire N__4840;
    wire N__4839;
    wire N__4838;
    wire N__4835;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4775;
    wire N__4772;
    wire N__4761;
    wire N__4750;
    wire N__4739;
    wire N__4736;
    wire N__4735;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4708;
    wire N__4705;
    wire N__4700;
    wire N__4695;
    wire N__4692;
    wire N__4689;
    wire N__4686;
    wire N__4683;
    wire N__4680;
    wire N__4677;
    wire N__4670;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4650;
    wire N__4647;
    wire N__4646;
    wire N__4645;
    wire N__4644;
    wire N__4643;
    wire N__4642;
    wire N__4641;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4624;
    wire N__4619;
    wire N__4612;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4593;
    wire N__4590;
    wire N__4587;
    wire N__4586;
    wire N__4585;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4569;
    wire N__4568;
    wire N__4567;
    wire N__4566;
    wire N__4565;
    wire N__4560;
    wire N__4553;
    wire N__4548;
    wire N__4547;
    wire N__4544;
    wire N__4543;
    wire N__4542;
    wire N__4539;
    wire N__4538;
    wire N__4537;
    wire N__4534;
    wire N__4531;
    wire N__4524;
    wire N__4521;
    wire N__4520;
    wire N__4519;
    wire N__4516;
    wire N__4511;
    wire N__4506;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4494;
    wire N__4491;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4449;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4401;
    wire N__4400;
    wire N__4399;
    wire N__4396;
    wire N__4393;
    wire N__4390;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4362;
    wire N__4359;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4302;
    wire N__4299;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4265;
    wire N__4264;
    wire N__4257;
    wire N__4254;
    wire N__4251;
    wire N__4248;
    wire N__4245;
    wire N__4242;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4170;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4158;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4110;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4098;
    wire N__4095;
    wire N__4092;
    wire N__4089;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4074;
    wire N__4071;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4047;
    wire N__4046;
    wire N__4045;
    wire N__4044;
    wire N__4039;
    wire N__4034;
    wire N__4029;
    wire N__4028;
    wire N__4027;
    wire N__4024;
    wire N__4019;
    wire N__4016;
    wire N__4011;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3989;
    wire N__3988;
    wire N__3987;
    wire N__3984;
    wire N__3979;
    wire N__3976;
    wire N__3969;
    wire N__3966;
    wire N__3963;
    wire N__3960;
    wire N__3957;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3926;
    wire N__3923;
    wire N__3920;
    wire N__3915;
    wire N__3914;
    wire N__3913;
    wire N__3912;
    wire N__3911;
    wire N__3908;
    wire N__3903;
    wire N__3896;
    wire N__3891;
    wire N__3888;
    wire N__3885;
    wire N__3882;
    wire N__3879;
    wire N__3878;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3843;
    wire N__3840;
    wire N__3837;
    wire N__3834;
    wire N__3831;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3819;
    wire N__3816;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3804;
    wire N__3801;
    wire N__3798;
    wire N__3795;
    wire N__3792;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3759;
    wire N__3756;
    wire N__3753;
    wire N__3752;
    wire N__3751;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3711;
    wire N__3708;
    wire N__3707;
    wire N__3704;
    wire N__3701;
    wire N__3696;
    wire N__3693;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3681;
    wire N__3678;
    wire N__3675;
    wire N__3672;
    wire N__3669;
    wire N__3666;
    wire N__3663;
    wire N__3660;
    wire N__3657;
    wire N__3654;
    wire N__3651;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3629;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3615;
    wire N__3612;
    wire N__3609;
    wire N__3606;
    wire N__3603;
    wire N__3600;
    wire N__3597;
    wire N__3594;
    wire N__3591;
    wire N__3588;
    wire N__3585;
    wire N__3582;
    wire N__3579;
    wire N__3576;
    wire N__3573;
    wire N__3570;
    wire N__3567;
    wire N__3564;
    wire N__3561;
    wire N__3558;
    wire N__3555;
    wire N__3552;
    wire N__3549;
    wire N__3546;
    wire N__3543;
    wire N__3540;
    wire N__3537;
    wire N__3534;
    wire N__3531;
    wire N__3528;
    wire N__3525;
    wire N__3522;
    wire N__3519;
    wire N__3516;
    wire N__3513;
    wire N__3510;
    wire N__3507;
    wire N__3504;
    wire N__3501;
    wire N__3498;
    wire N__3495;
    wire N__3492;
    wire N__3489;
    wire N__3486;
    wire N__3483;
    wire N__3480;
    wire N__3477;
    wire N__3474;
    wire N__3471;
    wire N__3468;
    wire N__3465;
    wire N__3462;
    wire N__3461;
    wire N__3458;
    wire N__3455;
    wire N__3450;
    wire N__3447;
    wire N__3444;
    wire N__3441;
    wire N__3438;
    wire N__3435;
    wire N__3432;
    wire N__3429;
    wire N__3426;
    wire N__3423;
    wire N__3420;
    wire N__3417;
    wire N__3414;
    wire N__3411;
    wire N__3408;
    wire N__3405;
    wire N__3404;
    wire N__3399;
    wire N__3396;
    wire N__3393;
    wire N__3390;
    wire N__3389;
    wire N__3386;
    wire N__3383;
    wire N__3378;
    wire N__3375;
    wire N__3372;
    wire N__3369;
    wire N__3366;
    wire N__3363;
    wire N__3360;
    wire N__3357;
    wire N__3354;
    wire N__3351;
    wire N__3348;
    wire N__3345;
    wire N__3342;
    wire N__3341;
    wire N__3338;
    wire N__3335;
    wire N__3332;
    wire N__3329;
    wire N__3326;
    wire N__3323;
    wire N__3320;
    wire N__3317;
    wire N__3314;
    wire N__3311;
    wire N__3308;
    wire N__3305;
    wire N__3302;
    wire N__3299;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3279;
    wire N__3276;
    wire N__3273;
    wire N__3270;
    wire N__3267;
    wire N__3264;
    wire N__3261;
    wire N__3260;
    wire N__3257;
    wire N__3254;
    wire N__3251;
    wire N__3248;
    wire N__3245;
    wire N__3242;
    wire N__3239;
    wire N__3236;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3222;
    wire N__3219;
    wire N__3216;
    wire N__3213;
    wire N__3210;
    wire N__3207;
    wire N__3204;
    wire N__3201;
    wire N__3198;
    wire N__3195;
    wire N__3192;
    wire N__3189;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3171;
    wire N__3168;
    wire N__3165;
    wire N__3162;
    wire N__3159;
    wire N__3156;
    wire N__3153;
    wire N__3150;
    wire N__3147;
    wire N__3144;
    wire N__3141;
    wire N__3138;
    wire N__3135;
    wire N__3132;
    wire N__3131;
    wire N__3128;
    wire N__3125;
    wire N__3122;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3104;
    wire N__3101;
    wire N__3098;
    wire N__3095;
    wire N__3092;
    wire N__3089;
    wire N__3084;
    wire N__3081;
    wire N__3078;
    wire N__3075;
    wire N__3072;
    wire N__3069;
    wire N__3066;
    wire N__3063;
    wire N__3060;
    wire N__3057;
    wire N__3054;
    wire N__3051;
    wire N__3048;
    wire N__3045;
    wire N__3042;
    wire N__3039;
    wire N__3036;
    wire N__3033;
    wire N__3030;
    wire N__3027;
    wire N__3024;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3011;
    wire N__3008;
    wire N__3005;
    wire N__3002;
    wire N__2999;
    wire N__2996;
    wire N__2993;
    wire N__2990;
    wire N__2985;
    wire N__2982;
    wire N__2979;
    wire N__2976;
    wire N__2973;
    wire N__2970;
    wire N__2967;
    wire N__2964;
    wire N__2961;
    wire N__2958;
    wire N__2955;
    wire N__2952;
    wire N__2949;
    wire N__2946;
    wire N__2943;
    wire N__2940;
    wire N__2937;
    wire N__2934;
    wire N__2931;
    wire N__2928;
    wire N__2925;
    wire N__2922;
    wire N__2919;
    wire N__2916;
    wire N__2915;
    wire N__2912;
    wire N__2909;
    wire N__2906;
    wire N__2903;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2886;
    wire N__2883;
    wire N__2880;
    wire N__2877;
    wire N__2874;
    wire N__2871;
    wire N__2868;
    wire N__2865;
    wire N__2862;
    wire N__2859;
    wire N__2856;
    wire N__2853;
    wire N__2850;
    wire N__2847;
    wire N__2844;
    wire N__2843;
    wire N__2840;
    wire N__2837;
    wire N__2834;
    wire N__2831;
    wire N__2826;
    wire N__2823;
    wire N__2820;
    wire N__2817;
    wire N__2814;
    wire N__2811;
    wire N__2808;
    wire N__2805;
    wire N__2802;
    wire N__2799;
    wire N__2796;
    wire N__2793;
    wire N__2790;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2778;
    wire N__2775;
    wire N__2772;
    wire N__2769;
    wire N__2766;
    wire N__2763;
    wire N__2760;
    wire N__2757;
    wire N__2754;
    wire N__2751;
    wire N__2748;
    wire N__2745;
    wire N__2742;
    wire N__2739;
    wire N__2736;
    wire N__2733;
    wire N__2730;
    wire N__2727;
    wire N__2724;
    wire N__2721;
    wire N__2718;
    wire N__2715;
    wire N__2712;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2700;
    wire N__2697;
    wire N__2694;
    wire N__2691;
    wire N__2688;
    wire N__2685;
    wire N__2682;
    wire N__2679;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2667;
    wire N__2664;
    wire N__2661;
    wire N__2658;
    wire N__2655;
    wire N__2652;
    wire N__2649;
    wire N__2646;
    wire N__2643;
    wire N__2640;
    wire N__2637;
    wire N__2634;
    wire N__2631;
    wire N__2628;
    wire N__2625;
    wire N__2622;
    wire N__2619;
    wire N__2616;
    wire N__2613;
    wire N__2610;
    wire N__2607;
    wire N__2604;
    wire N__2601;
    wire N__2598;
    wire N__2595;
    wire TCIn_c;
    wire TSn_in;
    wire GNDG0;
    wire VCCG0;
    wire TAn_in;
    wire RESETn_c_i;
    wire U111_CYCLE_SM_A_AMIGA_0_i_1;
    wire A_040_c_0;
    wire A_AMIGA_c_0;
    wire D_LL_AMIGA_in_4;
    wire un2_D_LL_AMIGA_4;
    wire D_LL_AMIGA_in_1;
    wire un2_D_LL_AMIGA_1;
    wire D_UM_040_in_0;
    wire D_LL_040_in_0;
    wire un1_D_UM_040_0;
    wire D_LM_AMIGA_in_3;
    wire N_119;
    wire D_LM_AMIGA_in_1;
    wire N_121;
    wire D_LL_040_in_6;
    wire D_UM_040_in_6;
    wire un1_D_UM_040_6;
    wire D_LM_AMIGA_in_2;
    wire N_120;
    wire D_LM_040_in_0;
    wire D_UU_040_in_0;
    wire un1_D_UU_040_0;
    wire D_UU_040_in_4;
    wire D_LM_040_in_4;
    wire un1_D_UU_040_4;
    wire D_UU_040_in_6;
    wire D_LM_040_in_6;
    wire un1_D_UU_040_6;
    wire D_LL_AMIGA_in_2;
    wire un2_D_LL_AMIGA_2;
    wire D_LL_AMIGA_in_3;
    wire un2_D_LL_AMIGA_3;
    wire A_040_c_1;
    wire D_LM_AMIGA_in_0;
    wire N_122;
    wire \U111_CYCLE_SM.A2_ENZ0 ;
    wire \U111_CYCLE_SM.N_151 ;
    wire D_UM_040_in_1;
    wire D_LL_040_in_1;
    wire un1_D_UM_040_1;
    wire D_LL_040_in_3;
    wire D_UM_040_in_3;
    wire un1_D_UM_040_3;
    wire D_LM_AMIGA_in_7;
    wire N_115;
    wire D_UU_AMIGA_in_2;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ;
    wire N_129;
    wire D_UU_040_in_2;
    wire D_LM_040_in_2;
    wire un1_D_UU_040_2;
    wire CPUBGn_c_i_0;
    wire D_LL_AMIGA_in_7;
    wire un2_D_LL_AMIGA_7;
    wire \U111_CYCLE_SM.N_112_cascade_ ;
    wire \U111_CYCLE_SM.N_144_cascade_ ;
    wire \U111_CYCLE_SM.N_142 ;
    wire \U111_CYCLE_SM.N_197 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ;
    wire \U111_CYCLE_SM.N_195_cascade_ ;
    wire \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_1_0 ;
    wire TBIn_c;
    wire \U111_CYCLE_SM.BURSTZ0 ;
    wire \U111_CYCLE_SM.BURST_COUNTZ0Z_0 ;
    wire \U111_CYCLE_SM.BURST_COUNTZ0Z_1 ;
    wire \U111_CYCLE_SM.N_109 ;
    wire \U111_CYCLE_SM.N_109_cascade_ ;
    wire \U111_CYCLE_SM.PORT_MISMATCHZ0 ;
    wire D_LM_AMIGA_in_5;
    wire N_117;
    wire D_LM_AMIGA_in_4;
    wire N_118;
    wire D_UM_AMIGA_in_1;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ;
    wire un1_D_UM_AMIGA_1;
    wire D_LM_AMIGA_in_6;
    wire N_116;
    wire N_102_i;
    wire BUFDIR_c;
    wire BBn_c;
    wire N_104;
    wire D_UU_AMIGA_in_3;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ;
    wire N_128;
    wire \U111_CYCLE_SM.N_195 ;
    wire \U111_CYCLE_SM.N_132 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ;
    wire \U111_CYCLE_SM.TS_ENZ0 ;
    wire TS_OUT;
    wire \INVU111_CYCLE_SM.TS_OUTC_net ;
    wire PORTSIZE_c;
    wire U111_CYCLE_SM_OFFBOARD_EN_0;
    wire \U111_CYCLE_SM.un4_TS_OUT_i_0_cascade_ ;
    wire \U111_CYCLE_SM.N_106 ;
    wire RESETn_c;
    wire \U111_CYCLE_SM.N_140 ;
    wire \U111_CYCLE_SM.N_107 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ;
    wire TACKn_in;
    wire \U111_CYCLE_SM.LATCH_EN_5 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ;
    wire \U111_CYCLE_SM.N_57 ;
    wire D_UM_AMIGA_in_7;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ;
    wire un1_D_UM_AMIGA_7;
    wire GB_BUFFER_CLK40_THRU_CO;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ;
    wire D_UU_AMIGA_in_6;
    wire N_124;
    wire D_UU_AMIGA_in_5;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ;
    wire N_126;
    wire D_UU_AMIGA_in_7;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ;
    wire N_123;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ;
    wire D_UU_AMIGA_in_4;
    wire N_127;
    wire TEAn_c;
    wire U111_CYCLE_SM_TEA_CPUn_0_i;
    wire D_UU_040_in_1;
    wire D_LM_040_in_1;
    wire un1_D_UU_040_1;
    wire D_UM_040_in_7;
    wire D_LL_040_in_7;
    wire un1_D_UM_040_7;
    wire D_UM_AMIGA_in_3;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ;
    wire un1_D_UM_AMIGA_3;
    wire D_LL_040_in_4;
    wire D_UM_040_in_4;
    wire un1_D_UM_040_4;
    wire D_LL_AMIGA_in_6;
    wire un2_D_LL_AMIGA_6;
    wire D_LL_AMIGA_in_5;
    wire un2_D_LL_AMIGA_5;
    wire TS_CPUn_in;
    wire \U111_CYCLE_SM.TS_DELAYZ0 ;
    wire \U111_CYCLE_SM.un4_TS_OUT_i_0 ;
    wire \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0 ;
    wire \U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ;
    wire \U111_CYCLE_SM.N_107_i ;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ;
    wire \U111_CYCLE_SM.LW_TRANSZ0 ;
    wire CLK40;
    wire RESETn_c_i_g;
    wire D_UU_AMIGA_in_1;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ;
    wire N_130;
    wire \U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ;
    wire D_UU_AMIGA_in_0;
    wire N_131;
    wire \U111_CYCLE_SM.TA_DISZ0 ;
    wire N_66;
    wire D_UM_AMIGA_in_5;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ;
    wire un1_D_UM_AMIGA_5;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ;
    wire D_UM_AMIGA_in_4;
    wire un1_D_UM_AMIGA_4;
    wire D_UU_040_in_5;
    wire D_LM_040_in_5;
    wire un1_D_UU_040_5;
    wire LBENn_c;
    wire LBENn_c_i;
    wire D_LL_AMIGA_in_0;
    wire un2_D_LL_AMIGA_0;
    wire \U111_CYCLE_SM.CYCLE_ENZ0 ;
    wire BGn_c;
    wire CPUBGn_c;
    wire \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ;
    wire CPUBGn_c_cascade_;
    wire RnW_c;
    wire N_62_i;
    wire D_UM_AMIGA_in_2;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ;
    wire un1_D_UM_AMIGA_2;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ;
    wire D_UM_AMIGA_in_0;
    wire un1_D_UM_AMIGA_0;
    wire \U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ;
    wire D_UM_AMIGA_in_6;
    wire \U111_CYCLE_SM.LATCH_ENZ0 ;
    wire N_125;
    wire D_LL_040_in_2;
    wire D_UM_040_in_2;
    wire un1_D_UM_040_2;
    wire CLK80;
    wire GB_BUFFER_CLK80_THRU_CO;
    wire D_UU_040_in_3;
    wire D_LM_040_in_3;
    wire un1_D_UU_040_3;
    wire D_UU_040_in_7;
    wire D_LM_040_in_7;
    wire un1_D_UU_040_7;
    wire CONSTANT_ONE_NET;
    wire D_LL_040_in_5;
    wire D_UM_040_in_5;
    wire \U111_CYCLE_SM.FLIP_WORDZ0 ;
    wire un1_D_UM_040_5;
    wire _gnd_net_;

    defparam pll_pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll_pll.TEST_MODE=1'b0;
    defparam pll_pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll_pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll_pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll_pll.FILTER_RANGE=3'b011;
    defparam pll_pll.FEEDBACK_PATH="SIMPLE";
    defparam pll_pll.FDA_RELATIVE=4'b0000;
    defparam pll_pll.FDA_FEEDBACK=4'b0000;
    defparam pll_pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll_pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll_pll.DIVR=4'b0000;
    defparam pll_pll.DIVQ=3'b011;
    defparam pll_pll.DIVF=7'b0001111;
    defparam pll_pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40_2F pll_pll (
            .SCLK(),
            .PLLOUTGLOBALA(CLK80),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALB(CLK40),
            .SDI(),
            .PLLOUTCOREA(),
            .BYPASS(),
            .RESETB(N__7998),
            .PLLOUTCOREB(),
            .LOCK(),
            .SDO(),
            .EXTFEEDBACK(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__9464));
    IO_PAD pll_iopad (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__9464),
            .PACKAGEPIN(CLK40_IN));
    IO_PAD LBENn_ibuf_iopad (
            .OE(N__9448),
            .DIN(N__9447),
            .DOUT(N__9446),
            .PACKAGEPIN(LBENn));
    defparam LBENn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam LBENn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO LBENn_ibuf_preio (
            .PADOEN(N__9448),
            .PADOUT(N__9447),
            .PADIN(N__9446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(LBENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_3_iopad (
            .OE(N__9439),
            .DIN(N__9438),
            .DOUT(N__9437),
            .PACKAGEPIN(D_UM_040[3]));
    defparam D_UM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_3_preio (
            .PADOEN(N__9439),
            .PADOUT(N__9438),
            .PADIN(N__9437),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7010),
            .DIN0(D_UM_040_in_3),
            .DOUT0(N__6015),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TAn_iobuf_iopad (
            .OE(N__9430),
            .DIN(N__9429),
            .DOUT(N__9428),
            .PACKAGEPIN(TAn));
    defparam TAn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TAn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TAn_iobuf_preio (
            .PADOEN(N__9430),
            .PADOUT(N__9429),
            .PADIN(N__9428),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6105),
            .DIN0(TAn_in),
            .DOUT0(N__4548),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_1_iopad (
            .OE(N__9421),
            .DIN(N__9420),
            .DOUT(N__9419),
            .PACKAGEPIN(D_LL_AMIGA[1]));
    defparam D_LL_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_1_preio (
            .PADOEN(N__9421),
            .PADOUT(N__9420),
            .PADIN(N__9419),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4910),
            .DIN0(D_LL_AMIGA_in_1),
            .DOUT0(N__3341),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_5_iopad (
            .OE(N__9412),
            .DIN(N__9411),
            .DOUT(N__9410),
            .PACKAGEPIN(D_UU_AMIGA[5]));
    defparam D_UU_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_5_preio (
            .PADOEN(N__9412),
            .PADOUT(N__9411),
            .PADIN(N__9410),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4931),
            .DIN0(D_UU_AMIGA_in_5),
            .DOUT0(N__7470),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_6_iopad (
            .OE(N__9403),
            .DIN(N__9402),
            .DOUT(N__9401),
            .PACKAGEPIN(D_UU_040[6]));
    defparam D_UU_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_6_preio (
            .PADOEN(N__9403),
            .PADOUT(N__9402),
            .PADIN(N__9401),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6973),
            .DIN0(D_UU_040_in_6),
            .DOUT0(N__5649),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CPUBGn_obuf_iopad (
            .OE(N__9394),
            .DIN(N__9393),
            .DOUT(N__9392),
            .PACKAGEPIN(CPUBGn));
    defparam CPUBGn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUBGn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CPUBGn_obuf_preio (
            .PADOEN(N__9394),
            .PADOUT(N__9393),
            .PADIN(N__9392),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7272),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_7_iopad (
            .OE(N__9385),
            .DIN(N__9384),
            .DOUT(N__9383),
            .PACKAGEPIN(D_LL_040[7]));
    defparam D_LL_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_7_preio (
            .PADOEN(N__9385),
            .PADOUT(N__9384),
            .PADIN(N__9383),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6850),
            .DIN0(D_LL_040_in_7),
            .DOUT0(N__3567),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_4_iopad (
            .OE(N__9376),
            .DIN(N__9375),
            .DOUT(N__9374),
            .PACKAGEPIN(D_LL_AMIGA[4]));
    defparam D_LL_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_4_preio (
            .PADOEN(N__9376),
            .PADOUT(N__9375),
            .PADIN(N__9374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4909),
            .DIN0(D_LL_AMIGA_in_4),
            .DOUT0(N__5999),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_3_iopad (
            .OE(N__9367),
            .DIN(N__9366),
            .DOUT(N__9365),
            .PACKAGEPIN(D_UM_AMIGA[3]));
    defparam D_UM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_3_preio (
            .PADOEN(N__9367),
            .PADOUT(N__9366),
            .PADIN(N__9365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4918),
            .DIN0(D_UM_AMIGA_in_3),
            .DOUT0(N__3816),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_3_iopad (
            .OE(N__9358),
            .DIN(N__9357),
            .DOUT(N__9356),
            .PACKAGEPIN(D_UU_040[3]));
    defparam D_UU_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_3_preio (
            .PADOEN(N__9358),
            .PADOUT(N__9357),
            .PADIN(N__9356),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7004),
            .DIN0(D_UU_040_in_3),
            .DOUT0(N__4158),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TEA_CPUn_obuf_iopad (
            .OE(N__9349),
            .DIN(N__9348),
            .DOUT(N__9347),
            .PACKAGEPIN(TEA_CPUn));
    defparam TEA_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TEA_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TEA_CPUn_obuf_preio (
            .PADOEN(N__9349),
            .PADOUT(N__9348),
            .PADIN(N__9347),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5310),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_1_iopad (
            .OE(N__9340),
            .DIN(N__9339),
            .DOUT(N__9338),
            .PACKAGEPIN(A_040[1]));
    defparam A_040_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_1_preio (
            .PADOEN(N__9340),
            .PADOUT(N__9339),
            .PADIN(N__9338),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_3_iopad (
            .OE(N__9331),
            .DIN(N__9330),
            .DOUT(N__9329),
            .PACKAGEPIN(D_LM_AMIGA[3]));
    defparam D_LM_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_3_preio (
            .PADOEN(N__9331),
            .PADOUT(N__9330),
            .PADIN(N__9329),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4708),
            .DIN0(D_LM_AMIGA_in_3),
            .DOUT0(N__8139),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_0_iopad (
            .OE(N__9322),
            .DIN(N__9321),
            .DOUT(N__9320),
            .PACKAGEPIN(D_LM_040[0]));
    defparam D_LM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_0_preio (
            .PADOEN(N__9322),
            .PADOUT(N__9321),
            .PADIN(N__9320),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6851),
            .DIN0(D_LM_040_in_0),
            .DOUT0(N__3429),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_6_iopad (
            .OE(N__9313),
            .DIN(N__9312),
            .DOUT(N__9311),
            .PACKAGEPIN(D_UM_AMIGA[6]));
    defparam D_UM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_6_preio (
            .PADOEN(N__9313),
            .PADOUT(N__9312),
            .PADIN(N__9311),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4930),
            .DIN0(D_UM_AMIGA_in_6),
            .DOUT0(N__3069),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_4_iopad (
            .OE(N__9304),
            .DIN(N__9303),
            .DOUT(N__9302),
            .PACKAGEPIN(D_LM_AMIGA[4]));
    defparam D_LM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_4_preio (
            .PADOEN(N__9304),
            .PADOUT(N__9303),
            .PADIN(N__9302),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4840),
            .DIN0(D_LM_AMIGA_in_4),
            .DOUT0(N__2925),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_1_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_1_iopad (
            .OE(N__9295),
            .DIN(N__9294),
            .DOUT(N__9293),
            .PACKAGEPIN(A_AMIGA[1]));
    defparam A_AMIGA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_1_preio (
            .PADOEN(N__9295),
            .PADOUT(N__9294),
            .PADIN(N__9293),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2760),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_7_iopad (
            .OE(N__9286),
            .DIN(N__9285),
            .DOUT(N__9284),
            .PACKAGEPIN(D_LM_040[7]));
    defparam D_LM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_7_preio (
            .PADOEN(N__9286),
            .PADOUT(N__9285),
            .PADIN(N__9284),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6970),
            .DIN0(D_LM_040_in_7),
            .DOUT0(N__3780),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_4_iopad (
            .OE(N__9277),
            .DIN(N__9276),
            .DOUT(N__9275),
            .PACKAGEPIN(D_UM_040[4]));
    defparam D_UM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_4_preio (
            .PADOEN(N__9277),
            .PADOUT(N__9276),
            .PADIN(N__9275),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7005),
            .DIN0(D_UM_040_in_4),
            .DOUT0(N__7542),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_obuf_iopad (
            .OE(N__9268),
            .DIN(N__9267),
            .DOUT(N__9266),
            .PACKAGEPIN(CLK40B));
    defparam CLK40B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_obuf_preio (
            .PADOEN(N__9268),
            .PADOUT(N__9267),
            .PADIN(N__9266),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5764),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_0_iopad (
            .OE(N__9259),
            .DIN(N__9258),
            .DOUT(N__9257),
            .PACKAGEPIN(D_UU_AMIGA[0]));
    defparam D_UU_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_0_preio (
            .PADOEN(N__9259),
            .PADOUT(N__9258),
            .PADIN(N__9257),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4878),
            .DIN0(D_UU_AMIGA_in_0),
            .DOUT0(N__2964),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_1_iopad (
            .OE(N__9250),
            .DIN(N__9249),
            .DOUT(N__9248),
            .PACKAGEPIN(D_UM_040[1]));
    defparam D_UM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_1_preio (
            .PADOEN(N__9250),
            .PADOUT(N__9249),
            .PADIN(N__9248),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6849),
            .DIN0(D_UM_040_in_1),
            .DOUT0(N__4347),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_ibuf_iopad (
            .OE(N__9241),
            .DIN(N__9240),
            .DOUT(N__9239),
            .PACKAGEPIN(TBIn));
    defparam TBIn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TBIn_ibuf_preio (
            .PADOEN(N__9241),
            .PADOUT(N__9240),
            .PADIN(N__9239),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TBIn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_4_iopad (
            .OE(N__9232),
            .DIN(N__9231),
            .DOUT(N__9230),
            .PACKAGEPIN(D_LL_040[4]));
    defparam D_LL_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_4_preio (
            .PADOEN(N__9232),
            .PADOUT(N__9231),
            .PADIN(N__9230),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6909),
            .DIN0(D_LL_040_in_4),
            .DOUT0(N__2706),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_7_iopad (
            .OE(N__9223),
            .DIN(N__9222),
            .DOUT(N__9221),
            .PACKAGEPIN(D_LL_AMIGA[7]));
    defparam D_LL_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_7_preio (
            .PADOEN(N__9223),
            .PADOUT(N__9222),
            .PADIN(N__9221),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4863),
            .DIN0(D_LL_AMIGA_in_7),
            .DOUT0(N__5199),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_7_iopad (
            .OE(N__9214),
            .DIN(N__9213),
            .DOUT(N__9212),
            .PACKAGEPIN(D_UU_AMIGA[7]));
    defparam D_UU_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_7_preio (
            .PADOEN(N__9214),
            .PADOUT(N__9213),
            .PADIN(N__9212),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4914),
            .DIN0(D_UU_AMIGA_in_7),
            .DOUT0(N__8013),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFDIR_obuf_iopad (
            .OE(N__9205),
            .DIN(N__9204),
            .DOUT(N__9203),
            .PACKAGEPIN(BUFDIR));
    defparam BUFDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFDIR_obuf_preio (
            .PADOEN(N__9205),
            .PADOUT(N__9204),
            .PADIN(N__9203),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4284),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_4_iopad (
            .OE(N__9196),
            .DIN(N__9195),
            .DOUT(N__9194),
            .PACKAGEPIN(D_UU_040[4]));
    defparam D_UU_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_4_preio (
            .PADOEN(N__9196),
            .PADOUT(N__9195),
            .PADIN(N__9194),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6936),
            .DIN0(D_UU_040_in_4),
            .DOUT0(N__5406),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__9187),
            .DIN(N__9186),
            .DOUT(N__9185),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__9187),
            .PADOUT(N__9186),
            .PADIN(N__9185),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_1_iopad (
            .OE(N__9178),
            .DIN(N__9177),
            .DOUT(N__9176),
            .PACKAGEPIN(D_LL_040[1]));
    defparam D_LL_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_1_preio (
            .PADOEN(N__9178),
            .PADOUT(N__9177),
            .PADIN(N__9176),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6908),
            .DIN0(D_LL_040_in_1),
            .DOUT0(N__2673),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_5_iopad (
            .OE(N__9169),
            .DIN(N__9168),
            .DOUT(N__9167),
            .PACKAGEPIN(D_UM_AMIGA[5]));
    defparam D_UM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_5_preio (
            .PADOEN(N__9169),
            .PADOUT(N__9168),
            .PADIN(N__9167),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4879),
            .DIN0(D_UM_AMIGA_in_5),
            .DOUT0(N__8574),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_1_iopad (
            .OE(N__9160),
            .DIN(N__9159),
            .DOUT(N__9158),
            .PACKAGEPIN(D_UU_040[1]));
    defparam D_UU_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_1_preio (
            .PADOEN(N__9160),
            .PADOUT(N__9159),
            .PADIN(N__9158),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7011),
            .DIN0(D_UU_040_in_1),
            .DOUT0(N__6243),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_1_iopad (
            .OE(N__9151),
            .DIN(N__9150),
            .DOUT(N__9149),
            .PACKAGEPIN(D_LM_AMIGA[1]));
    defparam D_LM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_1_preio (
            .PADOEN(N__9151),
            .PADOUT(N__9150),
            .PADIN(N__9149),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4775),
            .DIN0(D_LM_AMIGA_in_1),
            .DOUT0(N__5277),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_2_iopad (
            .OE(N__9142),
            .DIN(N__9141),
            .DOUT(N__9140),
            .PACKAGEPIN(D_LM_040[2]));
    defparam D_LM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_2_preio (
            .PADOEN(N__9142),
            .PADOUT(N__9141),
            .PADIN(N__9140),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6860),
            .DIN0(D_LM_040_in_2),
            .DOUT0(N__3045),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__9133),
            .DIN(N__9132),
            .DOUT(N__9131),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__9133),
            .PADOUT(N__9132),
            .PADIN(N__9131),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7374),
            .DIN0(TACKn_in),
            .DOUT0(N__2793),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_2_iopad (
            .OE(N__9124),
            .DIN(N__9123),
            .DOUT(N__9122),
            .PACKAGEPIN(D_UM_040[2]));
    defparam D_UM_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_2_preio (
            .PADOEN(N__9124),
            .PADOUT(N__9123),
            .PADIN(N__9122),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6924),
            .DIN0(D_UM_040_in_2),
            .DOUT0(N__6663),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMB_obuf_iopad (
            .OE(N__9115),
            .DIN(N__9114),
            .DOUT(N__9113),
            .PACKAGEPIN(CLKRAMB));
    defparam CLKRAMB_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMB_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMB_obuf_preio (
            .PADOEN(N__9115),
            .PADOUT(N__9114),
            .PADIN(N__9113),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8189),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_2_iopad (
            .OE(N__9106),
            .DIN(N__9105),
            .DOUT(N__9104),
            .PACKAGEPIN(D_LL_AMIGA[2]));
    defparam D_LL_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_2_preio (
            .PADOEN(N__9106),
            .PADOUT(N__9105),
            .PADIN(N__9104),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4735),
            .DIN0(D_LL_AMIGA_in_2),
            .DOUT0(N__8283),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_2_iopad (
            .OE(N__9097),
            .DIN(N__9096),
            .DOUT(N__9095),
            .PACKAGEPIN(D_UU_AMIGA[2]));
    defparam D_UU_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_2_preio (
            .PADOEN(N__9097),
            .PADOUT(N__9096),
            .PADIN(N__9095),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4877),
            .DIN0(D_UU_AMIGA_in_2),
            .DOUT0(N__3609),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TEAn_ibuf_iopad (
            .OE(N__9088),
            .DIN(N__9087),
            .DOUT(N__9086),
            .PACKAGEPIN(TEAn));
    defparam TEAn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TEAn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TEAn_ibuf_preio (
            .PADOEN(N__9088),
            .PADOUT(N__9087),
            .PADIN(N__9086),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TEAn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__9079),
            .DIN(N__9078),
            .DOUT(N__9077),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__9079),
            .PADOUT(N__9078),
            .PADIN(N__9077),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4296),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_6_iopad (
            .OE(N__9070),
            .DIN(N__9069),
            .DOUT(N__9068),
            .PACKAGEPIN(D_LL_040[6]));
    defparam D_LL_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_6_preio (
            .PADOEN(N__9070),
            .PADOUT(N__9069),
            .PADIN(N__9068),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6961),
            .DIN0(D_LL_040_in_6),
            .DOUT0(N__5901),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_5_iopad (
            .OE(N__9061),
            .DIN(N__9060),
            .DOUT(N__9059),
            .PACKAGEPIN(D_LL_AMIGA[5]));
    defparam D_LL_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_5_preio (
            .PADOEN(N__9061),
            .PADOUT(N__9060),
            .PADIN(N__9059),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4866),
            .DIN0(D_LL_AMIGA_in_5),
            .DOUT0(N__7983),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_0_iopad (
            .OE(N__9052),
            .DIN(N__9051),
            .DOUT(N__9050),
            .PACKAGEPIN(D_UM_AMIGA[0]));
    defparam D_UM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_0_preio (
            .PADOEN(N__9052),
            .PADOUT(N__9051),
            .PADIN(N__9050),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4839),
            .DIN0(D_UM_AMIGA_in_0),
            .DOUT0(N__3222),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_2_iopad (
            .OE(N__9043),
            .DIN(N__9042),
            .DOUT(N__9041),
            .PACKAGEPIN(D_UU_040[2]));
    defparam D_UU_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_2_preio (
            .PADOEN(N__9043),
            .PADOUT(N__9042),
            .PADIN(N__9041),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6852),
            .DIN0(D_UU_040_in_2),
            .DOUT0(N__3696),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_iobuf_iopad (
            .OE(N__9034),
            .DIN(N__9033),
            .DOUT(N__9032),
            .PACKAGEPIN(TSn));
    defparam TSn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TSn_iobuf_preio (
            .PADOEN(N__9034),
            .PADOUT(N__9033),
            .PADIN(N__9032),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3591),
            .DIN0(TSn_in),
            .DOUT0(N__4098),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_2_iopad (
            .OE(N__9025),
            .DIN(N__9024),
            .DOUT(N__9023),
            .PACKAGEPIN(D_LM_AMIGA[2]));
    defparam D_LM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_2_preio (
            .PADOEN(N__9025),
            .PADOUT(N__9024),
            .PADIN(N__9023),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4838),
            .DIN0(D_LM_AMIGA_in_2),
            .DOUT0(N__3651),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TS_CPUn_iobuf_iopad (
            .OE(N__9016),
            .DIN(N__9015),
            .DOUT(N__9014),
            .PACKAGEPIN(TS_CPUn));
    defparam TS_CPUn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TS_CPUn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TS_CPUn_iobuf_preio (
            .PADOEN(N__9016),
            .PADOUT(N__9015),
            .PADIN(N__9014),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7271),
            .DIN0(TS_CPUn_in),
            .DOUT0(N__2649),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK80_CPU_obuf_iopad (
            .OE(N__9007),
            .DIN(N__9006),
            .DOUT(N__9005),
            .PACKAGEPIN(CLK80_CPU));
    defparam CLK80_CPU_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK80_CPU_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK80_CPU_obuf_preio (
            .PADOEN(N__9007),
            .PADOUT(N__9006),
            .PADIN(N__9005),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8193),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_3_iopad (
            .OE(N__8998),
            .DIN(N__8997),
            .DOUT(N__8996),
            .PACKAGEPIN(D_LL_040[3]));
    defparam D_LL_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_3_preio (
            .PADOEN(N__8998),
            .PADOUT(N__8997),
            .PADIN(N__8996),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6994),
            .DIN0(D_LL_040_in_3),
            .DOUT0(N__3495),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_1_iopad (
            .OE(N__8989),
            .DIN(N__8988),
            .DOUT(N__8987),
            .PACKAGEPIN(D_LM_040[1]));
    defparam D_LM_040_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_1_preio (
            .PADOEN(N__8989),
            .PADOUT(N__8988),
            .PADIN(N__8987),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6859),
            .DIN0(D_LM_040_in_1),
            .DOUT0(N__3156),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_7_iopad (
            .OE(N__8980),
            .DIN(N__8979),
            .DOUT(N__8978),
            .PACKAGEPIN(D_UM_AMIGA[7]));
    defparam D_UM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_7_preio (
            .PADOEN(N__8980),
            .PADOUT(N__8979),
            .PADIN(N__8978),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4916),
            .DIN0(D_UM_AMIGA_in_7),
            .DOUT0(N__5151),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_7_iopad (
            .OE(N__8971),
            .DIN(N__8970),
            .DOUT(N__8969),
            .PACKAGEPIN(D_LM_AMIGA[7]));
    defparam D_LM_AMIGA_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_7_preio (
            .PADOEN(N__8971),
            .PADOUT(N__8970),
            .PADIN(N__8969),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4891),
            .DIN0(D_LM_AMIGA_in_7),
            .DOUT0(N__8055),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_ibuf_iopad (
            .OE(N__8962),
            .DIN(N__8961),
            .DOUT(N__8960),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PORTSIZE_ibuf_preio (
            .PADOEN(N__8962),
            .PADOUT(N__8961),
            .PADIN(N__8960),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PORTSIZE_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_AMIGA_obuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_AMIGA_obuf_0_iopad (
            .OE(N__8953),
            .DIN(N__8952),
            .DOUT(N__8951),
            .PACKAGEPIN(A_AMIGA[0]));
    defparam A_AMIGA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_AMIGA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO A_AMIGA_obuf_0_preio (
            .PADOEN(N__8953),
            .PADOUT(N__8952),
            .PADIN(N__8951),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2736),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_4_iopad (
            .OE(N__8944),
            .DIN(N__8943),
            .DOUT(N__8942),
            .PACKAGEPIN(D_LM_040[4]));
    defparam D_LM_040_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_4_preio (
            .PADOEN(N__8944),
            .PADOUT(N__8943),
            .PADIN(N__8942),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6927),
            .DIN0(D_LM_040_in_4),
            .DOUT0(N__4431),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_7_iopad (
            .OE(N__8935),
            .DIN(N__8934),
            .DOUT(N__8933),
            .PACKAGEPIN(D_UM_040[7]));
    defparam D_UM_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_7_preio (
            .PADOEN(N__8935),
            .PADOUT(N__8934),
            .PADIN(N__8933),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7009),
            .DIN0(D_UM_040_in_7),
            .DOUT0(N__4998),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__8926),
            .DIN(N__8925),
            .DOUT(N__8924),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__8926),
            .PADOUT(N__8925),
            .PADIN(N__8924),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_1_iopad (
            .OE(N__8917),
            .DIN(N__8916),
            .DOUT(N__8915),
            .PACKAGEPIN(D_UU_AMIGA[1]));
    defparam D_UU_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_1_preio (
            .PADOEN(N__8917),
            .PADOUT(N__8916),
            .PADIN(N__8915),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4917),
            .DIN0(D_UU_AMIGA_in_1),
            .DOUT0(N__5235),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__8908),
            .DIN(N__8907),
            .DOUT(N__8906),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__8908),
            .PADOUT(N__8907),
            .PADIN(N__8906),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5754),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_0_iopad (
            .OE(N__8899),
            .DIN(N__8898),
            .DOUT(N__8897),
            .PACKAGEPIN(D_UM_040[0]));
    defparam D_UM_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_0_preio (
            .PADOEN(N__8899),
            .PADOUT(N__8898),
            .PADIN(N__8897),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6925),
            .DIN0(D_UM_040_in_0),
            .DOUT0(N__8499),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_0_iopad (
            .OE(N__8890),
            .DIN(N__8889),
            .DOUT(N__8888),
            .PACKAGEPIN(D_LL_AMIGA[0]));
    defparam D_LL_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_0_preio (
            .PADOEN(N__8890),
            .PADOUT(N__8889),
            .PADIN(N__8888),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4929),
            .DIN0(D_LL_AMIGA_in_0),
            .DOUT0(N__3264),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_4_iopad (
            .OE(N__8881),
            .DIN(N__8880),
            .DOUT(N__8879),
            .PACKAGEPIN(D_UU_AMIGA[4]));
    defparam D_UU_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_4_preio (
            .PADOEN(N__8881),
            .PADOUT(N__8880),
            .PADIN(N__8879),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4876),
            .DIN0(D_UU_AMIGA_in_4),
            .DOUT0(N__2886),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_7_iopad (
            .OE(N__8872),
            .DIN(N__8871),
            .DOUT(N__8870),
            .PACKAGEPIN(D_UU_040[7]));
    defparam D_UU_040_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_7_preio (
            .PADOEN(N__8872),
            .PADOUT(N__8871),
            .PADIN(N__8870),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6972),
            .DIN0(D_UU_040_in_7),
            .DOUT0(N__5490),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__8863),
            .DIN(N__8862),
            .DOUT(N__8861),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__8863),
            .PADOUT(N__8862),
            .PADIN(N__8861),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BGn_ibuf_iopad (
            .OE(N__8854),
            .DIN(N__8853),
            .DOUT(N__8852),
            .PACKAGEPIN(BGn));
    defparam BGn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BGn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BGn_ibuf_preio (
            .PADOEN(N__8854),
            .PADOUT(N__8853),
            .PADIN(N__8852),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BGn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_0_iopad (
            .OE(N__8845),
            .DIN(N__8844),
            .DOUT(N__8843),
            .PACKAGEPIN(D_LL_040[0]));
    defparam D_LL_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_0_preio (
            .PADOEN(N__8845),
            .PADOUT(N__8844),
            .PADIN(N__8843),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6995),
            .DIN0(D_LL_040_in_0),
            .DOUT0(N__7347),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_2_iopad (
            .OE(N__8836),
            .DIN(N__8835),
            .DOUT(N__8834),
            .PACKAGEPIN(D_UM_AMIGA[2]));
    defparam D_UM_AMIGA_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_2_preio (
            .PADOEN(N__8836),
            .PADOUT(N__8835),
            .PADIN(N__8834),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4841),
            .DIN0(D_UM_AMIGA_in_2),
            .DOUT0(N__8226),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_0_iopad (
            .OE(N__8827),
            .DIN(N__8826),
            .DOUT(N__8825),
            .PACKAGEPIN(D_UU_040[0]));
    defparam D_UU_040_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_0_preio (
            .PADOEN(N__8827),
            .PADOUT(N__8826),
            .PADIN(N__8825),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6971),
            .DIN0(D_UU_040_in_0),
            .DOUT0(N__6159),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_ibuf_iopad (
            .OE(N__8818),
            .DIN(N__8817),
            .DOUT(N__8816),
            .PACKAGEPIN(TCIn));
    defparam TCIn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TCIn_ibuf_preio (
            .PADOEN(N__8818),
            .PADOUT(N__8817),
            .PADIN(N__8816),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TCIn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_040_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_040_ibuf_0_iopad (
            .OE(N__8809),
            .DIN(N__8808),
            .DOUT(N__8807),
            .PACKAGEPIN(A_040[0]));
    defparam A_040_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_040_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_040_ibuf_0_preio (
            .PADOEN(N__8809),
            .PADOUT(N__8808),
            .PADIN(N__8807),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_040_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_0_iopad (
            .OE(N__8800),
            .DIN(N__8799),
            .DOUT(N__8798),
            .PACKAGEPIN(D_LM_AMIGA[0]));
    defparam D_LM_AMIGA_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_0_preio (
            .PADOEN(N__8800),
            .PADOUT(N__8799),
            .PADIN(N__8798),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4864),
            .DIN0(D_LM_AMIGA_in_0),
            .DOUT0(N__3030),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBI_CPUn_obuf_iopad (
            .OE(N__8791),
            .DIN(N__8790),
            .DOUT(N__8789),
            .PACKAGEPIN(TBI_CPUn));
    defparam TBI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TBI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TBI_CPUn_obuf_preio (
            .PADOEN(N__8791),
            .PADOUT(N__8790),
            .PADIN(N__8789),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4070),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40A_obuf_iopad (
            .OE(N__8782),
            .DIN(N__8781),
            .DOUT(N__8780),
            .PACKAGEPIN(CLK40A));
    defparam CLK40A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40A_obuf_preio (
            .PADOEN(N__8782),
            .PADOUT(N__8781),
            .PADIN(N__8780),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5768),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_3_iopad (
            .OE(N__8773),
            .DIN(N__8772),
            .DOUT(N__8771),
            .PACKAGEPIN(D_LM_040[3]));
    defparam D_LM_040_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_3_preio (
            .PADOEN(N__8773),
            .PADOUT(N__8772),
            .PADIN(N__8771),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6969),
            .DIN0(D_LM_040_in_3),
            .DOUT0(N__3189),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_5_iopad (
            .OE(N__8764),
            .DIN(N__8763),
            .DOUT(N__8762),
            .PACKAGEPIN(D_LM_AMIGA[5]));
    defparam D_LM_AMIGA_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_5_preio (
            .PADOEN(N__8764),
            .PADOUT(N__8763),
            .PADIN(N__8762),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4889),
            .DIN0(D_LM_AMIGA_in_5),
            .DOUT0(N__7506),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_6_iopad (
            .OE(N__8755),
            .DIN(N__8754),
            .DOUT(N__8753),
            .PACKAGEPIN(D_LM_040[6]));
    defparam D_LM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_6_preio (
            .PADOEN(N__8755),
            .PADOUT(N__8754),
            .PADIN(N__8753),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6932),
            .DIN0(D_LM_040_in_6),
            .DOUT0(N__4308),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_5_iopad (
            .OE(N__8746),
            .DIN(N__8745),
            .DOUT(N__8744),
            .PACKAGEPIN(D_UM_040[5]));
    defparam D_UM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_5_preio (
            .PADOEN(N__8746),
            .PADOUT(N__8745),
            .PADIN(N__8744),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6996),
            .DIN0(D_UM_040_in_5),
            .DOUT0(N__7635),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_3_iopad (
            .OE(N__8737),
            .DIN(N__8736),
            .DOUT(N__8735),
            .PACKAGEPIN(D_LL_AMIGA[3]));
    defparam D_LL_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_3_preio (
            .PADOEN(N__8737),
            .PADOUT(N__8736),
            .PADIN(N__8735),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4734),
            .DIN0(D_LL_AMIGA_in_3),
            .DOUT0(N__3878),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_3_iopad (
            .OE(N__8728),
            .DIN(N__8727),
            .DOUT(N__8726),
            .PACKAGEPIN(D_UU_AMIGA[3]));
    defparam D_UU_AMIGA_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_3_preio (
            .PADOEN(N__8728),
            .PADOUT(N__8727),
            .PADIN(N__8726),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4932),
            .DIN0(D_UU_AMIGA_in_3),
            .DOUT0(N__8094),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_5_iopad (
            .OE(N__8719),
            .DIN(N__8718),
            .DOUT(N__8717),
            .PACKAGEPIN(D_LL_040[5]));
    defparam D_LL_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_5_preio (
            .PADOEN(N__8719),
            .PADOUT(N__8718),
            .PADIN(N__8717),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6960),
            .DIN0(D_LL_040_in_5),
            .DOUT0(N__5862),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_AMIGA_iobuf_6_iopad (
            .OE(N__8710),
            .DIN(N__8709),
            .DOUT(N__8708),
            .PACKAGEPIN(D_LL_AMIGA[6]));
    defparam D_LL_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_AMIGA_iobuf_6_preio (
            .PADOEN(N__8710),
            .PADOUT(N__8709),
            .PADIN(N__8708),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4865),
            .DIN0(D_LL_AMIGA_in_6),
            .DOUT0(N__3135),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_AMIGA_iobuf_6_iopad (
            .OE(N__8701),
            .DIN(N__8700),
            .DOUT(N__8699),
            .PACKAGEPIN(D_UU_AMIGA[6]));
    defparam D_UU_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_AMIGA_iobuf_6_preio (
            .PADOEN(N__8701),
            .PADOUT(N__8700),
            .PADIN(N__8699),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4915),
            .DIN0(D_UU_AMIGA_in_6),
            .DOUT0(N__2811),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_1_iopad (
            .OE(N__8692),
            .DIN(N__8691),
            .DOUT(N__8690),
            .PACKAGEPIN(D_UM_AMIGA[1]));
    defparam D_UM_AMIGA_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_1_preio (
            .PADOEN(N__8692),
            .PADOUT(N__8691),
            .PADIN(N__8690),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4890),
            .DIN0(D_UM_AMIGA_in_1),
            .DOUT0(N__3294),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UU_040_iobuf_5_iopad (
            .OE(N__8683),
            .DIN(N__8682),
            .DOUT(N__8681),
            .PACKAGEPIN(D_UU_040[5]));
    defparam D_UU_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_UU_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UU_040_iobuf_5_preio (
            .PADOEN(N__8683),
            .PADOUT(N__8682),
            .PADIN(N__8681),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6997),
            .DIN0(D_UU_040_in_5),
            .DOUT0(N__5565),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAMA_obuf_iopad (
            .OE(N__8674),
            .DIN(N__8673),
            .DOUT(N__8672),
            .PACKAGEPIN(CLKRAMA));
    defparam CLKRAMA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAMA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAMA_obuf_preio (
            .PADOEN(N__8674),
            .PADOUT(N__8673),
            .PADIN(N__8672),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5772),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LL_040_iobuf_2_iopad (
            .OE(N__8665),
            .DIN(N__8664),
            .DOUT(N__8663),
            .PACKAGEPIN(D_LL_040[2]));
    defparam D_LL_040_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam D_LL_040_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LL_040_iobuf_2_preio (
            .PADOEN(N__8665),
            .PADOUT(N__8664),
            .PADIN(N__8663),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6962),
            .DIN0(D_LL_040_in_2),
            .DOUT0(N__3534),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCI_CPUn_obuf_iopad (
            .OE(N__8656),
            .DIN(N__8655),
            .DOUT(N__8654),
            .PACKAGEPIN(TCI_CPUn));
    defparam TCI_CPUn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TCI_CPUn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TCI_CPUn_obuf_preio (
            .PADOEN(N__8656),
            .PADOUT(N__8655),
            .PADIN(N__8654),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2622),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BBn_ibuf_iopad (
            .OE(N__8647),
            .DIN(N__8646),
            .DOUT(N__8645),
            .PACKAGEPIN(BBn));
    defparam BBn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BBn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BBn_ibuf_preio (
            .PADOEN(N__8647),
            .PADOUT(N__8646),
            .PADIN(N__8645),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BBn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMAAn_obuf_iopad (
            .OE(N__8638),
            .DIN(N__8637),
            .DOUT(N__8636),
            .PACKAGEPIN(DMAAn));
    defparam DMAAn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMAAn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMAAn_obuf_preio (
            .PADOEN(N__8638),
            .PADOUT(N__8637),
            .PADIN(N__8636),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4245),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_AMIGA_iobuf_4_iopad (
            .OE(N__8629),
            .DIN(N__8628),
            .DOUT(N__8627),
            .PACKAGEPIN(D_UM_AMIGA[4]));
    defparam D_UM_AMIGA_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_AMIGA_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_AMIGA_iobuf_4_preio (
            .PADOEN(N__8629),
            .PADOUT(N__8628),
            .PADIN(N__8627),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4919),
            .DIN0(D_UM_AMIGA_in_4),
            .DOUT0(N__5937),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_AMIGA_iobuf_6_iopad (
            .OE(N__8620),
            .DIN(N__8619),
            .DOUT(N__8618),
            .PACKAGEPIN(D_LM_AMIGA[6]));
    defparam D_LM_AMIGA_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_AMIGA_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_AMIGA_iobuf_6_preio (
            .PADOEN(N__8620),
            .PADOUT(N__8619),
            .PADIN(N__8618),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4892),
            .DIN0(D_LM_AMIGA_in_6),
            .DOUT0(N__2850),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__8611),
            .DIN(N__8610),
            .DOUT(N__8609),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__8611),
            .PADOUT(N__8610),
            .PADIN(N__8609),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_LM_040_iobuf_5_iopad (
            .OE(N__8602),
            .DIN(N__8601),
            .DOUT(N__8600),
            .PACKAGEPIN(D_LM_040[5]));
    defparam D_LM_040_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_LM_040_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_LM_040_iobuf_5_preio (
            .PADOEN(N__8602),
            .PADOUT(N__8601),
            .PADIN(N__8600),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6926),
            .DIN0(D_LM_040_in_5),
            .DOUT0(N__3957),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_UM_040_iobuf_6_iopad (
            .OE(N__8593),
            .DIN(N__8592),
            .DOUT(N__8591),
            .PACKAGEPIN(D_UM_040[6]));
    defparam D_UM_040_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_UM_040_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_UM_040_iobuf_6_preio (
            .PADOEN(N__8593),
            .PADOUT(N__8592),
            .PADIN(N__8591),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6931),
            .DIN0(D_UM_040_in_6),
            .DOUT0(N__8304),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__2213 (
            .O(N__8574),
            .I(N__8571));
    LocalMux I__2212 (
            .O(N__8571),
            .I(N__8568));
    IoSpan4Mux I__2211 (
            .O(N__8568),
            .I(N__8565));
    Sp12to4 I__2210 (
            .O(N__8565),
            .I(N__8562));
    Span12Mux_s6_v I__2209 (
            .O(N__8562),
            .I(N__8559));
    Odrv12 I__2208 (
            .O(N__8559),
            .I(un1_D_UM_040_5));
    InMux I__2207 (
            .O(N__8556),
            .I(N__8552));
    InMux I__2206 (
            .O(N__8555),
            .I(N__8549));
    LocalMux I__2205 (
            .O(N__8552),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ));
    LocalMux I__2204 (
            .O(N__8549),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ));
    InMux I__2203 (
            .O(N__8544),
            .I(N__8541));
    LocalMux I__2202 (
            .O(N__8541),
            .I(N__8537));
    CascadeMux I__2201 (
            .O(N__8540),
            .I(N__8534));
    Span4Mux_v I__2200 (
            .O(N__8537),
            .I(N__8531));
    InMux I__2199 (
            .O(N__8534),
            .I(N__8528));
    Span4Mux_v I__2198 (
            .O(N__8531),
            .I(N__8523));
    LocalMux I__2197 (
            .O(N__8528),
            .I(N__8523));
    Span4Mux_v I__2196 (
            .O(N__8523),
            .I(N__8520));
    Span4Mux_h I__2195 (
            .O(N__8520),
            .I(N__8516));
    InMux I__2194 (
            .O(N__8519),
            .I(N__8513));
    Span4Mux_h I__2193 (
            .O(N__8516),
            .I(N__8510));
    LocalMux I__2192 (
            .O(N__8513),
            .I(N__8507));
    Sp12to4 I__2191 (
            .O(N__8510),
            .I(N__8502));
    Span12Mux_h I__2190 (
            .O(N__8507),
            .I(N__8502));
    Odrv12 I__2189 (
            .O(N__8502),
            .I(D_UM_AMIGA_in_0));
    IoInMux I__2188 (
            .O(N__8499),
            .I(N__8496));
    LocalMux I__2187 (
            .O(N__8496),
            .I(N__8493));
    IoSpan4Mux I__2186 (
            .O(N__8493),
            .I(N__8490));
    Span4Mux_s2_h I__2185 (
            .O(N__8490),
            .I(N__8487));
    Sp12to4 I__2184 (
            .O(N__8487),
            .I(N__8484));
    Span12Mux_s11_h I__2183 (
            .O(N__8484),
            .I(N__8481));
    Odrv12 I__2182 (
            .O(N__8481),
            .I(un1_D_UM_AMIGA_0));
    InMux I__2181 (
            .O(N__8478),
            .I(N__8474));
    InMux I__2180 (
            .O(N__8477),
            .I(N__8471));
    LocalMux I__2179 (
            .O(N__8474),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ));
    LocalMux I__2178 (
            .O(N__8471),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ));
    InMux I__2177 (
            .O(N__8466),
            .I(N__8462));
    CascadeMux I__2176 (
            .O(N__8465),
            .I(N__8459));
    LocalMux I__2175 (
            .O(N__8462),
            .I(N__8456));
    InMux I__2174 (
            .O(N__8459),
            .I(N__8453));
    Span4Mux_v I__2173 (
            .O(N__8456),
            .I(N__8447));
    LocalMux I__2172 (
            .O(N__8453),
            .I(N__8447));
    InMux I__2171 (
            .O(N__8452),
            .I(N__8444));
    Span4Mux_v I__2170 (
            .O(N__8447),
            .I(N__8441));
    LocalMux I__2169 (
            .O(N__8444),
            .I(N__8436));
    Sp12to4 I__2168 (
            .O(N__8441),
            .I(N__8436));
    Span12Mux_h I__2167 (
            .O(N__8436),
            .I(N__8433));
    Span12Mux_v I__2166 (
            .O(N__8433),
            .I(N__8430));
    Odrv12 I__2165 (
            .O(N__8430),
            .I(D_UM_AMIGA_in_6));
    InMux I__2164 (
            .O(N__8427),
            .I(N__8416));
    InMux I__2163 (
            .O(N__8426),
            .I(N__8416));
    InMux I__2162 (
            .O(N__8425),
            .I(N__8411));
    InMux I__2161 (
            .O(N__8424),
            .I(N__8411));
    InMux I__2160 (
            .O(N__8423),
            .I(N__8408));
    InMux I__2159 (
            .O(N__8422),
            .I(N__8405));
    InMux I__2158 (
            .O(N__8421),
            .I(N__8398));
    LocalMux I__2157 (
            .O(N__8416),
            .I(N__8393));
    LocalMux I__2156 (
            .O(N__8411),
            .I(N__8390));
    LocalMux I__2155 (
            .O(N__8408),
            .I(N__8385));
    LocalMux I__2154 (
            .O(N__8405),
            .I(N__8385));
    InMux I__2153 (
            .O(N__8404),
            .I(N__8382));
    InMux I__2152 (
            .O(N__8403),
            .I(N__8375));
    InMux I__2151 (
            .O(N__8402),
            .I(N__8375));
    InMux I__2150 (
            .O(N__8401),
            .I(N__8375));
    LocalMux I__2149 (
            .O(N__8398),
            .I(N__8372));
    InMux I__2148 (
            .O(N__8397),
            .I(N__8369));
    InMux I__2147 (
            .O(N__8396),
            .I(N__8366));
    Span4Mux_v I__2146 (
            .O(N__8393),
            .I(N__8360));
    Span4Mux_h I__2145 (
            .O(N__8390),
            .I(N__8351));
    Span4Mux_v I__2144 (
            .O(N__8385),
            .I(N__8351));
    LocalMux I__2143 (
            .O(N__8382),
            .I(N__8351));
    LocalMux I__2142 (
            .O(N__8375),
            .I(N__8351));
    Span4Mux_v I__2141 (
            .O(N__8372),
            .I(N__8346));
    LocalMux I__2140 (
            .O(N__8369),
            .I(N__8346));
    LocalMux I__2139 (
            .O(N__8366),
            .I(N__8343));
    InMux I__2138 (
            .O(N__8365),
            .I(N__8338));
    InMux I__2137 (
            .O(N__8364),
            .I(N__8338));
    CascadeMux I__2136 (
            .O(N__8363),
            .I(N__8334));
    Span4Mux_v I__2135 (
            .O(N__8360),
            .I(N__8331));
    Span4Mux_v I__2134 (
            .O(N__8351),
            .I(N__8328));
    Span4Mux_v I__2133 (
            .O(N__8346),
            .I(N__8321));
    Span4Mux_v I__2132 (
            .O(N__8343),
            .I(N__8321));
    LocalMux I__2131 (
            .O(N__8338),
            .I(N__8321));
    InMux I__2130 (
            .O(N__8337),
            .I(N__8318));
    InMux I__2129 (
            .O(N__8334),
            .I(N__8315));
    Odrv4 I__2128 (
            .O(N__8331),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    Odrv4 I__2127 (
            .O(N__8328),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    Odrv4 I__2126 (
            .O(N__8321),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    LocalMux I__2125 (
            .O(N__8318),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    LocalMux I__2124 (
            .O(N__8315),
            .I(\U111_CYCLE_SM.LATCH_ENZ0 ));
    IoInMux I__2123 (
            .O(N__8304),
            .I(N__8301));
    LocalMux I__2122 (
            .O(N__8301),
            .I(N__8298));
    IoSpan4Mux I__2121 (
            .O(N__8298),
            .I(N__8295));
    Span4Mux_s0_h I__2120 (
            .O(N__8295),
            .I(N__8292));
    Sp12to4 I__2119 (
            .O(N__8292),
            .I(N__8289));
    Span12Mux_s7_h I__2118 (
            .O(N__8289),
            .I(N__8286));
    Odrv12 I__2117 (
            .O(N__8286),
            .I(N_125));
    IoInMux I__2116 (
            .O(N__8283),
            .I(N__8280));
    LocalMux I__2115 (
            .O(N__8280),
            .I(N__8276));
    InMux I__2114 (
            .O(N__8279),
            .I(N__8273));
    IoSpan4Mux I__2113 (
            .O(N__8276),
            .I(N__8270));
    LocalMux I__2112 (
            .O(N__8273),
            .I(N__8267));
    Span4Mux_s2_h I__2111 (
            .O(N__8270),
            .I(N__8264));
    Span4Mux_v I__2110 (
            .O(N__8267),
            .I(N__8261));
    Sp12to4 I__2109 (
            .O(N__8264),
            .I(N__8258));
    Sp12to4 I__2108 (
            .O(N__8261),
            .I(N__8255));
    Span12Mux_h I__2107 (
            .O(N__8258),
            .I(N__8252));
    Span12Mux_h I__2106 (
            .O(N__8255),
            .I(N__8249));
    Span12Mux_h I__2105 (
            .O(N__8252),
            .I(N__8246));
    Span12Mux_v I__2104 (
            .O(N__8249),
            .I(N__8243));
    Odrv12 I__2103 (
            .O(N__8246),
            .I(D_LL_040_in_2));
    Odrv12 I__2102 (
            .O(N__8243),
            .I(D_LL_040_in_2));
    InMux I__2101 (
            .O(N__8238),
            .I(N__8235));
    LocalMux I__2100 (
            .O(N__8235),
            .I(N__8232));
    Span12Mux_h I__2099 (
            .O(N__8232),
            .I(N__8229));
    Odrv12 I__2098 (
            .O(N__8229),
            .I(D_UM_040_in_2));
    IoInMux I__2097 (
            .O(N__8226),
            .I(N__8223));
    LocalMux I__2096 (
            .O(N__8223),
            .I(N__8220));
    Span4Mux_s3_h I__2095 (
            .O(N__8220),
            .I(N__8217));
    Sp12to4 I__2094 (
            .O(N__8217),
            .I(N__8214));
    Span12Mux_v I__2093 (
            .O(N__8214),
            .I(N__8211));
    Span12Mux_h I__2092 (
            .O(N__8211),
            .I(N__8208));
    Odrv12 I__2091 (
            .O(N__8208),
            .I(un1_D_UM_040_2));
    InMux I__2090 (
            .O(N__8205),
            .I(N__8202));
    LocalMux I__2089 (
            .O(N__8202),
            .I(N__8199));
    Glb2LocalMux I__2088 (
            .O(N__8199),
            .I(N__8196));
    GlobalMux I__2087 (
            .O(N__8196),
            .I(CLK80));
    IoInMux I__2086 (
            .O(N__8193),
            .I(N__8190));
    LocalMux I__2085 (
            .O(N__8190),
            .I(N__8186));
    IoInMux I__2084 (
            .O(N__8189),
            .I(N__8183));
    IoSpan4Mux I__2083 (
            .O(N__8186),
            .I(N__8180));
    LocalMux I__2082 (
            .O(N__8183),
            .I(N__8177));
    Sp12to4 I__2081 (
            .O(N__8180),
            .I(N__8174));
    Span12Mux_s3_v I__2080 (
            .O(N__8177),
            .I(N__8171));
    Span12Mux_s7_h I__2079 (
            .O(N__8174),
            .I(N__8168));
    Span12Mux_v I__2078 (
            .O(N__8171),
            .I(N__8165));
    Odrv12 I__2077 (
            .O(N__8168),
            .I(GB_BUFFER_CLK80_THRU_CO));
    Odrv12 I__2076 (
            .O(N__8165),
            .I(GB_BUFFER_CLK80_THRU_CO));
    InMux I__2075 (
            .O(N__8160),
            .I(N__8157));
    LocalMux I__2074 (
            .O(N__8157),
            .I(N__8154));
    Span4Mux_v I__2073 (
            .O(N__8154),
            .I(N__8151));
    Span4Mux_h I__2072 (
            .O(N__8151),
            .I(N__8148));
    Sp12to4 I__2071 (
            .O(N__8148),
            .I(N__8145));
    Span12Mux_h I__2070 (
            .O(N__8145),
            .I(N__8142));
    Odrv12 I__2069 (
            .O(N__8142),
            .I(D_UU_040_in_3));
    IoInMux I__2068 (
            .O(N__8139),
            .I(N__8136));
    LocalMux I__2067 (
            .O(N__8136),
            .I(N__8133));
    IoSpan4Mux I__2066 (
            .O(N__8133),
            .I(N__8129));
    InMux I__2065 (
            .O(N__8132),
            .I(N__8126));
    IoSpan4Mux I__2064 (
            .O(N__8129),
            .I(N__8123));
    LocalMux I__2063 (
            .O(N__8126),
            .I(N__8120));
    Span4Mux_s2_h I__2062 (
            .O(N__8123),
            .I(N__8117));
    Span4Mux_v I__2061 (
            .O(N__8120),
            .I(N__8114));
    Sp12to4 I__2060 (
            .O(N__8117),
            .I(N__8111));
    Sp12to4 I__2059 (
            .O(N__8114),
            .I(N__8108));
    Span12Mux_h I__2058 (
            .O(N__8111),
            .I(N__8105));
    Span12Mux_h I__2057 (
            .O(N__8108),
            .I(N__8102));
    Span12Mux_h I__2056 (
            .O(N__8105),
            .I(N__8097));
    Span12Mux_v I__2055 (
            .O(N__8102),
            .I(N__8097));
    Odrv12 I__2054 (
            .O(N__8097),
            .I(D_LM_040_in_3));
    IoInMux I__2053 (
            .O(N__8094),
            .I(N__8091));
    LocalMux I__2052 (
            .O(N__8091),
            .I(N__8088));
    Span4Mux_s2_v I__2051 (
            .O(N__8088),
            .I(N__8085));
    Span4Mux_v I__2050 (
            .O(N__8085),
            .I(N__8082));
    Sp12to4 I__2049 (
            .O(N__8082),
            .I(N__8079));
    Span12Mux_s11_h I__2048 (
            .O(N__8079),
            .I(N__8076));
    Odrv12 I__2047 (
            .O(N__8076),
            .I(un1_D_UU_040_3));
    InMux I__2046 (
            .O(N__8073),
            .I(N__8070));
    LocalMux I__2045 (
            .O(N__8070),
            .I(N__8067));
    Span4Mux_v I__2044 (
            .O(N__8067),
            .I(N__8064));
    Sp12to4 I__2043 (
            .O(N__8064),
            .I(N__8061));
    Span12Mux_h I__2042 (
            .O(N__8061),
            .I(N__8058));
    Odrv12 I__2041 (
            .O(N__8058),
            .I(D_UU_040_in_7));
    IoInMux I__2040 (
            .O(N__8055),
            .I(N__8052));
    LocalMux I__2039 (
            .O(N__8052),
            .I(N__8049));
    IoSpan4Mux I__2038 (
            .O(N__8049),
            .I(N__8045));
    InMux I__2037 (
            .O(N__8048),
            .I(N__8042));
    Span4Mux_s2_h I__2036 (
            .O(N__8045),
            .I(N__8039));
    LocalMux I__2035 (
            .O(N__8042),
            .I(N__8036));
    Sp12to4 I__2034 (
            .O(N__8039),
            .I(N__8033));
    Span4Mux_v I__2033 (
            .O(N__8036),
            .I(N__8030));
    Span12Mux_h I__2032 (
            .O(N__8033),
            .I(N__8027));
    Sp12to4 I__2031 (
            .O(N__8030),
            .I(N__8024));
    Span12Mux_h I__2030 (
            .O(N__8027),
            .I(N__8021));
    Span12Mux_h I__2029 (
            .O(N__8024),
            .I(N__8018));
    Odrv12 I__2028 (
            .O(N__8021),
            .I(D_LM_040_in_7));
    Odrv12 I__2027 (
            .O(N__8018),
            .I(D_LM_040_in_7));
    IoInMux I__2026 (
            .O(N__8013),
            .I(N__8010));
    LocalMux I__2025 (
            .O(N__8010),
            .I(N__8007));
    Span12Mux_s8_v I__2024 (
            .O(N__8007),
            .I(N__8004));
    Span12Mux_h I__2023 (
            .O(N__8004),
            .I(N__8001));
    Odrv12 I__2022 (
            .O(N__8001),
            .I(un1_D_UU_040_7));
    IoInMux I__2021 (
            .O(N__7998),
            .I(N__7995));
    LocalMux I__2020 (
            .O(N__7995),
            .I(N__7992));
    Span4Mux_s2_v I__2019 (
            .O(N__7992),
            .I(N__7989));
    Span4Mux_v I__2018 (
            .O(N__7989),
            .I(N__7986));
    Odrv4 I__2017 (
            .O(N__7986),
            .I(CONSTANT_ONE_NET));
    IoInMux I__2016 (
            .O(N__7983),
            .I(N__7980));
    LocalMux I__2015 (
            .O(N__7980),
            .I(N__7977));
    IoSpan4Mux I__2014 (
            .O(N__7977),
            .I(N__7973));
    InMux I__2013 (
            .O(N__7976),
            .I(N__7970));
    Span4Mux_s2_h I__2012 (
            .O(N__7973),
            .I(N__7967));
    LocalMux I__2011 (
            .O(N__7970),
            .I(N__7964));
    Span4Mux_v I__2010 (
            .O(N__7967),
            .I(N__7961));
    Sp12to4 I__2009 (
            .O(N__7964),
            .I(N__7958));
    Sp12to4 I__2008 (
            .O(N__7961),
            .I(N__7955));
    Span12Mux_v I__2007 (
            .O(N__7958),
            .I(N__7952));
    Span12Mux_h I__2006 (
            .O(N__7955),
            .I(N__7947));
    Span12Mux_v I__2005 (
            .O(N__7952),
            .I(N__7947));
    Span12Mux_h I__2004 (
            .O(N__7947),
            .I(N__7944));
    Odrv12 I__2003 (
            .O(N__7944),
            .I(D_LL_040_in_5));
    InMux I__2002 (
            .O(N__7941),
            .I(N__7938));
    LocalMux I__2001 (
            .O(N__7938),
            .I(N__7935));
    Span4Mux_v I__2000 (
            .O(N__7935),
            .I(N__7932));
    Sp12to4 I__1999 (
            .O(N__7932),
            .I(N__7929));
    Span12Mux_h I__1998 (
            .O(N__7929),
            .I(N__7926));
    Odrv12 I__1997 (
            .O(N__7926),
            .I(D_UM_040_in_5));
    InMux I__1996 (
            .O(N__7923),
            .I(N__7910));
    InMux I__1995 (
            .O(N__7922),
            .I(N__7910));
    InMux I__1994 (
            .O(N__7921),
            .I(N__7910));
    InMux I__1993 (
            .O(N__7920),
            .I(N__7904));
    InMux I__1992 (
            .O(N__7919),
            .I(N__7904));
    InMux I__1991 (
            .O(N__7918),
            .I(N__7898));
    InMux I__1990 (
            .O(N__7917),
            .I(N__7890));
    LocalMux I__1989 (
            .O(N__7910),
            .I(N__7887));
    InMux I__1988 (
            .O(N__7909),
            .I(N__7884));
    LocalMux I__1987 (
            .O(N__7904),
            .I(N__7880));
    InMux I__1986 (
            .O(N__7903),
            .I(N__7877));
    InMux I__1985 (
            .O(N__7902),
            .I(N__7872));
    InMux I__1984 (
            .O(N__7901),
            .I(N__7872));
    LocalMux I__1983 (
            .O(N__7898),
            .I(N__7868));
    InMux I__1982 (
            .O(N__7897),
            .I(N__7861));
    InMux I__1981 (
            .O(N__7896),
            .I(N__7861));
    InMux I__1980 (
            .O(N__7895),
            .I(N__7861));
    InMux I__1979 (
            .O(N__7894),
            .I(N__7856));
    InMux I__1978 (
            .O(N__7893),
            .I(N__7856));
    LocalMux I__1977 (
            .O(N__7890),
            .I(N__7853));
    Span4Mux_v I__1976 (
            .O(N__7887),
            .I(N__7847));
    LocalMux I__1975 (
            .O(N__7884),
            .I(N__7844));
    InMux I__1974 (
            .O(N__7883),
            .I(N__7841));
    Span4Mux_v I__1973 (
            .O(N__7880),
            .I(N__7834));
    LocalMux I__1972 (
            .O(N__7877),
            .I(N__7834));
    LocalMux I__1971 (
            .O(N__7872),
            .I(N__7831));
    InMux I__1970 (
            .O(N__7871),
            .I(N__7828));
    Span4Mux_v I__1969 (
            .O(N__7868),
            .I(N__7825));
    LocalMux I__1968 (
            .O(N__7861),
            .I(N__7822));
    LocalMux I__1967 (
            .O(N__7856),
            .I(N__7819));
    Span4Mux_v I__1966 (
            .O(N__7853),
            .I(N__7814));
    InMux I__1965 (
            .O(N__7852),
            .I(N__7809));
    InMux I__1964 (
            .O(N__7851),
            .I(N__7809));
    InMux I__1963 (
            .O(N__7850),
            .I(N__7802));
    Span4Mux_h I__1962 (
            .O(N__7847),
            .I(N__7795));
    Span4Mux_v I__1961 (
            .O(N__7844),
            .I(N__7795));
    LocalMux I__1960 (
            .O(N__7841),
            .I(N__7795));
    InMux I__1959 (
            .O(N__7840),
            .I(N__7790));
    InMux I__1958 (
            .O(N__7839),
            .I(N__7790));
    Span4Mux_v I__1957 (
            .O(N__7834),
            .I(N__7787));
    Span4Mux_h I__1956 (
            .O(N__7831),
            .I(N__7782));
    LocalMux I__1955 (
            .O(N__7828),
            .I(N__7782));
    Span4Mux_h I__1954 (
            .O(N__7825),
            .I(N__7777));
    Span4Mux_v I__1953 (
            .O(N__7822),
            .I(N__7777));
    Span4Mux_v I__1952 (
            .O(N__7819),
            .I(N__7774));
    InMux I__1951 (
            .O(N__7818),
            .I(N__7769));
    InMux I__1950 (
            .O(N__7817),
            .I(N__7769));
    Span4Mux_h I__1949 (
            .O(N__7814),
            .I(N__7764));
    LocalMux I__1948 (
            .O(N__7809),
            .I(N__7764));
    InMux I__1947 (
            .O(N__7808),
            .I(N__7757));
    InMux I__1946 (
            .O(N__7807),
            .I(N__7757));
    InMux I__1945 (
            .O(N__7806),
            .I(N__7757));
    InMux I__1944 (
            .O(N__7805),
            .I(N__7754));
    LocalMux I__1943 (
            .O(N__7802),
            .I(N__7747));
    Span4Mux_v I__1942 (
            .O(N__7795),
            .I(N__7742));
    LocalMux I__1941 (
            .O(N__7790),
            .I(N__7742));
    Span4Mux_v I__1940 (
            .O(N__7787),
            .I(N__7737));
    Span4Mux_v I__1939 (
            .O(N__7782),
            .I(N__7737));
    Span4Mux_v I__1938 (
            .O(N__7777),
            .I(N__7730));
    Span4Mux_v I__1937 (
            .O(N__7774),
            .I(N__7730));
    LocalMux I__1936 (
            .O(N__7769),
            .I(N__7730));
    Sp12to4 I__1935 (
            .O(N__7764),
            .I(N__7723));
    LocalMux I__1934 (
            .O(N__7757),
            .I(N__7723));
    LocalMux I__1933 (
            .O(N__7754),
            .I(N__7723));
    InMux I__1932 (
            .O(N__7753),
            .I(N__7716));
    InMux I__1931 (
            .O(N__7752),
            .I(N__7716));
    InMux I__1930 (
            .O(N__7751),
            .I(N__7716));
    InMux I__1929 (
            .O(N__7750),
            .I(N__7713));
    Odrv12 I__1928 (
            .O(N__7747),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__1927 (
            .O(N__7742),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__1926 (
            .O(N__7737),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv4 I__1925 (
            .O(N__7730),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    Odrv12 I__1924 (
            .O(N__7723),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    LocalMux I__1923 (
            .O(N__7716),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    LocalMux I__1922 (
            .O(N__7713),
            .I(\U111_CYCLE_SM.FLIP_WORDZ0 ));
    InMux I__1921 (
            .O(N__7698),
            .I(N__7695));
    LocalMux I__1920 (
            .O(N__7695),
            .I(N__7691));
    CascadeMux I__1919 (
            .O(N__7694),
            .I(N__7688));
    Span4Mux_v I__1918 (
            .O(N__7691),
            .I(N__7685));
    InMux I__1917 (
            .O(N__7688),
            .I(N__7682));
    Span4Mux_v I__1916 (
            .O(N__7685),
            .I(N__7677));
    LocalMux I__1915 (
            .O(N__7682),
            .I(N__7677));
    Span4Mux_v I__1914 (
            .O(N__7677),
            .I(N__7674));
    Span4Mux_v I__1913 (
            .O(N__7674),
            .I(N__7671));
    Span4Mux_h I__1912 (
            .O(N__7671),
            .I(N__7667));
    InMux I__1911 (
            .O(N__7670),
            .I(N__7664));
    Sp12to4 I__1910 (
            .O(N__7667),
            .I(N__7659));
    LocalMux I__1909 (
            .O(N__7664),
            .I(N__7659));
    Span12Mux_h I__1908 (
            .O(N__7659),
            .I(N__7656));
    Odrv12 I__1907 (
            .O(N__7656),
            .I(D_UM_AMIGA_in_5));
    InMux I__1906 (
            .O(N__7653),
            .I(N__7650));
    LocalMux I__1905 (
            .O(N__7650),
            .I(N__7647));
    Span4Mux_v I__1904 (
            .O(N__7647),
            .I(N__7643));
    InMux I__1903 (
            .O(N__7646),
            .I(N__7640));
    Odrv4 I__1902 (
            .O(N__7643),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ));
    LocalMux I__1901 (
            .O(N__7640),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ));
    IoInMux I__1900 (
            .O(N__7635),
            .I(N__7632));
    LocalMux I__1899 (
            .O(N__7632),
            .I(N__7629));
    Span4Mux_s3_v I__1898 (
            .O(N__7629),
            .I(N__7626));
    Span4Mux_h I__1897 (
            .O(N__7626),
            .I(N__7623));
    Sp12to4 I__1896 (
            .O(N__7623),
            .I(N__7620));
    Span12Mux_s10_v I__1895 (
            .O(N__7620),
            .I(N__7617));
    Span12Mux_h I__1894 (
            .O(N__7617),
            .I(N__7614));
    Odrv12 I__1893 (
            .O(N__7614),
            .I(un1_D_UM_AMIGA_5));
    InMux I__1892 (
            .O(N__7611),
            .I(N__7608));
    LocalMux I__1891 (
            .O(N__7608),
            .I(N__7605));
    Span4Mux_v I__1890 (
            .O(N__7605),
            .I(N__7602));
    Span4Mux_v I__1889 (
            .O(N__7602),
            .I(N__7598));
    InMux I__1888 (
            .O(N__7601),
            .I(N__7595));
    Odrv4 I__1887 (
            .O(N__7598),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ));
    LocalMux I__1886 (
            .O(N__7595),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ));
    CascadeMux I__1885 (
            .O(N__7590),
            .I(N__7587));
    InMux I__1884 (
            .O(N__7587),
            .I(N__7582));
    InMux I__1883 (
            .O(N__7586),
            .I(N__7579));
    InMux I__1882 (
            .O(N__7585),
            .I(N__7576));
    LocalMux I__1881 (
            .O(N__7582),
            .I(N__7573));
    LocalMux I__1880 (
            .O(N__7579),
            .I(N__7570));
    LocalMux I__1879 (
            .O(N__7576),
            .I(N__7567));
    Span4Mux_h I__1878 (
            .O(N__7573),
            .I(N__7564));
    Span4Mux_v I__1877 (
            .O(N__7570),
            .I(N__7561));
    Span12Mux_v I__1876 (
            .O(N__7567),
            .I(N__7556));
    Sp12to4 I__1875 (
            .O(N__7564),
            .I(N__7556));
    Sp12to4 I__1874 (
            .O(N__7561),
            .I(N__7553));
    Span12Mux_v I__1873 (
            .O(N__7556),
            .I(N__7550));
    Span12Mux_h I__1872 (
            .O(N__7553),
            .I(N__7547));
    Odrv12 I__1871 (
            .O(N__7550),
            .I(D_UM_AMIGA_in_4));
    Odrv12 I__1870 (
            .O(N__7547),
            .I(D_UM_AMIGA_in_4));
    IoInMux I__1869 (
            .O(N__7542),
            .I(N__7539));
    LocalMux I__1868 (
            .O(N__7539),
            .I(N__7536));
    Span12Mux_s7_v I__1867 (
            .O(N__7536),
            .I(N__7533));
    Span12Mux_h I__1866 (
            .O(N__7533),
            .I(N__7530));
    Odrv12 I__1865 (
            .O(N__7530),
            .I(un1_D_UM_AMIGA_4));
    InMux I__1864 (
            .O(N__7527),
            .I(N__7524));
    LocalMux I__1863 (
            .O(N__7524),
            .I(N__7521));
    Span4Mux_h I__1862 (
            .O(N__7521),
            .I(N__7518));
    Sp12to4 I__1861 (
            .O(N__7518),
            .I(N__7515));
    Span12Mux_v I__1860 (
            .O(N__7515),
            .I(N__7512));
    Span12Mux_h I__1859 (
            .O(N__7512),
            .I(N__7509));
    Odrv12 I__1858 (
            .O(N__7509),
            .I(D_UU_040_in_5));
    IoInMux I__1857 (
            .O(N__7506),
            .I(N__7503));
    LocalMux I__1856 (
            .O(N__7503),
            .I(N__7500));
    IoSpan4Mux I__1855 (
            .O(N__7500),
            .I(N__7497));
    IoSpan4Mux I__1854 (
            .O(N__7497),
            .I(N__7494));
    Span4Mux_s2_h I__1853 (
            .O(N__7494),
            .I(N__7490));
    InMux I__1852 (
            .O(N__7493),
            .I(N__7487));
    Sp12to4 I__1851 (
            .O(N__7490),
            .I(N__7484));
    LocalMux I__1850 (
            .O(N__7487),
            .I(N__7481));
    Span12Mux_h I__1849 (
            .O(N__7484),
            .I(N__7476));
    Span12Mux_v I__1848 (
            .O(N__7481),
            .I(N__7476));
    Span12Mux_h I__1847 (
            .O(N__7476),
            .I(N__7473));
    Odrv12 I__1846 (
            .O(N__7473),
            .I(D_LM_040_in_5));
    IoInMux I__1845 (
            .O(N__7470),
            .I(N__7467));
    LocalMux I__1844 (
            .O(N__7467),
            .I(N__7464));
    IoSpan4Mux I__1843 (
            .O(N__7464),
            .I(N__7461));
    Span4Mux_s2_h I__1842 (
            .O(N__7461),
            .I(N__7458));
    Sp12to4 I__1841 (
            .O(N__7458),
            .I(N__7455));
    Span12Mux_h I__1840 (
            .O(N__7455),
            .I(N__7452));
    Odrv12 I__1839 (
            .O(N__7452),
            .I(un1_D_UU_040_5));
    InMux I__1838 (
            .O(N__7449),
            .I(N__7446));
    LocalMux I__1837 (
            .O(N__7446),
            .I(N__7442));
    InMux I__1836 (
            .O(N__7445),
            .I(N__7439));
    Span4Mux_v I__1835 (
            .O(N__7442),
            .I(N__7433));
    LocalMux I__1834 (
            .O(N__7439),
            .I(N__7433));
    CascadeMux I__1833 (
            .O(N__7438),
            .I(N__7430));
    Span4Mux_h I__1832 (
            .O(N__7433),
            .I(N__7427));
    InMux I__1831 (
            .O(N__7430),
            .I(N__7424));
    Span4Mux_v I__1830 (
            .O(N__7427),
            .I(N__7420));
    LocalMux I__1829 (
            .O(N__7424),
            .I(N__7417));
    InMux I__1828 (
            .O(N__7423),
            .I(N__7414));
    Span4Mux_v I__1827 (
            .O(N__7420),
            .I(N__7409));
    Span4Mux_h I__1826 (
            .O(N__7417),
            .I(N__7409));
    LocalMux I__1825 (
            .O(N__7414),
            .I(N__7405));
    Span4Mux_v I__1824 (
            .O(N__7409),
            .I(N__7402));
    InMux I__1823 (
            .O(N__7408),
            .I(N__7399));
    Span12Mux_h I__1822 (
            .O(N__7405),
            .I(N__7396));
    Span4Mux_v I__1821 (
            .O(N__7402),
            .I(N__7393));
    LocalMux I__1820 (
            .O(N__7399),
            .I(N__7390));
    Span12Mux_v I__1819 (
            .O(N__7396),
            .I(N__7387));
    Span4Mux_v I__1818 (
            .O(N__7393),
            .I(N__7384));
    Span4Mux_v I__1817 (
            .O(N__7390),
            .I(N__7381));
    Odrv12 I__1816 (
            .O(N__7387),
            .I(LBENn_c));
    Odrv4 I__1815 (
            .O(N__7384),
            .I(LBENn_c));
    Odrv4 I__1814 (
            .O(N__7381),
            .I(LBENn_c));
    IoInMux I__1813 (
            .O(N__7374),
            .I(N__7371));
    LocalMux I__1812 (
            .O(N__7371),
            .I(N__7368));
    Odrv12 I__1811 (
            .O(N__7368),
            .I(LBENn_c_i));
    InMux I__1810 (
            .O(N__7365),
            .I(N__7362));
    LocalMux I__1809 (
            .O(N__7362),
            .I(N__7359));
    Span4Mux_v I__1808 (
            .O(N__7359),
            .I(N__7356));
    Sp12to4 I__1807 (
            .O(N__7356),
            .I(N__7353));
    Span12Mux_h I__1806 (
            .O(N__7353),
            .I(N__7350));
    Odrv12 I__1805 (
            .O(N__7350),
            .I(D_LL_AMIGA_in_0));
    IoInMux I__1804 (
            .O(N__7347),
            .I(N__7344));
    LocalMux I__1803 (
            .O(N__7344),
            .I(N__7341));
    Span4Mux_s2_h I__1802 (
            .O(N__7341),
            .I(N__7338));
    Span4Mux_v I__1801 (
            .O(N__7338),
            .I(N__7335));
    Span4Mux_h I__1800 (
            .O(N__7335),
            .I(N__7332));
    Sp12to4 I__1799 (
            .O(N__7332),
            .I(N__7329));
    Span12Mux_h I__1798 (
            .O(N__7329),
            .I(N__7326));
    Odrv12 I__1797 (
            .O(N__7326),
            .I(un2_D_LL_AMIGA_0));
    InMux I__1796 (
            .O(N__7323),
            .I(N__7320));
    LocalMux I__1795 (
            .O(N__7320),
            .I(N__7315));
    InMux I__1794 (
            .O(N__7319),
            .I(N__7312));
    InMux I__1793 (
            .O(N__7318),
            .I(N__7309));
    Odrv12 I__1792 (
            .O(N__7315),
            .I(\U111_CYCLE_SM.CYCLE_ENZ0 ));
    LocalMux I__1791 (
            .O(N__7312),
            .I(\U111_CYCLE_SM.CYCLE_ENZ0 ));
    LocalMux I__1790 (
            .O(N__7309),
            .I(\U111_CYCLE_SM.CYCLE_ENZ0 ));
    InMux I__1789 (
            .O(N__7302),
            .I(N__7298));
    InMux I__1788 (
            .O(N__7301),
            .I(N__7295));
    LocalMux I__1787 (
            .O(N__7298),
            .I(N__7292));
    LocalMux I__1786 (
            .O(N__7295),
            .I(N__7289));
    Span4Mux_v I__1785 (
            .O(N__7292),
            .I(N__7286));
    Span4Mux_v I__1784 (
            .O(N__7289),
            .I(N__7283));
    Sp12to4 I__1783 (
            .O(N__7286),
            .I(N__7278));
    Sp12to4 I__1782 (
            .O(N__7283),
            .I(N__7278));
    Span12Mux_h I__1781 (
            .O(N__7278),
            .I(N__7275));
    Odrv12 I__1780 (
            .O(N__7275),
            .I(BGn_c));
    IoInMux I__1779 (
            .O(N__7272),
            .I(N__7268));
    IoInMux I__1778 (
            .O(N__7271),
            .I(N__7265));
    LocalMux I__1777 (
            .O(N__7268),
            .I(N__7262));
    LocalMux I__1776 (
            .O(N__7265),
            .I(N__7259));
    IoSpan4Mux I__1775 (
            .O(N__7262),
            .I(N__7253));
    IoSpan4Mux I__1774 (
            .O(N__7259),
            .I(N__7250));
    InMux I__1773 (
            .O(N__7258),
            .I(N__7247));
    InMux I__1772 (
            .O(N__7257),
            .I(N__7242));
    InMux I__1771 (
            .O(N__7256),
            .I(N__7242));
    Span4Mux_s2_h I__1770 (
            .O(N__7253),
            .I(N__7239));
    Span4Mux_s1_v I__1769 (
            .O(N__7250),
            .I(N__7236));
    LocalMux I__1768 (
            .O(N__7247),
            .I(N__7231));
    LocalMux I__1767 (
            .O(N__7242),
            .I(N__7231));
    Sp12to4 I__1766 (
            .O(N__7239),
            .I(N__7227));
    Span4Mux_v I__1765 (
            .O(N__7236),
            .I(N__7224));
    Span4Mux_v I__1764 (
            .O(N__7231),
            .I(N__7221));
    InMux I__1763 (
            .O(N__7230),
            .I(N__7218));
    Span12Mux_s9_h I__1762 (
            .O(N__7227),
            .I(N__7215));
    Span4Mux_v I__1761 (
            .O(N__7224),
            .I(N__7210));
    Span4Mux_h I__1760 (
            .O(N__7221),
            .I(N__7210));
    LocalMux I__1759 (
            .O(N__7218),
            .I(N__7207));
    Span12Mux_v I__1758 (
            .O(N__7215),
            .I(N__7204));
    Span4Mux_v I__1757 (
            .O(N__7210),
            .I(N__7201));
    Span4Mux_h I__1756 (
            .O(N__7207),
            .I(N__7198));
    Odrv12 I__1755 (
            .O(N__7204),
            .I(CPUBGn_c));
    Odrv4 I__1754 (
            .O(N__7201),
            .I(CPUBGn_c));
    Odrv4 I__1753 (
            .O(N__7198),
            .I(CPUBGn_c));
    InMux I__1752 (
            .O(N__7191),
            .I(N__7185));
    InMux I__1751 (
            .O(N__7190),
            .I(N__7178));
    InMux I__1750 (
            .O(N__7189),
            .I(N__7178));
    InMux I__1749 (
            .O(N__7188),
            .I(N__7178));
    LocalMux I__1748 (
            .O(N__7185),
            .I(N__7164));
    LocalMux I__1747 (
            .O(N__7178),
            .I(N__7161));
    InMux I__1746 (
            .O(N__7177),
            .I(N__7148));
    InMux I__1745 (
            .O(N__7176),
            .I(N__7148));
    InMux I__1744 (
            .O(N__7175),
            .I(N__7148));
    InMux I__1743 (
            .O(N__7174),
            .I(N__7148));
    InMux I__1742 (
            .O(N__7173),
            .I(N__7148));
    InMux I__1741 (
            .O(N__7172),
            .I(N__7148));
    InMux I__1740 (
            .O(N__7171),
            .I(N__7141));
    InMux I__1739 (
            .O(N__7170),
            .I(N__7141));
    InMux I__1738 (
            .O(N__7169),
            .I(N__7141));
    InMux I__1737 (
            .O(N__7168),
            .I(N__7134));
    InMux I__1736 (
            .O(N__7167),
            .I(N__7131));
    Span4Mux_v I__1735 (
            .O(N__7164),
            .I(N__7128));
    Span4Mux_h I__1734 (
            .O(N__7161),
            .I(N__7125));
    LocalMux I__1733 (
            .O(N__7148),
            .I(N__7122));
    LocalMux I__1732 (
            .O(N__7141),
            .I(N__7119));
    InMux I__1731 (
            .O(N__7140),
            .I(N__7112));
    InMux I__1730 (
            .O(N__7139),
            .I(N__7112));
    InMux I__1729 (
            .O(N__7138),
            .I(N__7112));
    InMux I__1728 (
            .O(N__7137),
            .I(N__7109));
    LocalMux I__1727 (
            .O(N__7134),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    LocalMux I__1726 (
            .O(N__7131),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    Odrv4 I__1725 (
            .O(N__7128),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    Odrv4 I__1724 (
            .O(N__7125),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    Odrv4 I__1723 (
            .O(N__7122),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    Odrv4 I__1722 (
            .O(N__7119),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    LocalMux I__1721 (
            .O(N__7112),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    LocalMux I__1720 (
            .O(N__7109),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ));
    CascadeMux I__1719 (
            .O(N__7092),
            .I(CPUBGn_c_cascade_));
    CascadeMux I__1718 (
            .O(N__7089),
            .I(N__7084));
    CascadeMux I__1717 (
            .O(N__7088),
            .I(N__7081));
    CascadeMux I__1716 (
            .O(N__7087),
            .I(N__7078));
    InMux I__1715 (
            .O(N__7084),
            .I(N__7075));
    InMux I__1714 (
            .O(N__7081),
            .I(N__7072));
    InMux I__1713 (
            .O(N__7078),
            .I(N__7069));
    LocalMux I__1712 (
            .O(N__7075),
            .I(N__7064));
    LocalMux I__1711 (
            .O(N__7072),
            .I(N__7059));
    LocalMux I__1710 (
            .O(N__7069),
            .I(N__7059));
    InMux I__1709 (
            .O(N__7068),
            .I(N__7056));
    InMux I__1708 (
            .O(N__7067),
            .I(N__7053));
    Span4Mux_v I__1707 (
            .O(N__7064),
            .I(N__7050));
    Span4Mux_h I__1706 (
            .O(N__7059),
            .I(N__7047));
    LocalMux I__1705 (
            .O(N__7056),
            .I(N__7044));
    LocalMux I__1704 (
            .O(N__7053),
            .I(N__7041));
    Span4Mux_v I__1703 (
            .O(N__7050),
            .I(N__7038));
    Span4Mux_v I__1702 (
            .O(N__7047),
            .I(N__7035));
    Sp12to4 I__1701 (
            .O(N__7044),
            .I(N__7032));
    Span12Mux_s11_v I__1700 (
            .O(N__7041),
            .I(N__7029));
    Sp12to4 I__1699 (
            .O(N__7038),
            .I(N__7022));
    Sp12to4 I__1698 (
            .O(N__7035),
            .I(N__7022));
    Span12Mux_v I__1697 (
            .O(N__7032),
            .I(N__7022));
    Span12Mux_h I__1696 (
            .O(N__7029),
            .I(N__7019));
    Span12Mux_h I__1695 (
            .O(N__7022),
            .I(N__7016));
    Odrv12 I__1694 (
            .O(N__7019),
            .I(RnW_c));
    Odrv12 I__1693 (
            .O(N__7016),
            .I(RnW_c));
    IoInMux I__1692 (
            .O(N__7011),
            .I(N__7006));
    IoInMux I__1691 (
            .O(N__7010),
            .I(N__7001));
    IoInMux I__1690 (
            .O(N__7009),
            .I(N__6998));
    LocalMux I__1689 (
            .O(N__7006),
            .I(N__6991));
    IoInMux I__1688 (
            .O(N__7005),
            .I(N__6988));
    IoInMux I__1687 (
            .O(N__7004),
            .I(N__6985));
    LocalMux I__1686 (
            .O(N__7001),
            .I(N__6980));
    LocalMux I__1685 (
            .O(N__6998),
            .I(N__6980));
    IoInMux I__1684 (
            .O(N__6997),
            .I(N__6977));
    IoInMux I__1683 (
            .O(N__6996),
            .I(N__6974));
    IoInMux I__1682 (
            .O(N__6995),
            .I(N__6966));
    IoInMux I__1681 (
            .O(N__6994),
            .I(N__6963));
    IoSpan4Mux I__1680 (
            .O(N__6991),
            .I(N__6953));
    LocalMux I__1679 (
            .O(N__6988),
            .I(N__6953));
    LocalMux I__1678 (
            .O(N__6985),
            .I(N__6953));
    Span4Mux_s2_h I__1677 (
            .O(N__6980),
            .I(N__6946));
    LocalMux I__1676 (
            .O(N__6977),
            .I(N__6946));
    LocalMux I__1675 (
            .O(N__6974),
            .I(N__6946));
    IoInMux I__1674 (
            .O(N__6973),
            .I(N__6943));
    IoInMux I__1673 (
            .O(N__6972),
            .I(N__6940));
    IoInMux I__1672 (
            .O(N__6971),
            .I(N__6937));
    IoInMux I__1671 (
            .O(N__6970),
            .I(N__6933));
    IoInMux I__1670 (
            .O(N__6969),
            .I(N__6928));
    LocalMux I__1669 (
            .O(N__6966),
            .I(N__6919));
    LocalMux I__1668 (
            .O(N__6963),
            .I(N__6919));
    IoInMux I__1667 (
            .O(N__6962),
            .I(N__6916));
    IoInMux I__1666 (
            .O(N__6961),
            .I(N__6913));
    IoInMux I__1665 (
            .O(N__6960),
            .I(N__6910));
    IoSpan4Mux I__1664 (
            .O(N__6953),
            .I(N__6897));
    IoSpan4Mux I__1663 (
            .O(N__6946),
            .I(N__6897));
    LocalMux I__1662 (
            .O(N__6943),
            .I(N__6897));
    LocalMux I__1661 (
            .O(N__6940),
            .I(N__6897));
    LocalMux I__1660 (
            .O(N__6937),
            .I(N__6897));
    IoInMux I__1659 (
            .O(N__6936),
            .I(N__6894));
    LocalMux I__1658 (
            .O(N__6933),
            .I(N__6891));
    IoInMux I__1657 (
            .O(N__6932),
            .I(N__6888));
    IoInMux I__1656 (
            .O(N__6931),
            .I(N__6885));
    LocalMux I__1655 (
            .O(N__6928),
            .I(N__6882));
    IoInMux I__1654 (
            .O(N__6927),
            .I(N__6879));
    IoInMux I__1653 (
            .O(N__6926),
            .I(N__6876));
    IoInMux I__1652 (
            .O(N__6925),
            .I(N__6873));
    IoInMux I__1651 (
            .O(N__6924),
            .I(N__6870));
    IoSpan4Mux I__1650 (
            .O(N__6919),
            .I(N__6861));
    LocalMux I__1649 (
            .O(N__6916),
            .I(N__6861));
    LocalMux I__1648 (
            .O(N__6913),
            .I(N__6861));
    LocalMux I__1647 (
            .O(N__6910),
            .I(N__6861));
    IoInMux I__1646 (
            .O(N__6909),
            .I(N__6856));
    IoInMux I__1645 (
            .O(N__6908),
            .I(N__6853));
    IoSpan4Mux I__1644 (
            .O(N__6897),
            .I(N__6844));
    LocalMux I__1643 (
            .O(N__6894),
            .I(N__6844));
    IoSpan4Mux I__1642 (
            .O(N__6891),
            .I(N__6837));
    LocalMux I__1641 (
            .O(N__6888),
            .I(N__6837));
    LocalMux I__1640 (
            .O(N__6885),
            .I(N__6837));
    IoSpan4Mux I__1639 (
            .O(N__6882),
            .I(N__6826));
    LocalMux I__1638 (
            .O(N__6879),
            .I(N__6826));
    LocalMux I__1637 (
            .O(N__6876),
            .I(N__6826));
    LocalMux I__1636 (
            .O(N__6873),
            .I(N__6826));
    LocalMux I__1635 (
            .O(N__6870),
            .I(N__6826));
    IoSpan4Mux I__1634 (
            .O(N__6861),
            .I(N__6823));
    IoInMux I__1633 (
            .O(N__6860),
            .I(N__6820));
    IoInMux I__1632 (
            .O(N__6859),
            .I(N__6817));
    LocalMux I__1631 (
            .O(N__6856),
            .I(N__6812));
    LocalMux I__1630 (
            .O(N__6853),
            .I(N__6812));
    IoInMux I__1629 (
            .O(N__6852),
            .I(N__6809));
    IoInMux I__1628 (
            .O(N__6851),
            .I(N__6806));
    IoInMux I__1627 (
            .O(N__6850),
            .I(N__6803));
    IoInMux I__1626 (
            .O(N__6849),
            .I(N__6800));
    Span4Mux_s2_v I__1625 (
            .O(N__6844),
            .I(N__6797));
    IoSpan4Mux I__1624 (
            .O(N__6837),
            .I(N__6792));
    IoSpan4Mux I__1623 (
            .O(N__6826),
            .I(N__6792));
    Span4Mux_s3_h I__1622 (
            .O(N__6823),
            .I(N__6789));
    LocalMux I__1621 (
            .O(N__6820),
            .I(N__6784));
    LocalMux I__1620 (
            .O(N__6817),
            .I(N__6784));
    Span12Mux_s5_h I__1619 (
            .O(N__6812),
            .I(N__6781));
    LocalMux I__1618 (
            .O(N__6809),
            .I(N__6778));
    LocalMux I__1617 (
            .O(N__6806),
            .I(N__6773));
    LocalMux I__1616 (
            .O(N__6803),
            .I(N__6773));
    LocalMux I__1615 (
            .O(N__6800),
            .I(N__6770));
    Span4Mux_h I__1614 (
            .O(N__6797),
            .I(N__6767));
    Span4Mux_s2_h I__1613 (
            .O(N__6792),
            .I(N__6764));
    Sp12to4 I__1612 (
            .O(N__6789),
            .I(N__6759));
    Span12Mux_s5_h I__1611 (
            .O(N__6784),
            .I(N__6759));
    Span12Mux_h I__1610 (
            .O(N__6781),
            .I(N__6756));
    Span12Mux_s6_v I__1609 (
            .O(N__6778),
            .I(N__6753));
    Span12Mux_s10_h I__1608 (
            .O(N__6773),
            .I(N__6750));
    Span12Mux_s10_h I__1607 (
            .O(N__6770),
            .I(N__6745));
    Sp12to4 I__1606 (
            .O(N__6767),
            .I(N__6745));
    Sp12to4 I__1605 (
            .O(N__6764),
            .I(N__6742));
    Span12Mux_h I__1604 (
            .O(N__6759),
            .I(N__6739));
    Span12Mux_v I__1603 (
            .O(N__6756),
            .I(N__6734));
    Span12Mux_h I__1602 (
            .O(N__6753),
            .I(N__6734));
    Span12Mux_v I__1601 (
            .O(N__6750),
            .I(N__6727));
    Span12Mux_v I__1600 (
            .O(N__6745),
            .I(N__6727));
    Span12Mux_s10_h I__1599 (
            .O(N__6742),
            .I(N__6727));
    Odrv12 I__1598 (
            .O(N__6739),
            .I(N_62_i));
    Odrv12 I__1597 (
            .O(N__6734),
            .I(N_62_i));
    Odrv12 I__1596 (
            .O(N__6727),
            .I(N_62_i));
    InMux I__1595 (
            .O(N__6720),
            .I(N__6717));
    LocalMux I__1594 (
            .O(N__6717),
            .I(N__6714));
    Span4Mux_v I__1593 (
            .O(N__6714),
            .I(N__6709));
    InMux I__1592 (
            .O(N__6713),
            .I(N__6706));
    CascadeMux I__1591 (
            .O(N__6712),
            .I(N__6703));
    Span4Mux_v I__1590 (
            .O(N__6709),
            .I(N__6700));
    LocalMux I__1589 (
            .O(N__6706),
            .I(N__6697));
    InMux I__1588 (
            .O(N__6703),
            .I(N__6694));
    Span4Mux_v I__1587 (
            .O(N__6700),
            .I(N__6689));
    Span4Mux_v I__1586 (
            .O(N__6697),
            .I(N__6689));
    LocalMux I__1585 (
            .O(N__6694),
            .I(N__6686));
    Sp12to4 I__1584 (
            .O(N__6689),
            .I(N__6681));
    Span12Mux_v I__1583 (
            .O(N__6686),
            .I(N__6681));
    Span12Mux_h I__1582 (
            .O(N__6681),
            .I(N__6678));
    Odrv12 I__1581 (
            .O(N__6678),
            .I(D_UM_AMIGA_in_2));
    InMux I__1580 (
            .O(N__6675),
            .I(N__6671));
    InMux I__1579 (
            .O(N__6674),
            .I(N__6668));
    LocalMux I__1578 (
            .O(N__6671),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ));
    LocalMux I__1577 (
            .O(N__6668),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ));
    IoInMux I__1576 (
            .O(N__6663),
            .I(N__6660));
    LocalMux I__1575 (
            .O(N__6660),
            .I(N__6657));
    IoSpan4Mux I__1574 (
            .O(N__6657),
            .I(N__6654));
    Span4Mux_s0_h I__1573 (
            .O(N__6654),
            .I(N__6651));
    Span4Mux_h I__1572 (
            .O(N__6651),
            .I(N__6648));
    Sp12to4 I__1571 (
            .O(N__6648),
            .I(N__6645));
    Odrv12 I__1570 (
            .O(N__6645),
            .I(un1_D_UM_AMIGA_2));
    InMux I__1569 (
            .O(N__6642),
            .I(N__6636));
    InMux I__1568 (
            .O(N__6641),
            .I(N__6636));
    LocalMux I__1567 (
            .O(N__6636),
            .I(N__6632));
    InMux I__1566 (
            .O(N__6635),
            .I(N__6629));
    Span4Mux_v I__1565 (
            .O(N__6632),
            .I(N__6621));
    LocalMux I__1564 (
            .O(N__6629),
            .I(N__6621));
    InMux I__1563 (
            .O(N__6628),
            .I(N__6618));
    InMux I__1562 (
            .O(N__6627),
            .I(N__6613));
    InMux I__1561 (
            .O(N__6626),
            .I(N__6613));
    Odrv4 I__1560 (
            .O(N__6621),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1559 (
            .O(N__6618),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    LocalMux I__1558 (
            .O(N__6613),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ));
    InMux I__1557 (
            .O(N__6606),
            .I(N__6597));
    InMux I__1556 (
            .O(N__6605),
            .I(N__6585));
    InMux I__1555 (
            .O(N__6604),
            .I(N__6580));
    InMux I__1554 (
            .O(N__6603),
            .I(N__6580));
    InMux I__1553 (
            .O(N__6602),
            .I(N__6577));
    InMux I__1552 (
            .O(N__6601),
            .I(N__6572));
    InMux I__1551 (
            .O(N__6600),
            .I(N__6572));
    LocalMux I__1550 (
            .O(N__6597),
            .I(N__6569));
    InMux I__1549 (
            .O(N__6596),
            .I(N__6556));
    InMux I__1548 (
            .O(N__6595),
            .I(N__6556));
    InMux I__1547 (
            .O(N__6594),
            .I(N__6556));
    InMux I__1546 (
            .O(N__6593),
            .I(N__6556));
    InMux I__1545 (
            .O(N__6592),
            .I(N__6556));
    InMux I__1544 (
            .O(N__6591),
            .I(N__6556));
    InMux I__1543 (
            .O(N__6590),
            .I(N__6549));
    InMux I__1542 (
            .O(N__6589),
            .I(N__6549));
    InMux I__1541 (
            .O(N__6588),
            .I(N__6549));
    LocalMux I__1540 (
            .O(N__6585),
            .I(\U111_CYCLE_SM.N_107_i ));
    LocalMux I__1539 (
            .O(N__6580),
            .I(\U111_CYCLE_SM.N_107_i ));
    LocalMux I__1538 (
            .O(N__6577),
            .I(\U111_CYCLE_SM.N_107_i ));
    LocalMux I__1537 (
            .O(N__6572),
            .I(\U111_CYCLE_SM.N_107_i ));
    Odrv4 I__1536 (
            .O(N__6569),
            .I(\U111_CYCLE_SM.N_107_i ));
    LocalMux I__1535 (
            .O(N__6556),
            .I(\U111_CYCLE_SM.N_107_i ));
    LocalMux I__1534 (
            .O(N__6549),
            .I(\U111_CYCLE_SM.N_107_i ));
    InMux I__1533 (
            .O(N__6534),
            .I(N__6530));
    InMux I__1532 (
            .O(N__6533),
            .I(N__6527));
    LocalMux I__1531 (
            .O(N__6530),
            .I(N__6524));
    LocalMux I__1530 (
            .O(N__6527),
            .I(N__6521));
    Span12Mux_h I__1529 (
            .O(N__6524),
            .I(N__6518));
    Sp12to4 I__1528 (
            .O(N__6521),
            .I(N__6515));
    Span12Mux_h I__1527 (
            .O(N__6518),
            .I(N__6512));
    Span12Mux_v I__1526 (
            .O(N__6515),
            .I(N__6509));
    Span12Mux_v I__1525 (
            .O(N__6512),
            .I(N__6506));
    Span12Mux_h I__1524 (
            .O(N__6509),
            .I(N__6503));
    Odrv12 I__1523 (
            .O(N__6506),
            .I(SIZ_c_1));
    Odrv12 I__1522 (
            .O(N__6503),
            .I(SIZ_c_1));
    InMux I__1521 (
            .O(N__6498),
            .I(N__6494));
    CascadeMux I__1520 (
            .O(N__6497),
            .I(N__6491));
    LocalMux I__1519 (
            .O(N__6494),
            .I(N__6488));
    InMux I__1518 (
            .O(N__6491),
            .I(N__6485));
    Span4Mux_h I__1517 (
            .O(N__6488),
            .I(N__6480));
    LocalMux I__1516 (
            .O(N__6485),
            .I(N__6480));
    Span4Mux_v I__1515 (
            .O(N__6480),
            .I(N__6477));
    Span4Mux_v I__1514 (
            .O(N__6477),
            .I(N__6474));
    Sp12to4 I__1513 (
            .O(N__6474),
            .I(N__6471));
    Span12Mux_h I__1512 (
            .O(N__6471),
            .I(N__6468));
    Odrv12 I__1511 (
            .O(N__6468),
            .I(SIZ_c_0));
    CascadeMux I__1510 (
            .O(N__6465),
            .I(N__6459));
    CascadeMux I__1509 (
            .O(N__6464),
            .I(N__6454));
    CascadeMux I__1508 (
            .O(N__6463),
            .I(N__6450));
    InMux I__1507 (
            .O(N__6462),
            .I(N__6447));
    InMux I__1506 (
            .O(N__6459),
            .I(N__6444));
    InMux I__1505 (
            .O(N__6458),
            .I(N__6441));
    InMux I__1504 (
            .O(N__6457),
            .I(N__6438));
    InMux I__1503 (
            .O(N__6454),
            .I(N__6433));
    InMux I__1502 (
            .O(N__6453),
            .I(N__6433));
    InMux I__1501 (
            .O(N__6450),
            .I(N__6430));
    LocalMux I__1500 (
            .O(N__6447),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    LocalMux I__1499 (
            .O(N__6444),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    LocalMux I__1498 (
            .O(N__6441),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    LocalMux I__1497 (
            .O(N__6438),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    LocalMux I__1496 (
            .O(N__6433),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    LocalMux I__1495 (
            .O(N__6430),
            .I(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ));
    InMux I__1494 (
            .O(N__6417),
            .I(N__6414));
    LocalMux I__1493 (
            .O(N__6414),
            .I(N__6410));
    InMux I__1492 (
            .O(N__6413),
            .I(N__6406));
    Span4Mux_h I__1491 (
            .O(N__6410),
            .I(N__6403));
    InMux I__1490 (
            .O(N__6409),
            .I(N__6400));
    LocalMux I__1489 (
            .O(N__6406),
            .I(N__6397));
    Odrv4 I__1488 (
            .O(N__6403),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    LocalMux I__1487 (
            .O(N__6400),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    Odrv4 I__1486 (
            .O(N__6397),
            .I(\U111_CYCLE_SM.LW_TRANSZ0 ));
    InMux I__1485 (
            .O(N__6390),
            .I(N__6387));
    LocalMux I__1484 (
            .O(N__6387),
            .I(N__6371));
    ClkMux I__1483 (
            .O(N__6386),
            .I(N__6342));
    ClkMux I__1482 (
            .O(N__6385),
            .I(N__6342));
    ClkMux I__1481 (
            .O(N__6384),
            .I(N__6342));
    ClkMux I__1480 (
            .O(N__6383),
            .I(N__6342));
    ClkMux I__1479 (
            .O(N__6382),
            .I(N__6342));
    ClkMux I__1478 (
            .O(N__6381),
            .I(N__6342));
    ClkMux I__1477 (
            .O(N__6380),
            .I(N__6342));
    ClkMux I__1476 (
            .O(N__6379),
            .I(N__6342));
    ClkMux I__1475 (
            .O(N__6378),
            .I(N__6342));
    ClkMux I__1474 (
            .O(N__6377),
            .I(N__6342));
    ClkMux I__1473 (
            .O(N__6376),
            .I(N__6342));
    ClkMux I__1472 (
            .O(N__6375),
            .I(N__6342));
    ClkMux I__1471 (
            .O(N__6374),
            .I(N__6342));
    Glb2LocalMux I__1470 (
            .O(N__6371),
            .I(N__6342));
    GlobalMux I__1469 (
            .O(N__6342),
            .I(CLK40));
    SRMux I__1468 (
            .O(N__6339),
            .I(N__6312));
    SRMux I__1467 (
            .O(N__6338),
            .I(N__6312));
    SRMux I__1466 (
            .O(N__6337),
            .I(N__6312));
    SRMux I__1465 (
            .O(N__6336),
            .I(N__6312));
    SRMux I__1464 (
            .O(N__6335),
            .I(N__6312));
    SRMux I__1463 (
            .O(N__6334),
            .I(N__6312));
    SRMux I__1462 (
            .O(N__6333),
            .I(N__6312));
    SRMux I__1461 (
            .O(N__6332),
            .I(N__6312));
    SRMux I__1460 (
            .O(N__6331),
            .I(N__6312));
    GlobalMux I__1459 (
            .O(N__6312),
            .I(N__6309));
    gio2CtrlBuf I__1458 (
            .O(N__6309),
            .I(RESETn_c_i_g));
    CascadeMux I__1457 (
            .O(N__6306),
            .I(N__6303));
    InMux I__1456 (
            .O(N__6303),
            .I(N__6300));
    LocalMux I__1455 (
            .O(N__6300),
            .I(N__6296));
    InMux I__1454 (
            .O(N__6299),
            .I(N__6293));
    Span4Mux_v I__1453 (
            .O(N__6296),
            .I(N__6289));
    LocalMux I__1452 (
            .O(N__6293),
            .I(N__6286));
    InMux I__1451 (
            .O(N__6292),
            .I(N__6283));
    Span4Mux_h I__1450 (
            .O(N__6289),
            .I(N__6278));
    Span4Mux_v I__1449 (
            .O(N__6286),
            .I(N__6278));
    LocalMux I__1448 (
            .O(N__6283),
            .I(N__6275));
    Span4Mux_v I__1447 (
            .O(N__6278),
            .I(N__6272));
    Span4Mux_v I__1446 (
            .O(N__6275),
            .I(N__6269));
    Span4Mux_v I__1445 (
            .O(N__6272),
            .I(N__6264));
    Span4Mux_h I__1444 (
            .O(N__6269),
            .I(N__6264));
    Sp12to4 I__1443 (
            .O(N__6264),
            .I(N__6261));
    Odrv12 I__1442 (
            .O(N__6261),
            .I(D_UU_AMIGA_in_1));
    InMux I__1441 (
            .O(N__6258),
            .I(N__6255));
    LocalMux I__1440 (
            .O(N__6255),
            .I(N__6251));
    InMux I__1439 (
            .O(N__6254),
            .I(N__6248));
    Odrv12 I__1438 (
            .O(N__6251),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ));
    LocalMux I__1437 (
            .O(N__6248),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ));
    IoInMux I__1436 (
            .O(N__6243),
            .I(N__6240));
    LocalMux I__1435 (
            .O(N__6240),
            .I(N__6237));
    IoSpan4Mux I__1434 (
            .O(N__6237),
            .I(N__6234));
    Span4Mux_s1_h I__1433 (
            .O(N__6234),
            .I(N__6231));
    Span4Mux_v I__1432 (
            .O(N__6231),
            .I(N__6228));
    Sp12to4 I__1431 (
            .O(N__6228),
            .I(N__6225));
    Span12Mux_s10_h I__1430 (
            .O(N__6225),
            .I(N__6222));
    Odrv12 I__1429 (
            .O(N__6222),
            .I(N_130));
    InMux I__1428 (
            .O(N__6219),
            .I(N__6216));
    LocalMux I__1427 (
            .O(N__6216),
            .I(N__6212));
    InMux I__1426 (
            .O(N__6215),
            .I(N__6209));
    Odrv12 I__1425 (
            .O(N__6212),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ));
    LocalMux I__1424 (
            .O(N__6209),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ));
    InMux I__1423 (
            .O(N__6204),
            .I(N__6201));
    LocalMux I__1422 (
            .O(N__6201),
            .I(N__6197));
    CascadeMux I__1421 (
            .O(N__6200),
            .I(N__6194));
    Span4Mux_v I__1420 (
            .O(N__6197),
            .I(N__6191));
    InMux I__1419 (
            .O(N__6194),
            .I(N__6188));
    Span4Mux_h I__1418 (
            .O(N__6191),
            .I(N__6183));
    LocalMux I__1417 (
            .O(N__6188),
            .I(N__6183));
    Span4Mux_v I__1416 (
            .O(N__6183),
            .I(N__6179));
    InMux I__1415 (
            .O(N__6182),
            .I(N__6176));
    Span4Mux_v I__1414 (
            .O(N__6179),
            .I(N__6171));
    LocalMux I__1413 (
            .O(N__6176),
            .I(N__6171));
    Span4Mux_v I__1412 (
            .O(N__6171),
            .I(N__6168));
    Sp12to4 I__1411 (
            .O(N__6168),
            .I(N__6165));
    Span12Mux_h I__1410 (
            .O(N__6165),
            .I(N__6162));
    Odrv12 I__1409 (
            .O(N__6162),
            .I(D_UU_AMIGA_in_0));
    IoInMux I__1408 (
            .O(N__6159),
            .I(N__6156));
    LocalMux I__1407 (
            .O(N__6156),
            .I(N__6153));
    Span4Mux_s3_v I__1406 (
            .O(N__6153),
            .I(N__6150));
    Span4Mux_v I__1405 (
            .O(N__6150),
            .I(N__6147));
    Sp12to4 I__1404 (
            .O(N__6147),
            .I(N__6144));
    Span12Mux_h I__1403 (
            .O(N__6144),
            .I(N__6141));
    Odrv12 I__1402 (
            .O(N__6141),
            .I(N_131));
    InMux I__1401 (
            .O(N__6138),
            .I(N__6134));
    InMux I__1400 (
            .O(N__6137),
            .I(N__6131));
    LocalMux I__1399 (
            .O(N__6134),
            .I(N__6127));
    LocalMux I__1398 (
            .O(N__6131),
            .I(N__6124));
    CascadeMux I__1397 (
            .O(N__6130),
            .I(N__6121));
    Span4Mux_v I__1396 (
            .O(N__6127),
            .I(N__6118));
    Span4Mux_v I__1395 (
            .O(N__6124),
            .I(N__6115));
    InMux I__1394 (
            .O(N__6121),
            .I(N__6112));
    Odrv4 I__1393 (
            .O(N__6118),
            .I(\U111_CYCLE_SM.TA_DISZ0 ));
    Odrv4 I__1392 (
            .O(N__6115),
            .I(\U111_CYCLE_SM.TA_DISZ0 ));
    LocalMux I__1391 (
            .O(N__6112),
            .I(\U111_CYCLE_SM.TA_DISZ0 ));
    IoInMux I__1390 (
            .O(N__6105),
            .I(N__6102));
    LocalMux I__1389 (
            .O(N__6102),
            .I(N__6099));
    IoSpan4Mux I__1388 (
            .O(N__6099),
            .I(N__6096));
    Span4Mux_s0_v I__1387 (
            .O(N__6096),
            .I(N__6093));
    Span4Mux_v I__1386 (
            .O(N__6093),
            .I(N__6090));
    Span4Mux_v I__1385 (
            .O(N__6090),
            .I(N__6087));
    Odrv4 I__1384 (
            .O(N__6087),
            .I(N_66));
    CascadeMux I__1383 (
            .O(N__6084),
            .I(N__6081));
    InMux I__1382 (
            .O(N__6081),
            .I(N__6077));
    InMux I__1381 (
            .O(N__6080),
            .I(N__6074));
    LocalMux I__1380 (
            .O(N__6077),
            .I(N__6071));
    LocalMux I__1379 (
            .O(N__6074),
            .I(N__6067));
    Span4Mux_v I__1378 (
            .O(N__6071),
            .I(N__6064));
    InMux I__1377 (
            .O(N__6070),
            .I(N__6061));
    Span4Mux_h I__1376 (
            .O(N__6067),
            .I(N__6058));
    Span4Mux_v I__1375 (
            .O(N__6064),
            .I(N__6053));
    LocalMux I__1374 (
            .O(N__6061),
            .I(N__6053));
    Span4Mux_v I__1373 (
            .O(N__6058),
            .I(N__6050));
    Span4Mux_v I__1372 (
            .O(N__6053),
            .I(N__6047));
    Sp12to4 I__1371 (
            .O(N__6050),
            .I(N__6044));
    Span4Mux_h I__1370 (
            .O(N__6047),
            .I(N__6041));
    Span12Mux_v I__1369 (
            .O(N__6044),
            .I(N__6036));
    Sp12to4 I__1368 (
            .O(N__6041),
            .I(N__6036));
    Odrv12 I__1367 (
            .O(N__6036),
            .I(D_UM_AMIGA_in_3));
    InMux I__1366 (
            .O(N__6033),
            .I(N__6030));
    LocalMux I__1365 (
            .O(N__6030),
            .I(N__6027));
    Span4Mux_v I__1364 (
            .O(N__6027),
            .I(N__6023));
    InMux I__1363 (
            .O(N__6026),
            .I(N__6020));
    Odrv4 I__1362 (
            .O(N__6023),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ));
    LocalMux I__1361 (
            .O(N__6020),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ));
    IoInMux I__1360 (
            .O(N__6015),
            .I(N__6012));
    LocalMux I__1359 (
            .O(N__6012),
            .I(N__6009));
    Span12Mux_s7_h I__1358 (
            .O(N__6009),
            .I(N__6006));
    Span12Mux_h I__1357 (
            .O(N__6006),
            .I(N__6003));
    Odrv12 I__1356 (
            .O(N__6003),
            .I(un1_D_UM_AMIGA_3));
    InMux I__1355 (
            .O(N__6000),
            .I(N__5996));
    IoInMux I__1354 (
            .O(N__5999),
            .I(N__5993));
    LocalMux I__1353 (
            .O(N__5996),
            .I(N__5990));
    LocalMux I__1352 (
            .O(N__5993),
            .I(N__5987));
    Span4Mux_v I__1351 (
            .O(N__5990),
            .I(N__5984));
    Span4Mux_s2_h I__1350 (
            .O(N__5987),
            .I(N__5981));
    Sp12to4 I__1349 (
            .O(N__5984),
            .I(N__5978));
    Span4Mux_v I__1348 (
            .O(N__5981),
            .I(N__5975));
    Span12Mux_v I__1347 (
            .O(N__5978),
            .I(N__5972));
    Sp12to4 I__1346 (
            .O(N__5975),
            .I(N__5969));
    Span12Mux_v I__1345 (
            .O(N__5972),
            .I(N__5964));
    Span12Mux_h I__1344 (
            .O(N__5969),
            .I(N__5964));
    Span12Mux_h I__1343 (
            .O(N__5964),
            .I(N__5961));
    Odrv12 I__1342 (
            .O(N__5961),
            .I(D_LL_040_in_4));
    InMux I__1341 (
            .O(N__5958),
            .I(N__5955));
    LocalMux I__1340 (
            .O(N__5955),
            .I(N__5952));
    Span4Mux_v I__1339 (
            .O(N__5952),
            .I(N__5949));
    Span4Mux_h I__1338 (
            .O(N__5949),
            .I(N__5946));
    Sp12to4 I__1337 (
            .O(N__5946),
            .I(N__5943));
    Span12Mux_h I__1336 (
            .O(N__5943),
            .I(N__5940));
    Odrv12 I__1335 (
            .O(N__5940),
            .I(D_UM_040_in_4));
    IoInMux I__1334 (
            .O(N__5937),
            .I(N__5934));
    LocalMux I__1333 (
            .O(N__5934),
            .I(N__5931));
    IoSpan4Mux I__1332 (
            .O(N__5931),
            .I(N__5928));
    Sp12to4 I__1331 (
            .O(N__5928),
            .I(N__5925));
    Span12Mux_h I__1330 (
            .O(N__5925),
            .I(N__5922));
    Odrv12 I__1329 (
            .O(N__5922),
            .I(un1_D_UM_040_4));
    InMux I__1328 (
            .O(N__5919),
            .I(N__5916));
    LocalMux I__1327 (
            .O(N__5916),
            .I(N__5913));
    Span4Mux_v I__1326 (
            .O(N__5913),
            .I(N__5910));
    Sp12to4 I__1325 (
            .O(N__5910),
            .I(N__5907));
    Span12Mux_h I__1324 (
            .O(N__5907),
            .I(N__5904));
    Odrv12 I__1323 (
            .O(N__5904),
            .I(D_LL_AMIGA_in_6));
    IoInMux I__1322 (
            .O(N__5901),
            .I(N__5898));
    LocalMux I__1321 (
            .O(N__5898),
            .I(N__5895));
    Span4Mux_s2_h I__1320 (
            .O(N__5895),
            .I(N__5892));
    Span4Mux_h I__1319 (
            .O(N__5892),
            .I(N__5889));
    Sp12to4 I__1318 (
            .O(N__5889),
            .I(N__5886));
    Span12Mux_s10_v I__1317 (
            .O(N__5886),
            .I(N__5883));
    Span12Mux_h I__1316 (
            .O(N__5883),
            .I(N__5880));
    Odrv12 I__1315 (
            .O(N__5880),
            .I(un2_D_LL_AMIGA_6));
    InMux I__1314 (
            .O(N__5877),
            .I(N__5874));
    LocalMux I__1313 (
            .O(N__5874),
            .I(N__5871));
    Span12Mux_v I__1312 (
            .O(N__5871),
            .I(N__5868));
    Span12Mux_h I__1311 (
            .O(N__5868),
            .I(N__5865));
    Odrv12 I__1310 (
            .O(N__5865),
            .I(D_LL_AMIGA_in_5));
    IoInMux I__1309 (
            .O(N__5862),
            .I(N__5859));
    LocalMux I__1308 (
            .O(N__5859),
            .I(N__5856));
    Span4Mux_s3_h I__1307 (
            .O(N__5856),
            .I(N__5853));
    Span4Mux_v I__1306 (
            .O(N__5853),
            .I(N__5850));
    Span4Mux_v I__1305 (
            .O(N__5850),
            .I(N__5847));
    Span4Mux_h I__1304 (
            .O(N__5847),
            .I(N__5844));
    Sp12to4 I__1303 (
            .O(N__5844),
            .I(N__5841));
    Odrv12 I__1302 (
            .O(N__5841),
            .I(un2_D_LL_AMIGA_5));
    InMux I__1301 (
            .O(N__5838),
            .I(N__5835));
    LocalMux I__1300 (
            .O(N__5835),
            .I(N__5832));
    Span4Mux_v I__1299 (
            .O(N__5832),
            .I(N__5829));
    Span4Mux_h I__1298 (
            .O(N__5829),
            .I(N__5826));
    Sp12to4 I__1297 (
            .O(N__5826),
            .I(N__5823));
    Span12Mux_v I__1296 (
            .O(N__5823),
            .I(N__5820));
    Odrv12 I__1295 (
            .O(N__5820),
            .I(TS_CPUn_in));
    CascadeMux I__1294 (
            .O(N__5817),
            .I(N__5813));
    InMux I__1293 (
            .O(N__5816),
            .I(N__5810));
    InMux I__1292 (
            .O(N__5813),
            .I(N__5807));
    LocalMux I__1291 (
            .O(N__5810),
            .I(\U111_CYCLE_SM.TS_DELAYZ0 ));
    LocalMux I__1290 (
            .O(N__5807),
            .I(\U111_CYCLE_SM.TS_DELAYZ0 ));
    InMux I__1289 (
            .O(N__5802),
            .I(N__5797));
    InMux I__1288 (
            .O(N__5801),
            .I(N__5794));
    InMux I__1287 (
            .O(N__5800),
            .I(N__5791));
    LocalMux I__1286 (
            .O(N__5797),
            .I(\U111_CYCLE_SM.un4_TS_OUT_i_0 ));
    LocalMux I__1285 (
            .O(N__5794),
            .I(\U111_CYCLE_SM.un4_TS_OUT_i_0 ));
    LocalMux I__1284 (
            .O(N__5791),
            .I(\U111_CYCLE_SM.un4_TS_OUT_i_0 ));
    InMux I__1283 (
            .O(N__5784),
            .I(N__5780));
    InMux I__1282 (
            .O(N__5783),
            .I(N__5777));
    LocalMux I__1281 (
            .O(N__5780),
            .I(\U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0 ));
    LocalMux I__1280 (
            .O(N__5777),
            .I(\U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0 ));
    IoInMux I__1279 (
            .O(N__5772),
            .I(N__5769));
    LocalMux I__1278 (
            .O(N__5769),
            .I(N__5765));
    IoInMux I__1277 (
            .O(N__5768),
            .I(N__5761));
    IoSpan4Mux I__1276 (
            .O(N__5765),
            .I(N__5758));
    IoInMux I__1275 (
            .O(N__5764),
            .I(N__5755));
    LocalMux I__1274 (
            .O(N__5761),
            .I(N__5751));
    IoSpan4Mux I__1273 (
            .O(N__5758),
            .I(N__5746));
    LocalMux I__1272 (
            .O(N__5755),
            .I(N__5746));
    IoInMux I__1271 (
            .O(N__5754),
            .I(N__5743));
    IoSpan4Mux I__1270 (
            .O(N__5751),
            .I(N__5740));
    IoSpan4Mux I__1269 (
            .O(N__5746),
            .I(N__5737));
    LocalMux I__1268 (
            .O(N__5743),
            .I(N__5734));
    Sp12to4 I__1267 (
            .O(N__5740),
            .I(N__5731));
    Span4Mux_s0_v I__1266 (
            .O(N__5737),
            .I(N__5728));
    Span4Mux_s1_h I__1265 (
            .O(N__5734),
            .I(N__5725));
    Span12Mux_s7_h I__1264 (
            .O(N__5731),
            .I(N__5722));
    Sp12to4 I__1263 (
            .O(N__5728),
            .I(N__5719));
    Sp12to4 I__1262 (
            .O(N__5725),
            .I(N__5716));
    Span12Mux_h I__1261 (
            .O(N__5722),
            .I(N__5711));
    Span12Mux_v I__1260 (
            .O(N__5719),
            .I(N__5711));
    Span12Mux_v I__1259 (
            .O(N__5716),
            .I(N__5708));
    Odrv12 I__1258 (
            .O(N__5711),
            .I(GB_BUFFER_CLK40_THRU_CO));
    Odrv12 I__1257 (
            .O(N__5708),
            .I(GB_BUFFER_CLK40_THRU_CO));
    InMux I__1256 (
            .O(N__5703),
            .I(N__5700));
    LocalMux I__1255 (
            .O(N__5700),
            .I(N__5696));
    InMux I__1254 (
            .O(N__5699),
            .I(N__5693));
    Odrv12 I__1253 (
            .O(N__5696),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ));
    LocalMux I__1252 (
            .O(N__5693),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ));
    CascadeMux I__1251 (
            .O(N__5688),
            .I(N__5685));
    InMux I__1250 (
            .O(N__5685),
            .I(N__5682));
    LocalMux I__1249 (
            .O(N__5682),
            .I(N__5678));
    InMux I__1248 (
            .O(N__5681),
            .I(N__5675));
    Span4Mux_v I__1247 (
            .O(N__5678),
            .I(N__5672));
    LocalMux I__1246 (
            .O(N__5675),
            .I(N__5669));
    Span4Mux_v I__1245 (
            .O(N__5672),
            .I(N__5663));
    Span4Mux_v I__1244 (
            .O(N__5669),
            .I(N__5663));
    InMux I__1243 (
            .O(N__5668),
            .I(N__5660));
    Sp12to4 I__1242 (
            .O(N__5663),
            .I(N__5655));
    LocalMux I__1241 (
            .O(N__5660),
            .I(N__5655));
    Span12Mux_h I__1240 (
            .O(N__5655),
            .I(N__5652));
    Odrv12 I__1239 (
            .O(N__5652),
            .I(D_UU_AMIGA_in_6));
    IoInMux I__1238 (
            .O(N__5649),
            .I(N__5646));
    LocalMux I__1237 (
            .O(N__5646),
            .I(N__5643));
    Span4Mux_s3_v I__1236 (
            .O(N__5643),
            .I(N__5640));
    Span4Mux_h I__1235 (
            .O(N__5640),
            .I(N__5637));
    Sp12to4 I__1234 (
            .O(N__5637),
            .I(N__5634));
    Span12Mux_s11_v I__1233 (
            .O(N__5634),
            .I(N__5631));
    Span12Mux_h I__1232 (
            .O(N__5631),
            .I(N__5628));
    Odrv12 I__1231 (
            .O(N__5628),
            .I(N_124));
    CascadeMux I__1230 (
            .O(N__5625),
            .I(N__5622));
    InMux I__1229 (
            .O(N__5622),
            .I(N__5619));
    LocalMux I__1228 (
            .O(N__5619),
            .I(N__5615));
    InMux I__1227 (
            .O(N__5618),
            .I(N__5612));
    Span4Mux_v I__1226 (
            .O(N__5615),
            .I(N__5606));
    LocalMux I__1225 (
            .O(N__5612),
            .I(N__5606));
    InMux I__1224 (
            .O(N__5611),
            .I(N__5603));
    Span4Mux_v I__1223 (
            .O(N__5606),
            .I(N__5600));
    LocalMux I__1222 (
            .O(N__5603),
            .I(N__5597));
    Span4Mux_v I__1221 (
            .O(N__5600),
            .I(N__5592));
    Span4Mux_v I__1220 (
            .O(N__5597),
            .I(N__5592));
    Span4Mux_v I__1219 (
            .O(N__5592),
            .I(N__5589));
    Span4Mux_h I__1218 (
            .O(N__5589),
            .I(N__5586));
    Sp12to4 I__1217 (
            .O(N__5586),
            .I(N__5583));
    Odrv12 I__1216 (
            .O(N__5583),
            .I(D_UU_AMIGA_in_5));
    InMux I__1215 (
            .O(N__5580),
            .I(N__5577));
    LocalMux I__1214 (
            .O(N__5577),
            .I(N__5573));
    InMux I__1213 (
            .O(N__5576),
            .I(N__5570));
    Odrv12 I__1212 (
            .O(N__5573),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ));
    LocalMux I__1211 (
            .O(N__5570),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ));
    IoInMux I__1210 (
            .O(N__5565),
            .I(N__5562));
    LocalMux I__1209 (
            .O(N__5562),
            .I(N__5559));
    Span4Mux_s1_v I__1208 (
            .O(N__5559),
            .I(N__5556));
    Span4Mux_h I__1207 (
            .O(N__5556),
            .I(N__5553));
    Span4Mux_v I__1206 (
            .O(N__5553),
            .I(N__5550));
    Span4Mux_v I__1205 (
            .O(N__5550),
            .I(N__5547));
    Sp12to4 I__1204 (
            .O(N__5547),
            .I(N__5544));
    Odrv12 I__1203 (
            .O(N__5544),
            .I(N_126));
    InMux I__1202 (
            .O(N__5541),
            .I(N__5537));
    InMux I__1201 (
            .O(N__5540),
            .I(N__5534));
    LocalMux I__1200 (
            .O(N__5537),
            .I(N__5531));
    LocalMux I__1199 (
            .O(N__5534),
            .I(N__5528));
    Span4Mux_v I__1198 (
            .O(N__5531),
            .I(N__5522));
    Span4Mux_v I__1197 (
            .O(N__5528),
            .I(N__5522));
    InMux I__1196 (
            .O(N__5527),
            .I(N__5519));
    Sp12to4 I__1195 (
            .O(N__5522),
            .I(N__5514));
    LocalMux I__1194 (
            .O(N__5519),
            .I(N__5514));
    Span12Mux_h I__1193 (
            .O(N__5514),
            .I(N__5511));
    Odrv12 I__1192 (
            .O(N__5511),
            .I(D_UU_AMIGA_in_7));
    InMux I__1191 (
            .O(N__5508),
            .I(N__5504));
    CascadeMux I__1190 (
            .O(N__5507),
            .I(N__5501));
    LocalMux I__1189 (
            .O(N__5504),
            .I(N__5498));
    InMux I__1188 (
            .O(N__5501),
            .I(N__5495));
    Odrv12 I__1187 (
            .O(N__5498),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ));
    LocalMux I__1186 (
            .O(N__5495),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ));
    IoInMux I__1185 (
            .O(N__5490),
            .I(N__5487));
    LocalMux I__1184 (
            .O(N__5487),
            .I(N__5484));
    IoSpan4Mux I__1183 (
            .O(N__5484),
            .I(N__5481));
    IoSpan4Mux I__1182 (
            .O(N__5481),
            .I(N__5478));
    Span4Mux_s1_v I__1181 (
            .O(N__5478),
            .I(N__5475));
    Sp12to4 I__1180 (
            .O(N__5475),
            .I(N__5472));
    Span12Mux_s9_v I__1179 (
            .O(N__5472),
            .I(N__5469));
    Odrv12 I__1178 (
            .O(N__5469),
            .I(N_123));
    InMux I__1177 (
            .O(N__5466),
            .I(N__5463));
    LocalMux I__1176 (
            .O(N__5463),
            .I(N__5459));
    InMux I__1175 (
            .O(N__5462),
            .I(N__5456));
    Odrv12 I__1174 (
            .O(N__5459),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ));
    LocalMux I__1173 (
            .O(N__5456),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ));
    CascadeMux I__1172 (
            .O(N__5451),
            .I(N__5448));
    InMux I__1171 (
            .O(N__5448),
            .I(N__5445));
    LocalMux I__1170 (
            .O(N__5445),
            .I(N__5441));
    InMux I__1169 (
            .O(N__5444),
            .I(N__5437));
    Span4Mux_v I__1168 (
            .O(N__5441),
            .I(N__5434));
    InMux I__1167 (
            .O(N__5440),
            .I(N__5431));
    LocalMux I__1166 (
            .O(N__5437),
            .I(N__5428));
    Span4Mux_h I__1165 (
            .O(N__5434),
            .I(N__5423));
    LocalMux I__1164 (
            .O(N__5431),
            .I(N__5423));
    Span4Mux_v I__1163 (
            .O(N__5428),
            .I(N__5420));
    Span4Mux_v I__1162 (
            .O(N__5423),
            .I(N__5417));
    Sp12to4 I__1161 (
            .O(N__5420),
            .I(N__5412));
    Sp12to4 I__1160 (
            .O(N__5417),
            .I(N__5412));
    Span12Mux_h I__1159 (
            .O(N__5412),
            .I(N__5409));
    Odrv12 I__1158 (
            .O(N__5409),
            .I(D_UU_AMIGA_in_4));
    IoInMux I__1157 (
            .O(N__5406),
            .I(N__5403));
    LocalMux I__1156 (
            .O(N__5403),
            .I(N__5400));
    Span4Mux_s0_v I__1155 (
            .O(N__5400),
            .I(N__5397));
    Sp12to4 I__1154 (
            .O(N__5397),
            .I(N__5394));
    Span12Mux_h I__1153 (
            .O(N__5394),
            .I(N__5391));
    Odrv12 I__1152 (
            .O(N__5391),
            .I(N_127));
    InMux I__1151 (
            .O(N__5388),
            .I(N__5385));
    LocalMux I__1150 (
            .O(N__5385),
            .I(N__5377));
    InMux I__1149 (
            .O(N__5384),
            .I(N__5370));
    InMux I__1148 (
            .O(N__5383),
            .I(N__5370));
    InMux I__1147 (
            .O(N__5382),
            .I(N__5370));
    InMux I__1146 (
            .O(N__5381),
            .I(N__5367));
    InMux I__1145 (
            .O(N__5380),
            .I(N__5364));
    Span4Mux_v I__1144 (
            .O(N__5377),
            .I(N__5361));
    LocalMux I__1143 (
            .O(N__5370),
            .I(N__5358));
    LocalMux I__1142 (
            .O(N__5367),
            .I(N__5355));
    LocalMux I__1141 (
            .O(N__5364),
            .I(N__5352));
    Sp12to4 I__1140 (
            .O(N__5361),
            .I(N__5347));
    Span4Mux_h I__1139 (
            .O(N__5358),
            .I(N__5344));
    Span4Mux_v I__1138 (
            .O(N__5355),
            .I(N__5339));
    Span4Mux_v I__1137 (
            .O(N__5352),
            .I(N__5339));
    InMux I__1136 (
            .O(N__5351),
            .I(N__5334));
    InMux I__1135 (
            .O(N__5350),
            .I(N__5334));
    Span12Mux_h I__1134 (
            .O(N__5347),
            .I(N__5331));
    Span4Mux_v I__1133 (
            .O(N__5344),
            .I(N__5328));
    Sp12to4 I__1132 (
            .O(N__5339),
            .I(N__5323));
    LocalMux I__1131 (
            .O(N__5334),
            .I(N__5323));
    Span12Mux_v I__1130 (
            .O(N__5331),
            .I(N__5316));
    Sp12to4 I__1129 (
            .O(N__5328),
            .I(N__5316));
    Span12Mux_h I__1128 (
            .O(N__5323),
            .I(N__5316));
    Span12Mux_v I__1127 (
            .O(N__5316),
            .I(N__5313));
    Odrv12 I__1126 (
            .O(N__5313),
            .I(TEAn_c));
    IoInMux I__1125 (
            .O(N__5310),
            .I(N__5307));
    LocalMux I__1124 (
            .O(N__5307),
            .I(N__5304));
    Span12Mux_s8_v I__1123 (
            .O(N__5304),
            .I(N__5301));
    Odrv12 I__1122 (
            .O(N__5301),
            .I(U111_CYCLE_SM_TEA_CPUn_0_i));
    InMux I__1121 (
            .O(N__5298),
            .I(N__5295));
    LocalMux I__1120 (
            .O(N__5295),
            .I(N__5292));
    Span4Mux_v I__1119 (
            .O(N__5292),
            .I(N__5289));
    Span4Mux_v I__1118 (
            .O(N__5289),
            .I(N__5286));
    Sp12to4 I__1117 (
            .O(N__5286),
            .I(N__5283));
    Span12Mux_h I__1116 (
            .O(N__5283),
            .I(N__5280));
    Odrv12 I__1115 (
            .O(N__5280),
            .I(D_UU_040_in_1));
    IoInMux I__1114 (
            .O(N__5277),
            .I(N__5273));
    InMux I__1113 (
            .O(N__5276),
            .I(N__5270));
    LocalMux I__1112 (
            .O(N__5273),
            .I(N__5267));
    LocalMux I__1111 (
            .O(N__5270),
            .I(N__5264));
    Span4Mux_s3_h I__1110 (
            .O(N__5267),
            .I(N__5261));
    Span4Mux_h I__1109 (
            .O(N__5264),
            .I(N__5258));
    Sp12to4 I__1108 (
            .O(N__5261),
            .I(N__5255));
    Sp12to4 I__1107 (
            .O(N__5258),
            .I(N__5252));
    Span12Mux_v I__1106 (
            .O(N__5255),
            .I(N__5249));
    Span12Mux_v I__1105 (
            .O(N__5252),
            .I(N__5246));
    Span12Mux_h I__1104 (
            .O(N__5249),
            .I(N__5241));
    Span12Mux_v I__1103 (
            .O(N__5246),
            .I(N__5241));
    Span12Mux_h I__1102 (
            .O(N__5241),
            .I(N__5238));
    Odrv12 I__1101 (
            .O(N__5238),
            .I(D_LM_040_in_1));
    IoInMux I__1100 (
            .O(N__5235),
            .I(N__5232));
    LocalMux I__1099 (
            .O(N__5232),
            .I(N__5229));
    Span12Mux_s0_h I__1098 (
            .O(N__5229),
            .I(N__5226));
    Span12Mux_h I__1097 (
            .O(N__5226),
            .I(N__5223));
    Odrv12 I__1096 (
            .O(N__5223),
            .I(un1_D_UU_040_1));
    InMux I__1095 (
            .O(N__5220),
            .I(N__5217));
    LocalMux I__1094 (
            .O(N__5217),
            .I(N__5214));
    Span4Mux_v I__1093 (
            .O(N__5214),
            .I(N__5211));
    Span4Mux_v I__1092 (
            .O(N__5211),
            .I(N__5208));
    Sp12to4 I__1091 (
            .O(N__5208),
            .I(N__5205));
    Span12Mux_h I__1090 (
            .O(N__5205),
            .I(N__5202));
    Odrv12 I__1089 (
            .O(N__5202),
            .I(D_UM_040_in_7));
    IoInMux I__1088 (
            .O(N__5199),
            .I(N__5195));
    InMux I__1087 (
            .O(N__5198),
            .I(N__5192));
    LocalMux I__1086 (
            .O(N__5195),
            .I(N__5189));
    LocalMux I__1085 (
            .O(N__5192),
            .I(N__5186));
    IoSpan4Mux I__1084 (
            .O(N__5189),
            .I(N__5183));
    Span4Mux_h I__1083 (
            .O(N__5186),
            .I(N__5180));
    Span4Mux_s3_h I__1082 (
            .O(N__5183),
            .I(N__5177));
    Sp12to4 I__1081 (
            .O(N__5180),
            .I(N__5174));
    Sp12to4 I__1080 (
            .O(N__5177),
            .I(N__5171));
    Span12Mux_v I__1079 (
            .O(N__5174),
            .I(N__5168));
    Span12Mux_v I__1078 (
            .O(N__5171),
            .I(N__5165));
    Span12Mux_h I__1077 (
            .O(N__5168),
            .I(N__5162));
    Span12Mux_h I__1076 (
            .O(N__5165),
            .I(N__5159));
    Span12Mux_v I__1075 (
            .O(N__5162),
            .I(N__5154));
    Span12Mux_h I__1074 (
            .O(N__5159),
            .I(N__5154));
    Odrv12 I__1073 (
            .O(N__5154),
            .I(D_LL_040_in_7));
    IoInMux I__1072 (
            .O(N__5151),
            .I(N__5148));
    LocalMux I__1071 (
            .O(N__5148),
            .I(N__5145));
    IoSpan4Mux I__1070 (
            .O(N__5145),
            .I(N__5142));
    Sp12to4 I__1069 (
            .O(N__5142),
            .I(N__5139));
    Span12Mux_s6_h I__1068 (
            .O(N__5139),
            .I(N__5136));
    Odrv12 I__1067 (
            .O(N__5136),
            .I(un1_D_UM_040_7));
    InMux I__1066 (
            .O(N__5133),
            .I(N__5130));
    LocalMux I__1065 (
            .O(N__5130),
            .I(N__5127));
    Odrv4 I__1064 (
            .O(N__5127),
            .I(\U111_CYCLE_SM.LATCH_EN_5 ));
    InMux I__1063 (
            .O(N__5124),
            .I(N__5116));
    InMux I__1062 (
            .O(N__5123),
            .I(N__5116));
    InMux I__1061 (
            .O(N__5122),
            .I(N__5109));
    InMux I__1060 (
            .O(N__5121),
            .I(N__5109));
    LocalMux I__1059 (
            .O(N__5116),
            .I(N__5106));
    InMux I__1058 (
            .O(N__5115),
            .I(N__5101));
    InMux I__1057 (
            .O(N__5114),
            .I(N__5101));
    LocalMux I__1056 (
            .O(N__5109),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    Odrv4 I__1055 (
            .O(N__5106),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    LocalMux I__1054 (
            .O(N__5101),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ));
    InMux I__1053 (
            .O(N__5094),
            .I(N__5090));
    InMux I__1052 (
            .O(N__5093),
            .I(N__5083));
    LocalMux I__1051 (
            .O(N__5090),
            .I(N__5080));
    InMux I__1050 (
            .O(N__5089),
            .I(N__5075));
    InMux I__1049 (
            .O(N__5088),
            .I(N__5075));
    InMux I__1048 (
            .O(N__5087),
            .I(N__5072));
    InMux I__1047 (
            .O(N__5086),
            .I(N__5069));
    LocalMux I__1046 (
            .O(N__5083),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    Odrv4 I__1045 (
            .O(N__5080),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1044 (
            .O(N__5075),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1043 (
            .O(N__5072),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    LocalMux I__1042 (
            .O(N__5069),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ));
    InMux I__1041 (
            .O(N__5058),
            .I(N__5055));
    LocalMux I__1040 (
            .O(N__5055),
            .I(N__5052));
    Odrv4 I__1039 (
            .O(N__5052),
            .I(\U111_CYCLE_SM.N_57 ));
    InMux I__1038 (
            .O(N__5049),
            .I(N__5046));
    LocalMux I__1037 (
            .O(N__5046),
            .I(N__5041));
    InMux I__1036 (
            .O(N__5045),
            .I(N__5038));
    InMux I__1035 (
            .O(N__5044),
            .I(N__5035));
    Span4Mux_v I__1034 (
            .O(N__5041),
            .I(N__5028));
    LocalMux I__1033 (
            .O(N__5038),
            .I(N__5028));
    LocalMux I__1032 (
            .O(N__5035),
            .I(N__5028));
    Span4Mux_v I__1031 (
            .O(N__5028),
            .I(N__5025));
    Span4Mux_v I__1030 (
            .O(N__5025),
            .I(N__5022));
    Span4Mux_v I__1029 (
            .O(N__5022),
            .I(N__5019));
    Sp12to4 I__1028 (
            .O(N__5019),
            .I(N__5016));
    Odrv12 I__1027 (
            .O(N__5016),
            .I(D_UM_AMIGA_in_7));
    CascadeMux I__1026 (
            .O(N__5013),
            .I(N__5009));
    InMux I__1025 (
            .O(N__5012),
            .I(N__5006));
    InMux I__1024 (
            .O(N__5009),
            .I(N__5003));
    LocalMux I__1023 (
            .O(N__5006),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ));
    LocalMux I__1022 (
            .O(N__5003),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ));
    IoInMux I__1021 (
            .O(N__4998),
            .I(N__4995));
    LocalMux I__1020 (
            .O(N__4995),
            .I(N__4992));
    Span4Mux_s0_h I__1019 (
            .O(N__4992),
            .I(N__4989));
    Sp12to4 I__1018 (
            .O(N__4989),
            .I(N__4986));
    Span12Mux_v I__1017 (
            .O(N__4986),
            .I(N__4983));
    Span12Mux_h I__1016 (
            .O(N__4983),
            .I(N__4980));
    Odrv12 I__1015 (
            .O(N__4980),
            .I(un1_D_UM_AMIGA_7));
    CascadeMux I__1014 (
            .O(N__4977),
            .I(N__4974));
    InMux I__1013 (
            .O(N__4974),
            .I(N__4970));
    InMux I__1012 (
            .O(N__4973),
            .I(N__4967));
    LocalMux I__1011 (
            .O(N__4970),
            .I(N__4964));
    LocalMux I__1010 (
            .O(N__4967),
            .I(N__4961));
    Span4Mux_v I__1009 (
            .O(N__4964),
            .I(N__4957));
    Span4Mux_v I__1008 (
            .O(N__4961),
            .I(N__4954));
    InMux I__1007 (
            .O(N__4960),
            .I(N__4951));
    Span4Mux_h I__1006 (
            .O(N__4957),
            .I(N__4948));
    Sp12to4 I__1005 (
            .O(N__4954),
            .I(N__4943));
    LocalMux I__1004 (
            .O(N__4951),
            .I(N__4943));
    Sp12to4 I__1003 (
            .O(N__4948),
            .I(N__4938));
    Span12Mux_h I__1002 (
            .O(N__4943),
            .I(N__4938));
    Span12Mux_v I__1001 (
            .O(N__4938),
            .I(N__4935));
    Odrv12 I__1000 (
            .O(N__4935),
            .I(PORTSIZE_c));
    IoInMux I__999 (
            .O(N__4932),
            .I(N__4926));
    IoInMux I__998 (
            .O(N__4931),
            .I(N__4923));
    IoInMux I__997 (
            .O(N__4930),
            .I(N__4920));
    IoInMux I__996 (
            .O(N__4929),
            .I(N__4911));
    LocalMux I__995 (
            .O(N__4926),
            .I(N__4902));
    LocalMux I__994 (
            .O(N__4923),
            .I(N__4902));
    LocalMux I__993 (
            .O(N__4920),
            .I(N__4902));
    IoInMux I__992 (
            .O(N__4919),
            .I(N__4899));
    IoInMux I__991 (
            .O(N__4918),
            .I(N__4896));
    IoInMux I__990 (
            .O(N__4917),
            .I(N__4893));
    IoInMux I__989 (
            .O(N__4916),
            .I(N__4886));
    IoInMux I__988 (
            .O(N__4915),
            .I(N__4883));
    IoInMux I__987 (
            .O(N__4914),
            .I(N__4880));
    LocalMux I__986 (
            .O(N__4911),
            .I(N__4873));
    IoInMux I__985 (
            .O(N__4910),
            .I(N__4870));
    IoInMux I__984 (
            .O(N__4909),
            .I(N__4867));
    IoSpan4Mux I__983 (
            .O(N__4902),
            .I(N__4854));
    LocalMux I__982 (
            .O(N__4899),
            .I(N__4854));
    LocalMux I__981 (
            .O(N__4896),
            .I(N__4854));
    LocalMux I__980 (
            .O(N__4893),
            .I(N__4854));
    IoInMux I__979 (
            .O(N__4892),
            .I(N__4851));
    IoInMux I__978 (
            .O(N__4891),
            .I(N__4848));
    IoInMux I__977 (
            .O(N__4890),
            .I(N__4845));
    IoInMux I__976 (
            .O(N__4889),
            .I(N__4842));
    LocalMux I__975 (
            .O(N__4886),
            .I(N__4835));
    LocalMux I__974 (
            .O(N__4883),
            .I(N__4830));
    LocalMux I__973 (
            .O(N__4880),
            .I(N__4830));
    IoInMux I__972 (
            .O(N__4879),
            .I(N__4827));
    IoInMux I__971 (
            .O(N__4878),
            .I(N__4824));
    IoInMux I__970 (
            .O(N__4877),
            .I(N__4821));
    IoInMux I__969 (
            .O(N__4876),
            .I(N__4818));
    IoSpan4Mux I__968 (
            .O(N__4873),
            .I(N__4811));
    LocalMux I__967 (
            .O(N__4870),
            .I(N__4811));
    LocalMux I__966 (
            .O(N__4867),
            .I(N__4811));
    IoInMux I__965 (
            .O(N__4866),
            .I(N__4808));
    IoInMux I__964 (
            .O(N__4865),
            .I(N__4805));
    IoInMux I__963 (
            .O(N__4864),
            .I(N__4802));
    IoInMux I__962 (
            .O(N__4863),
            .I(N__4799));
    IoSpan4Mux I__961 (
            .O(N__4854),
            .I(N__4788));
    LocalMux I__960 (
            .O(N__4851),
            .I(N__4788));
    LocalMux I__959 (
            .O(N__4848),
            .I(N__4788));
    LocalMux I__958 (
            .O(N__4845),
            .I(N__4788));
    LocalMux I__957 (
            .O(N__4842),
            .I(N__4788));
    IoInMux I__956 (
            .O(N__4841),
            .I(N__4785));
    IoInMux I__955 (
            .O(N__4840),
            .I(N__4782));
    IoInMux I__954 (
            .O(N__4839),
            .I(N__4779));
    IoInMux I__953 (
            .O(N__4838),
            .I(N__4776));
    IoSpan4Mux I__952 (
            .O(N__4835),
            .I(N__4772));
    IoSpan4Mux I__951 (
            .O(N__4830),
            .I(N__4761));
    LocalMux I__950 (
            .O(N__4827),
            .I(N__4761));
    LocalMux I__949 (
            .O(N__4824),
            .I(N__4761));
    LocalMux I__948 (
            .O(N__4821),
            .I(N__4761));
    LocalMux I__947 (
            .O(N__4818),
            .I(N__4761));
    IoSpan4Mux I__946 (
            .O(N__4811),
            .I(N__4750));
    LocalMux I__945 (
            .O(N__4808),
            .I(N__4750));
    LocalMux I__944 (
            .O(N__4805),
            .I(N__4750));
    LocalMux I__943 (
            .O(N__4802),
            .I(N__4750));
    LocalMux I__942 (
            .O(N__4799),
            .I(N__4750));
    IoSpan4Mux I__941 (
            .O(N__4788),
            .I(N__4739));
    LocalMux I__940 (
            .O(N__4785),
            .I(N__4739));
    LocalMux I__939 (
            .O(N__4782),
            .I(N__4739));
    LocalMux I__938 (
            .O(N__4779),
            .I(N__4739));
    LocalMux I__937 (
            .O(N__4776),
            .I(N__4739));
    IoInMux I__936 (
            .O(N__4775),
            .I(N__4736));
    Span4Mux_s0_h I__935 (
            .O(N__4772),
            .I(N__4731));
    IoSpan4Mux I__934 (
            .O(N__4761),
            .I(N__4728));
    IoSpan4Mux I__933 (
            .O(N__4750),
            .I(N__4721));
    IoSpan4Mux I__932 (
            .O(N__4739),
            .I(N__4721));
    LocalMux I__931 (
            .O(N__4736),
            .I(N__4721));
    IoInMux I__930 (
            .O(N__4735),
            .I(N__4718));
    IoInMux I__929 (
            .O(N__4734),
            .I(N__4715));
    Span4Mux_h I__928 (
            .O(N__4731),
            .I(N__4712));
    Span4Mux_s3_v I__927 (
            .O(N__4728),
            .I(N__4709));
    IoSpan4Mux I__926 (
            .O(N__4721),
            .I(N__4705));
    LocalMux I__925 (
            .O(N__4718),
            .I(N__4700));
    LocalMux I__924 (
            .O(N__4715),
            .I(N__4700));
    Span4Mux_h I__923 (
            .O(N__4712),
            .I(N__4695));
    Span4Mux_v I__922 (
            .O(N__4709),
            .I(N__4695));
    IoInMux I__921 (
            .O(N__4708),
            .I(N__4692));
    Sp12to4 I__920 (
            .O(N__4705),
            .I(N__4689));
    Span12Mux_s8_h I__919 (
            .O(N__4700),
            .I(N__4686));
    Sp12to4 I__918 (
            .O(N__4695),
            .I(N__4683));
    LocalMux I__917 (
            .O(N__4692),
            .I(N__4680));
    Span12Mux_h I__916 (
            .O(N__4689),
            .I(N__4677));
    Span12Mux_v I__915 (
            .O(N__4686),
            .I(N__4670));
    Span12Mux_v I__914 (
            .O(N__4683),
            .I(N__4670));
    Span12Mux_s8_h I__913 (
            .O(N__4680),
            .I(N__4670));
    Odrv12 I__912 (
            .O(N__4677),
            .I(U111_CYCLE_SM_OFFBOARD_EN_0));
    Odrv12 I__911 (
            .O(N__4670),
            .I(U111_CYCLE_SM_OFFBOARD_EN_0));
    CascadeMux I__910 (
            .O(N__4665),
            .I(\U111_CYCLE_SM.un4_TS_OUT_i_0_cascade_ ));
    InMux I__909 (
            .O(N__4662),
            .I(N__4659));
    LocalMux I__908 (
            .O(N__4659),
            .I(\U111_CYCLE_SM.N_106 ));
    CascadeMux I__907 (
            .O(N__4656),
            .I(N__4653));
    InMux I__906 (
            .O(N__4653),
            .I(N__4650));
    LocalMux I__905 (
            .O(N__4650),
            .I(N__4647));
    Span4Mux_v I__904 (
            .O(N__4647),
            .I(N__4637));
    InMux I__903 (
            .O(N__4646),
            .I(N__4634));
    InMux I__902 (
            .O(N__4645),
            .I(N__4631));
    InMux I__901 (
            .O(N__4644),
            .I(N__4624));
    InMux I__900 (
            .O(N__4643),
            .I(N__4624));
    InMux I__899 (
            .O(N__4642),
            .I(N__4624));
    InMux I__898 (
            .O(N__4641),
            .I(N__4619));
    InMux I__897 (
            .O(N__4640),
            .I(N__4619));
    Sp12to4 I__896 (
            .O(N__4637),
            .I(N__4612));
    LocalMux I__895 (
            .O(N__4634),
            .I(N__4612));
    LocalMux I__894 (
            .O(N__4631),
            .I(N__4612));
    LocalMux I__893 (
            .O(N__4624),
            .I(N__4607));
    LocalMux I__892 (
            .O(N__4619),
            .I(N__4607));
    Span12Mux_h I__891 (
            .O(N__4612),
            .I(N__4604));
    Span12Mux_v I__890 (
            .O(N__4607),
            .I(N__4601));
    Span12Mux_v I__889 (
            .O(N__4604),
            .I(N__4598));
    Odrv12 I__888 (
            .O(N__4601),
            .I(RESETn_c));
    Odrv12 I__887 (
            .O(N__4598),
            .I(RESETn_c));
    InMux I__886 (
            .O(N__4593),
            .I(N__4590));
    LocalMux I__885 (
            .O(N__4590),
            .I(\U111_CYCLE_SM.N_140 ));
    InMux I__884 (
            .O(N__4587),
            .I(N__4582));
    InMux I__883 (
            .O(N__4586),
            .I(N__4579));
    InMux I__882 (
            .O(N__4585),
            .I(N__4576));
    LocalMux I__881 (
            .O(N__4582),
            .I(\U111_CYCLE_SM.N_107 ));
    LocalMux I__880 (
            .O(N__4579),
            .I(\U111_CYCLE_SM.N_107 ));
    LocalMux I__879 (
            .O(N__4576),
            .I(\U111_CYCLE_SM.N_107 ));
    InMux I__878 (
            .O(N__4569),
            .I(N__4560));
    InMux I__877 (
            .O(N__4568),
            .I(N__4560));
    InMux I__876 (
            .O(N__4567),
            .I(N__4553));
    InMux I__875 (
            .O(N__4566),
            .I(N__4553));
    InMux I__874 (
            .O(N__4565),
            .I(N__4553));
    LocalMux I__873 (
            .O(N__4560),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    LocalMux I__872 (
            .O(N__4553),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ));
    IoInMux I__871 (
            .O(N__4548),
            .I(N__4544));
    CascadeMux I__870 (
            .O(N__4547),
            .I(N__4539));
    LocalMux I__869 (
            .O(N__4544),
            .I(N__4534));
    InMux I__868 (
            .O(N__4543),
            .I(N__4531));
    InMux I__867 (
            .O(N__4542),
            .I(N__4524));
    InMux I__866 (
            .O(N__4539),
            .I(N__4524));
    InMux I__865 (
            .O(N__4538),
            .I(N__4524));
    CascadeMux I__864 (
            .O(N__4537),
            .I(N__4521));
    Span4Mux_s1_v I__863 (
            .O(N__4534),
            .I(N__4516));
    LocalMux I__862 (
            .O(N__4531),
            .I(N__4511));
    LocalMux I__861 (
            .O(N__4524),
            .I(N__4511));
    InMux I__860 (
            .O(N__4521),
            .I(N__4506));
    InMux I__859 (
            .O(N__4520),
            .I(N__4506));
    CascadeMux I__858 (
            .O(N__4519),
            .I(N__4503));
    Span4Mux_v I__857 (
            .O(N__4516),
            .I(N__4500));
    Span4Mux_v I__856 (
            .O(N__4511),
            .I(N__4497));
    LocalMux I__855 (
            .O(N__4506),
            .I(N__4494));
    InMux I__854 (
            .O(N__4503),
            .I(N__4491));
    Sp12to4 I__853 (
            .O(N__4500),
            .I(N__4487));
    Span4Mux_h I__852 (
            .O(N__4497),
            .I(N__4484));
    Span4Mux_h I__851 (
            .O(N__4494),
            .I(N__4481));
    LocalMux I__850 (
            .O(N__4491),
            .I(N__4478));
    InMux I__849 (
            .O(N__4490),
            .I(N__4475));
    Span12Mux_h I__848 (
            .O(N__4487),
            .I(N__4472));
    Sp12to4 I__847 (
            .O(N__4484),
            .I(N__4469));
    Span4Mux_v I__846 (
            .O(N__4481),
            .I(N__4466));
    Span4Mux_h I__845 (
            .O(N__4478),
            .I(N__4463));
    LocalMux I__844 (
            .O(N__4475),
            .I(N__4460));
    Span12Mux_v I__843 (
            .O(N__4472),
            .I(N__4449));
    Span12Mux_h I__842 (
            .O(N__4469),
            .I(N__4449));
    Sp12to4 I__841 (
            .O(N__4466),
            .I(N__4449));
    Sp12to4 I__840 (
            .O(N__4463),
            .I(N__4449));
    Span12Mux_h I__839 (
            .O(N__4460),
            .I(N__4449));
    Span12Mux_v I__838 (
            .O(N__4449),
            .I(N__4446));
    Odrv12 I__837 (
            .O(N__4446),
            .I(TACKn_in));
    InMux I__836 (
            .O(N__4443),
            .I(N__4440));
    LocalMux I__835 (
            .O(N__4440),
            .I(N__4437));
    Span12Mux_v I__834 (
            .O(N__4437),
            .I(N__4434));
    Odrv12 I__833 (
            .O(N__4434),
            .I(D_LM_AMIGA_in_4));
    IoInMux I__832 (
            .O(N__4431),
            .I(N__4428));
    LocalMux I__831 (
            .O(N__4428),
            .I(N__4425));
    IoSpan4Mux I__830 (
            .O(N__4425),
            .I(N__4422));
    Span4Mux_s3_h I__829 (
            .O(N__4422),
            .I(N__4419));
    Span4Mux_v I__828 (
            .O(N__4419),
            .I(N__4416));
    Span4Mux_h I__827 (
            .O(N__4416),
            .I(N__4413));
    Sp12to4 I__826 (
            .O(N__4413),
            .I(N__4410));
    Odrv12 I__825 (
            .O(N__4410),
            .I(N_118));
    CascadeMux I__824 (
            .O(N__4407),
            .I(N__4404));
    InMux I__823 (
            .O(N__4404),
            .I(N__4401));
    LocalMux I__822 (
            .O(N__4401),
            .I(N__4396));
    InMux I__821 (
            .O(N__4400),
            .I(N__4393));
    InMux I__820 (
            .O(N__4399),
            .I(N__4390));
    Span4Mux_h I__819 (
            .O(N__4396),
            .I(N__4385));
    LocalMux I__818 (
            .O(N__4393),
            .I(N__4385));
    LocalMux I__817 (
            .O(N__4390),
            .I(N__4382));
    Span4Mux_v I__816 (
            .O(N__4385),
            .I(N__4379));
    Sp12to4 I__815 (
            .O(N__4382),
            .I(N__4376));
    Sp12to4 I__814 (
            .O(N__4379),
            .I(N__4373));
    Span12Mux_v I__813 (
            .O(N__4376),
            .I(N__4370));
    Span12Mux_h I__812 (
            .O(N__4373),
            .I(N__4367));
    Odrv12 I__811 (
            .O(N__4370),
            .I(D_UM_AMIGA_in_1));
    Odrv12 I__810 (
            .O(N__4367),
            .I(D_UM_AMIGA_in_1));
    InMux I__809 (
            .O(N__4362),
            .I(N__4359));
    LocalMux I__808 (
            .O(N__4359),
            .I(N__4355));
    InMux I__807 (
            .O(N__4358),
            .I(N__4352));
    Odrv12 I__806 (
            .O(N__4355),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ));
    LocalMux I__805 (
            .O(N__4352),
            .I(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ));
    IoInMux I__804 (
            .O(N__4347),
            .I(N__4344));
    LocalMux I__803 (
            .O(N__4344),
            .I(N__4341));
    IoSpan4Mux I__802 (
            .O(N__4341),
            .I(N__4338));
    IoSpan4Mux I__801 (
            .O(N__4338),
            .I(N__4335));
    Sp12to4 I__800 (
            .O(N__4335),
            .I(N__4332));
    Span12Mux_s9_h I__799 (
            .O(N__4332),
            .I(N__4329));
    Odrv12 I__798 (
            .O(N__4329),
            .I(un1_D_UM_AMIGA_1));
    InMux I__797 (
            .O(N__4326),
            .I(N__4323));
    LocalMux I__796 (
            .O(N__4323),
            .I(N__4320));
    Span4Mux_h I__795 (
            .O(N__4320),
            .I(N__4317));
    Span4Mux_v I__794 (
            .O(N__4317),
            .I(N__4314));
    Sp12to4 I__793 (
            .O(N__4314),
            .I(N__4311));
    Odrv12 I__792 (
            .O(N__4311),
            .I(D_LM_AMIGA_in_6));
    IoInMux I__791 (
            .O(N__4308),
            .I(N__4305));
    LocalMux I__790 (
            .O(N__4305),
            .I(N__4302));
    Span12Mux_s10_h I__789 (
            .O(N__4302),
            .I(N__4299));
    Odrv12 I__788 (
            .O(N__4299),
            .I(N_116));
    IoInMux I__787 (
            .O(N__4296),
            .I(N__4293));
    LocalMux I__786 (
            .O(N__4293),
            .I(N__4290));
    Span12Mux_s6_v I__785 (
            .O(N__4290),
            .I(N__4287));
    Odrv12 I__784 (
            .O(N__4287),
            .I(N_102_i));
    IoInMux I__783 (
            .O(N__4284),
            .I(N__4281));
    LocalMux I__782 (
            .O(N__4281),
            .I(N__4278));
    IoSpan4Mux I__781 (
            .O(N__4278),
            .I(N__4275));
    Span4Mux_s3_v I__780 (
            .O(N__4275),
            .I(N__4272));
    Span4Mux_h I__779 (
            .O(N__4272),
            .I(N__4269));
    Odrv4 I__778 (
            .O(N__4269),
            .I(BUFDIR_c));
    InMux I__777 (
            .O(N__4266),
            .I(N__4257));
    InMux I__776 (
            .O(N__4265),
            .I(N__4257));
    InMux I__775 (
            .O(N__4264),
            .I(N__4257));
    LocalMux I__774 (
            .O(N__4257),
            .I(N__4254));
    Span4Mux_h I__773 (
            .O(N__4254),
            .I(N__4251));
    Span4Mux_v I__772 (
            .O(N__4251),
            .I(N__4248));
    Odrv4 I__771 (
            .O(N__4248),
            .I(BBn_c));
    IoInMux I__770 (
            .O(N__4245),
            .I(N__4242));
    LocalMux I__769 (
            .O(N__4242),
            .I(N__4239));
    Span4Mux_s3_v I__768 (
            .O(N__4239),
            .I(N__4236));
    Span4Mux_h I__767 (
            .O(N__4236),
            .I(N__4233));
    Odrv4 I__766 (
            .O(N__4233),
            .I(N_104));
    CascadeMux I__765 (
            .O(N__4230),
            .I(N__4226));
    InMux I__764 (
            .O(N__4229),
            .I(N__4223));
    InMux I__763 (
            .O(N__4226),
            .I(N__4220));
    LocalMux I__762 (
            .O(N__4223),
            .I(N__4217));
    LocalMux I__761 (
            .O(N__4220),
            .I(N__4214));
    Span4Mux_v I__760 (
            .O(N__4217),
            .I(N__4210));
    Span4Mux_v I__759 (
            .O(N__4214),
            .I(N__4207));
    InMux I__758 (
            .O(N__4213),
            .I(N__4204));
    Span4Mux_v I__757 (
            .O(N__4210),
            .I(N__4201));
    Span4Mux_v I__756 (
            .O(N__4207),
            .I(N__4196));
    LocalMux I__755 (
            .O(N__4204),
            .I(N__4196));
    Span4Mux_v I__754 (
            .O(N__4201),
            .I(N__4193));
    Span4Mux_v I__753 (
            .O(N__4196),
            .I(N__4190));
    Sp12to4 I__752 (
            .O(N__4193),
            .I(N__4185));
    Sp12to4 I__751 (
            .O(N__4190),
            .I(N__4185));
    Span12Mux_h I__750 (
            .O(N__4185),
            .I(N__4182));
    Odrv12 I__749 (
            .O(N__4182),
            .I(D_UU_AMIGA_in_3));
    InMux I__748 (
            .O(N__4179),
            .I(N__4176));
    LocalMux I__747 (
            .O(N__4176),
            .I(N__4173));
    Span4Mux_v I__746 (
            .O(N__4173),
            .I(N__4170));
    Span4Mux_v I__745 (
            .O(N__4170),
            .I(N__4166));
    InMux I__744 (
            .O(N__4169),
            .I(N__4163));
    Odrv4 I__743 (
            .O(N__4166),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ));
    LocalMux I__742 (
            .O(N__4163),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ));
    IoInMux I__741 (
            .O(N__4158),
            .I(N__4155));
    LocalMux I__740 (
            .O(N__4155),
            .I(N__4152));
    Span4Mux_s2_v I__739 (
            .O(N__4152),
            .I(N__4149));
    Span4Mux_v I__738 (
            .O(N__4149),
            .I(N__4146));
    Sp12to4 I__737 (
            .O(N__4146),
            .I(N__4143));
    Span12Mux_s10_h I__736 (
            .O(N__4143),
            .I(N__4140));
    Odrv12 I__735 (
            .O(N__4140),
            .I(N_128));
    InMux I__734 (
            .O(N__4137),
            .I(N__4134));
    LocalMux I__733 (
            .O(N__4134),
            .I(\U111_CYCLE_SM.N_195 ));
    InMux I__732 (
            .O(N__4131),
            .I(N__4128));
    LocalMux I__731 (
            .O(N__4128),
            .I(\U111_CYCLE_SM.N_132 ));
    CascadeMux I__730 (
            .O(N__4125),
            .I(N__4121));
    InMux I__729 (
            .O(N__4124),
            .I(N__4118));
    InMux I__728 (
            .O(N__4121),
            .I(N__4115));
    LocalMux I__727 (
            .O(N__4118),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ));
    LocalMux I__726 (
            .O(N__4115),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ));
    InMux I__725 (
            .O(N__4110),
            .I(N__4106));
    InMux I__724 (
            .O(N__4109),
            .I(N__4103));
    LocalMux I__723 (
            .O(N__4106),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    LocalMux I__722 (
            .O(N__4103),
            .I(\U111_CYCLE_SM.TS_ENZ0 ));
    IoInMux I__721 (
            .O(N__4098),
            .I(N__4095));
    LocalMux I__720 (
            .O(N__4095),
            .I(N__4092));
    Span4Mux_s3_v I__719 (
            .O(N__4092),
            .I(N__4089));
    Sp12to4 I__718 (
            .O(N__4089),
            .I(N__4086));
    Span12Mux_h I__717 (
            .O(N__4086),
            .I(N__4083));
    Odrv12 I__716 (
            .O(N__4083),
            .I(TS_OUT));
    InMux I__715 (
            .O(N__4080),
            .I(N__4077));
    LocalMux I__714 (
            .O(N__4077),
            .I(N__4074));
    Span4Mux_v I__713 (
            .O(N__4074),
            .I(N__4071));
    Sp12to4 I__712 (
            .O(N__4071),
            .I(N__4067));
    IoInMux I__711 (
            .O(N__4070),
            .I(N__4064));
    Span12Mux_h I__710 (
            .O(N__4067),
            .I(N__4061));
    LocalMux I__709 (
            .O(N__4064),
            .I(N__4058));
    Span12Mux_v I__708 (
            .O(N__4061),
            .I(N__4055));
    IoSpan4Mux I__707 (
            .O(N__4058),
            .I(N__4052));
    Odrv12 I__706 (
            .O(N__4055),
            .I(TBIn_c));
    Odrv4 I__705 (
            .O(N__4052),
            .I(TBIn_c));
    InMux I__704 (
            .O(N__4047),
            .I(N__4039));
    InMux I__703 (
            .O(N__4046),
            .I(N__4039));
    InMux I__702 (
            .O(N__4045),
            .I(N__4034));
    InMux I__701 (
            .O(N__4044),
            .I(N__4034));
    LocalMux I__700 (
            .O(N__4039),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    LocalMux I__699 (
            .O(N__4034),
            .I(\U111_CYCLE_SM.BURSTZ0 ));
    CascadeMux I__698 (
            .O(N__4029),
            .I(N__4024));
    InMux I__697 (
            .O(N__4028),
            .I(N__4019));
    InMux I__696 (
            .O(N__4027),
            .I(N__4019));
    InMux I__695 (
            .O(N__4024),
            .I(N__4016));
    LocalMux I__694 (
            .O(N__4019),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    LocalMux I__693 (
            .O(N__4016),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ));
    InMux I__692 (
            .O(N__4011),
            .I(N__4007));
    InMux I__691 (
            .O(N__4010),
            .I(N__4004));
    LocalMux I__690 (
            .O(N__4007),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ));
    LocalMux I__689 (
            .O(N__4004),
            .I(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ));
    InMux I__688 (
            .O(N__3999),
            .I(N__3996));
    LocalMux I__687 (
            .O(N__3996),
            .I(\U111_CYCLE_SM.N_109 ));
    CascadeMux I__686 (
            .O(N__3993),
            .I(\U111_CYCLE_SM.N_109_cascade_ ));
    InMux I__685 (
            .O(N__3990),
            .I(N__3984));
    InMux I__684 (
            .O(N__3989),
            .I(N__3979));
    InMux I__683 (
            .O(N__3988),
            .I(N__3979));
    InMux I__682 (
            .O(N__3987),
            .I(N__3976));
    LocalMux I__681 (
            .O(N__3984),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    LocalMux I__680 (
            .O(N__3979),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    LocalMux I__679 (
            .O(N__3976),
            .I(\U111_CYCLE_SM.PORT_MISMATCHZ0 ));
    InMux I__678 (
            .O(N__3969),
            .I(N__3966));
    LocalMux I__677 (
            .O(N__3966),
            .I(N__3963));
    Span12Mux_v I__676 (
            .O(N__3963),
            .I(N__3960));
    Odrv12 I__675 (
            .O(N__3960),
            .I(D_LM_AMIGA_in_5));
    IoInMux I__674 (
            .O(N__3957),
            .I(N__3954));
    LocalMux I__673 (
            .O(N__3954),
            .I(N__3951));
    Span4Mux_s3_h I__672 (
            .O(N__3951),
            .I(N__3948));
    Span4Mux_v I__671 (
            .O(N__3948),
            .I(N__3945));
    Sp12to4 I__670 (
            .O(N__3945),
            .I(N__3942));
    Span12Mux_h I__669 (
            .O(N__3942),
            .I(N__3939));
    Odrv12 I__668 (
            .O(N__3939),
            .I(N_117));
    CascadeMux I__667 (
            .O(N__3936),
            .I(\U111_CYCLE_SM.N_144_cascade_ ));
    InMux I__666 (
            .O(N__3933),
            .I(N__3930));
    LocalMux I__665 (
            .O(N__3930),
            .I(\U111_CYCLE_SM.N_142 ));
    InMux I__664 (
            .O(N__3927),
            .I(N__3923));
    InMux I__663 (
            .O(N__3926),
            .I(N__3920));
    LocalMux I__662 (
            .O(N__3923),
            .I(\U111_CYCLE_SM.N_197 ));
    LocalMux I__661 (
            .O(N__3920),
            .I(\U111_CYCLE_SM.N_197 ));
    CascadeMux I__660 (
            .O(N__3915),
            .I(N__3908));
    InMux I__659 (
            .O(N__3914),
            .I(N__3903));
    InMux I__658 (
            .O(N__3913),
            .I(N__3903));
    InMux I__657 (
            .O(N__3912),
            .I(N__3896));
    InMux I__656 (
            .O(N__3911),
            .I(N__3896));
    InMux I__655 (
            .O(N__3908),
            .I(N__3896));
    LocalMux I__654 (
            .O(N__3903),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    LocalMux I__653 (
            .O(N__3896),
            .I(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ));
    CascadeMux I__652 (
            .O(N__3891),
            .I(\U111_CYCLE_SM.N_195_cascade_ ));
    InMux I__651 (
            .O(N__3888),
            .I(N__3885));
    LocalMux I__650 (
            .O(N__3885),
            .I(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_1_0 ));
    InMux I__649 (
            .O(N__3882),
            .I(N__3879));
    LocalMux I__648 (
            .O(N__3879),
            .I(N__3875));
    IoInMux I__647 (
            .O(N__3878),
            .I(N__3872));
    Span4Mux_v I__646 (
            .O(N__3875),
            .I(N__3869));
    LocalMux I__645 (
            .O(N__3872),
            .I(N__3866));
    Span4Mux_h I__644 (
            .O(N__3869),
            .I(N__3863));
    Span4Mux_s3_h I__643 (
            .O(N__3866),
            .I(N__3860));
    Span4Mux_v I__642 (
            .O(N__3863),
            .I(N__3857));
    Sp12to4 I__641 (
            .O(N__3860),
            .I(N__3854));
    Sp12to4 I__640 (
            .O(N__3857),
            .I(N__3851));
    Span12Mux_v I__639 (
            .O(N__3854),
            .I(N__3848));
    Span12Mux_v I__638 (
            .O(N__3851),
            .I(N__3843));
    Span12Mux_h I__637 (
            .O(N__3848),
            .I(N__3843));
    Span12Mux_h I__636 (
            .O(N__3843),
            .I(N__3840));
    Odrv12 I__635 (
            .O(N__3840),
            .I(D_LL_040_in_3));
    InMux I__634 (
            .O(N__3837),
            .I(N__3834));
    LocalMux I__633 (
            .O(N__3834),
            .I(N__3831));
    Span4Mux_v I__632 (
            .O(N__3831),
            .I(N__3828));
    Sp12to4 I__631 (
            .O(N__3828),
            .I(N__3825));
    Span12Mux_h I__630 (
            .O(N__3825),
            .I(N__3822));
    Span12Mux_v I__629 (
            .O(N__3822),
            .I(N__3819));
    Odrv12 I__628 (
            .O(N__3819),
            .I(D_UM_040_in_3));
    IoInMux I__627 (
            .O(N__3816),
            .I(N__3813));
    LocalMux I__626 (
            .O(N__3813),
            .I(N__3810));
    IoSpan4Mux I__625 (
            .O(N__3810),
            .I(N__3807));
    Span4Mux_s2_h I__624 (
            .O(N__3807),
            .I(N__3804));
    Span4Mux_h I__623 (
            .O(N__3804),
            .I(N__3801));
    Span4Mux_h I__622 (
            .O(N__3801),
            .I(N__3798));
    Odrv4 I__621 (
            .O(N__3798),
            .I(un1_D_UM_040_3));
    InMux I__620 (
            .O(N__3795),
            .I(N__3792));
    LocalMux I__619 (
            .O(N__3792),
            .I(N__3789));
    Sp12to4 I__618 (
            .O(N__3789),
            .I(N__3786));
    Span12Mux_v I__617 (
            .O(N__3786),
            .I(N__3783));
    Odrv12 I__616 (
            .O(N__3783),
            .I(D_LM_AMIGA_in_7));
    IoInMux I__615 (
            .O(N__3780),
            .I(N__3777));
    LocalMux I__614 (
            .O(N__3777),
            .I(N__3774));
    IoSpan4Mux I__613 (
            .O(N__3774),
            .I(N__3771));
    Span4Mux_s2_h I__612 (
            .O(N__3771),
            .I(N__3768));
    Sp12to4 I__611 (
            .O(N__3768),
            .I(N__3765));
    Span12Mux_s9_h I__610 (
            .O(N__3765),
            .I(N__3762));
    Odrv12 I__609 (
            .O(N__3762),
            .I(N_115));
    CascadeMux I__608 (
            .O(N__3759),
            .I(N__3756));
    InMux I__607 (
            .O(N__3756),
            .I(N__3753));
    LocalMux I__606 (
            .O(N__3753),
            .I(N__3748));
    InMux I__605 (
            .O(N__3752),
            .I(N__3745));
    InMux I__604 (
            .O(N__3751),
            .I(N__3742));
    Span4Mux_h I__603 (
            .O(N__3748),
            .I(N__3737));
    LocalMux I__602 (
            .O(N__3745),
            .I(N__3737));
    LocalMux I__601 (
            .O(N__3742),
            .I(N__3734));
    Span4Mux_v I__600 (
            .O(N__3737),
            .I(N__3731));
    Span4Mux_v I__599 (
            .O(N__3734),
            .I(N__3728));
    Span4Mux_h I__598 (
            .O(N__3731),
            .I(N__3725));
    IoSpan4Mux I__597 (
            .O(N__3728),
            .I(N__3722));
    Sp12to4 I__596 (
            .O(N__3725),
            .I(N__3719));
    IoSpan4Mux I__595 (
            .O(N__3722),
            .I(N__3716));
    Odrv12 I__594 (
            .O(N__3719),
            .I(D_UU_AMIGA_in_2));
    Odrv4 I__593 (
            .O(N__3716),
            .I(D_UU_AMIGA_in_2));
    InMux I__592 (
            .O(N__3711),
            .I(N__3708));
    LocalMux I__591 (
            .O(N__3708),
            .I(N__3704));
    InMux I__590 (
            .O(N__3707),
            .I(N__3701));
    Odrv12 I__589 (
            .O(N__3704),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ));
    LocalMux I__588 (
            .O(N__3701),
            .I(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ));
    IoInMux I__587 (
            .O(N__3696),
            .I(N__3693));
    LocalMux I__586 (
            .O(N__3693),
            .I(N__3690));
    Span4Mux_s3_v I__585 (
            .O(N__3690),
            .I(N__3687));
    Span4Mux_h I__584 (
            .O(N__3687),
            .I(N__3684));
    Span4Mux_h I__583 (
            .O(N__3684),
            .I(N__3681));
    Span4Mux_h I__582 (
            .O(N__3681),
            .I(N__3678));
    Span4Mux_h I__581 (
            .O(N__3678),
            .I(N__3675));
    Odrv4 I__580 (
            .O(N__3675),
            .I(N_129));
    InMux I__579 (
            .O(N__3672),
            .I(N__3669));
    LocalMux I__578 (
            .O(N__3669),
            .I(N__3666));
    Span4Mux_v I__577 (
            .O(N__3666),
            .I(N__3663));
    Span4Mux_h I__576 (
            .O(N__3663),
            .I(N__3660));
    Sp12to4 I__575 (
            .O(N__3660),
            .I(N__3657));
    Span12Mux_h I__574 (
            .O(N__3657),
            .I(N__3654));
    Odrv12 I__573 (
            .O(N__3654),
            .I(D_UU_040_in_2));
    IoInMux I__572 (
            .O(N__3651),
            .I(N__3647));
    InMux I__571 (
            .O(N__3650),
            .I(N__3644));
    LocalMux I__570 (
            .O(N__3647),
            .I(N__3641));
    LocalMux I__569 (
            .O(N__3644),
            .I(N__3638));
    Span4Mux_s1_h I__568 (
            .O(N__3641),
            .I(N__3635));
    Span4Mux_h I__567 (
            .O(N__3638),
            .I(N__3632));
    Sp12to4 I__566 (
            .O(N__3635),
            .I(N__3629));
    Sp12to4 I__565 (
            .O(N__3632),
            .I(N__3626));
    Span12Mux_v I__564 (
            .O(N__3629),
            .I(N__3623));
    Span12Mux_v I__563 (
            .O(N__3626),
            .I(N__3620));
    Span12Mux_h I__562 (
            .O(N__3623),
            .I(N__3615));
    Span12Mux_v I__561 (
            .O(N__3620),
            .I(N__3615));
    Span12Mux_h I__560 (
            .O(N__3615),
            .I(N__3612));
    Odrv12 I__559 (
            .O(N__3612),
            .I(D_LM_040_in_2));
    IoInMux I__558 (
            .O(N__3609),
            .I(N__3606));
    LocalMux I__557 (
            .O(N__3606),
            .I(N__3603));
    IoSpan4Mux I__556 (
            .O(N__3603),
            .I(N__3600));
    Span4Mux_s2_v I__555 (
            .O(N__3600),
            .I(N__3597));
    Span4Mux_v I__554 (
            .O(N__3597),
            .I(N__3594));
    Odrv4 I__553 (
            .O(N__3594),
            .I(un1_D_UU_040_2));
    IoInMux I__552 (
            .O(N__3591),
            .I(N__3588));
    LocalMux I__551 (
            .O(N__3588),
            .I(N__3585));
    Span12Mux_s11_v I__550 (
            .O(N__3585),
            .I(N__3582));
    Odrv12 I__549 (
            .O(N__3582),
            .I(CPUBGn_c_i_0));
    InMux I__548 (
            .O(N__3579),
            .I(N__3576));
    LocalMux I__547 (
            .O(N__3576),
            .I(N__3573));
    Span12Mux_v I__546 (
            .O(N__3573),
            .I(N__3570));
    Odrv12 I__545 (
            .O(N__3570),
            .I(D_LL_AMIGA_in_7));
    IoInMux I__544 (
            .O(N__3567),
            .I(N__3564));
    LocalMux I__543 (
            .O(N__3564),
            .I(N__3561));
    Span12Mux_s8_h I__542 (
            .O(N__3561),
            .I(N__3558));
    Span12Mux_h I__541 (
            .O(N__3558),
            .I(N__3555));
    Odrv12 I__540 (
            .O(N__3555),
            .I(un2_D_LL_AMIGA_7));
    CascadeMux I__539 (
            .O(N__3552),
            .I(\U111_CYCLE_SM.N_112_cascade_ ));
    InMux I__538 (
            .O(N__3549),
            .I(N__3546));
    LocalMux I__537 (
            .O(N__3546),
            .I(N__3543));
    Span4Mux_v I__536 (
            .O(N__3543),
            .I(N__3540));
    Sp12to4 I__535 (
            .O(N__3540),
            .I(N__3537));
    Odrv12 I__534 (
            .O(N__3537),
            .I(D_LL_AMIGA_in_2));
    IoInMux I__533 (
            .O(N__3534),
            .I(N__3531));
    LocalMux I__532 (
            .O(N__3531),
            .I(N__3528));
    IoSpan4Mux I__531 (
            .O(N__3528),
            .I(N__3525));
    IoSpan4Mux I__530 (
            .O(N__3525),
            .I(N__3522));
    Sp12to4 I__529 (
            .O(N__3522),
            .I(N__3519));
    Span12Mux_s9_h I__528 (
            .O(N__3519),
            .I(N__3516));
    Span12Mux_h I__527 (
            .O(N__3516),
            .I(N__3513));
    Odrv12 I__526 (
            .O(N__3513),
            .I(un2_D_LL_AMIGA_2));
    InMux I__525 (
            .O(N__3510),
            .I(N__3507));
    LocalMux I__524 (
            .O(N__3507),
            .I(N__3504));
    Span4Mux_v I__523 (
            .O(N__3504),
            .I(N__3501));
    Sp12to4 I__522 (
            .O(N__3501),
            .I(N__3498));
    Odrv12 I__521 (
            .O(N__3498),
            .I(D_LL_AMIGA_in_3));
    IoInMux I__520 (
            .O(N__3495),
            .I(N__3492));
    LocalMux I__519 (
            .O(N__3492),
            .I(N__3489));
    Span4Mux_s2_h I__518 (
            .O(N__3489),
            .I(N__3486));
    Span4Mux_v I__517 (
            .O(N__3486),
            .I(N__3483));
    Span4Mux_v I__516 (
            .O(N__3483),
            .I(N__3480));
    Sp12to4 I__515 (
            .O(N__3480),
            .I(N__3477));
    Span12Mux_s11_h I__514 (
            .O(N__3477),
            .I(N__3474));
    Odrv12 I__513 (
            .O(N__3474),
            .I(un2_D_LL_AMIGA_3));
    InMux I__512 (
            .O(N__3471),
            .I(N__3468));
    LocalMux I__511 (
            .O(N__3468),
            .I(N__3465));
    Span4Mux_v I__510 (
            .O(N__3465),
            .I(N__3462));
    Span4Mux_v I__509 (
            .O(N__3462),
            .I(N__3458));
    InMux I__508 (
            .O(N__3461),
            .I(N__3455));
    Sp12to4 I__507 (
            .O(N__3458),
            .I(N__3450));
    LocalMux I__506 (
            .O(N__3455),
            .I(N__3450));
    Span12Mux_h I__505 (
            .O(N__3450),
            .I(N__3447));
    Odrv12 I__504 (
            .O(N__3447),
            .I(A_040_c_1));
    InMux I__503 (
            .O(N__3444),
            .I(N__3441));
    LocalMux I__502 (
            .O(N__3441),
            .I(N__3438));
    Span4Mux_v I__501 (
            .O(N__3438),
            .I(N__3435));
    Sp12to4 I__500 (
            .O(N__3435),
            .I(N__3432));
    Odrv12 I__499 (
            .O(N__3432),
            .I(D_LM_AMIGA_in_0));
    IoInMux I__498 (
            .O(N__3429),
            .I(N__3426));
    LocalMux I__497 (
            .O(N__3426),
            .I(N__3423));
    Span4Mux_s2_h I__496 (
            .O(N__3423),
            .I(N__3420));
    Span4Mux_v I__495 (
            .O(N__3420),
            .I(N__3417));
    Span4Mux_v I__494 (
            .O(N__3417),
            .I(N__3414));
    Sp12to4 I__493 (
            .O(N__3414),
            .I(N__3411));
    Span12Mux_s11_h I__492 (
            .O(N__3411),
            .I(N__3408));
    Odrv12 I__491 (
            .O(N__3408),
            .I(N_122));
    InMux I__490 (
            .O(N__3405),
            .I(N__3399));
    InMux I__489 (
            .O(N__3404),
            .I(N__3399));
    LocalMux I__488 (
            .O(N__3399),
            .I(N__3396));
    Span4Mux_v I__487 (
            .O(N__3396),
            .I(N__3393));
    Span4Mux_v I__486 (
            .O(N__3393),
            .I(N__3390));
    Span4Mux_h I__485 (
            .O(N__3390),
            .I(N__3386));
    InMux I__484 (
            .O(N__3389),
            .I(N__3383));
    Odrv4 I__483 (
            .O(N__3386),
            .I(\U111_CYCLE_SM.A2_ENZ0 ));
    LocalMux I__482 (
            .O(N__3383),
            .I(\U111_CYCLE_SM.A2_ENZ0 ));
    CascadeMux I__481 (
            .O(N__3378),
            .I(N__3375));
    InMux I__480 (
            .O(N__3375),
            .I(N__3372));
    LocalMux I__479 (
            .O(N__3372),
            .I(N__3369));
    Odrv4 I__478 (
            .O(N__3369),
            .I(\U111_CYCLE_SM.N_151 ));
    InMux I__477 (
            .O(N__3366),
            .I(N__3363));
    LocalMux I__476 (
            .O(N__3363),
            .I(N__3360));
    Span4Mux_v I__475 (
            .O(N__3360),
            .I(N__3357));
    Sp12to4 I__474 (
            .O(N__3357),
            .I(N__3354));
    Span12Mux_h I__473 (
            .O(N__3354),
            .I(N__3351));
    Span12Mux_h I__472 (
            .O(N__3351),
            .I(N__3348));
    Span12Mux_v I__471 (
            .O(N__3348),
            .I(N__3345));
    Odrv12 I__470 (
            .O(N__3345),
            .I(D_UM_040_in_1));
    InMux I__469 (
            .O(N__3342),
            .I(N__3338));
    IoInMux I__468 (
            .O(N__3341),
            .I(N__3335));
    LocalMux I__467 (
            .O(N__3338),
            .I(N__3332));
    LocalMux I__466 (
            .O(N__3335),
            .I(N__3329));
    Span4Mux_v I__465 (
            .O(N__3332),
            .I(N__3326));
    Span4Mux_s3_h I__464 (
            .O(N__3329),
            .I(N__3323));
    Span4Mux_v I__463 (
            .O(N__3326),
            .I(N__3320));
    Sp12to4 I__462 (
            .O(N__3323),
            .I(N__3317));
    Sp12to4 I__461 (
            .O(N__3320),
            .I(N__3314));
    Span12Mux_v I__460 (
            .O(N__3317),
            .I(N__3311));
    Span12Mux_v I__459 (
            .O(N__3314),
            .I(N__3308));
    Span12Mux_h I__458 (
            .O(N__3311),
            .I(N__3305));
    Span12Mux_h I__457 (
            .O(N__3308),
            .I(N__3302));
    Span12Mux_h I__456 (
            .O(N__3305),
            .I(N__3299));
    Odrv12 I__455 (
            .O(N__3302),
            .I(D_LL_040_in_1));
    Odrv12 I__454 (
            .O(N__3299),
            .I(D_LL_040_in_1));
    IoInMux I__453 (
            .O(N__3294),
            .I(N__3291));
    LocalMux I__452 (
            .O(N__3291),
            .I(N__3288));
    Span12Mux_s10_h I__451 (
            .O(N__3288),
            .I(N__3285));
    Odrv12 I__450 (
            .O(N__3285),
            .I(un1_D_UM_040_1));
    InMux I__449 (
            .O(N__3282),
            .I(N__3279));
    LocalMux I__448 (
            .O(N__3279),
            .I(N__3276));
    Span4Mux_v I__447 (
            .O(N__3276),
            .I(N__3273));
    Sp12to4 I__446 (
            .O(N__3273),
            .I(N__3270));
    Span12Mux_h I__445 (
            .O(N__3270),
            .I(N__3267));
    Odrv12 I__444 (
            .O(N__3267),
            .I(D_UM_040_in_0));
    IoInMux I__443 (
            .O(N__3264),
            .I(N__3261));
    LocalMux I__442 (
            .O(N__3261),
            .I(N__3257));
    InMux I__441 (
            .O(N__3260),
            .I(N__3254));
    IoSpan4Mux I__440 (
            .O(N__3257),
            .I(N__3251));
    LocalMux I__439 (
            .O(N__3254),
            .I(N__3248));
    Span4Mux_s2_h I__438 (
            .O(N__3251),
            .I(N__3245));
    Span12Mux_v I__437 (
            .O(N__3248),
            .I(N__3242));
    Sp12to4 I__436 (
            .O(N__3245),
            .I(N__3239));
    Span12Mux_v I__435 (
            .O(N__3242),
            .I(N__3236));
    Span12Mux_h I__434 (
            .O(N__3239),
            .I(N__3233));
    Span12Mux_h I__433 (
            .O(N__3236),
            .I(N__3230));
    Span12Mux_h I__432 (
            .O(N__3233),
            .I(N__3227));
    Odrv12 I__431 (
            .O(N__3230),
            .I(D_LL_040_in_0));
    Odrv12 I__430 (
            .O(N__3227),
            .I(D_LL_040_in_0));
    IoInMux I__429 (
            .O(N__3222),
            .I(N__3219));
    LocalMux I__428 (
            .O(N__3219),
            .I(N__3216));
    IoSpan4Mux I__427 (
            .O(N__3216),
            .I(N__3213));
    Span4Mux_s3_h I__426 (
            .O(N__3213),
            .I(N__3210));
    Span4Mux_h I__425 (
            .O(N__3210),
            .I(N__3207));
    Odrv4 I__424 (
            .O(N__3207),
            .I(un1_D_UM_040_0));
    InMux I__423 (
            .O(N__3204),
            .I(N__3201));
    LocalMux I__422 (
            .O(N__3201),
            .I(N__3198));
    Span4Mux_v I__421 (
            .O(N__3198),
            .I(N__3195));
    Sp12to4 I__420 (
            .O(N__3195),
            .I(N__3192));
    Odrv12 I__419 (
            .O(N__3192),
            .I(D_LM_AMIGA_in_3));
    IoInMux I__418 (
            .O(N__3189),
            .I(N__3186));
    LocalMux I__417 (
            .O(N__3186),
            .I(N__3183));
    IoSpan4Mux I__416 (
            .O(N__3183),
            .I(N__3180));
    Span4Mux_s1_h I__415 (
            .O(N__3180),
            .I(N__3177));
    Span4Mux_v I__414 (
            .O(N__3177),
            .I(N__3174));
    Sp12to4 I__413 (
            .O(N__3174),
            .I(N__3171));
    Span12Mux_s10_h I__412 (
            .O(N__3171),
            .I(N__3168));
    Odrv12 I__411 (
            .O(N__3168),
            .I(N_119));
    InMux I__410 (
            .O(N__3165),
            .I(N__3162));
    LocalMux I__409 (
            .O(N__3162),
            .I(N__3159));
    Odrv12 I__408 (
            .O(N__3159),
            .I(D_LM_AMIGA_in_1));
    IoInMux I__407 (
            .O(N__3156),
            .I(N__3153));
    LocalMux I__406 (
            .O(N__3153),
            .I(N__3150));
    Span4Mux_s0_h I__405 (
            .O(N__3150),
            .I(N__3147));
    Sp12to4 I__404 (
            .O(N__3147),
            .I(N__3144));
    Span12Mux_v I__403 (
            .O(N__3144),
            .I(N__3141));
    Span12Mux_h I__402 (
            .O(N__3141),
            .I(N__3138));
    Odrv12 I__401 (
            .O(N__3138),
            .I(N_121));
    IoInMux I__400 (
            .O(N__3135),
            .I(N__3132));
    LocalMux I__399 (
            .O(N__3132),
            .I(N__3128));
    InMux I__398 (
            .O(N__3131),
            .I(N__3125));
    IoSpan4Mux I__397 (
            .O(N__3128),
            .I(N__3122));
    LocalMux I__396 (
            .O(N__3125),
            .I(N__3119));
    Span4Mux_s0_h I__395 (
            .O(N__3122),
            .I(N__3116));
    Span4Mux_v I__394 (
            .O(N__3119),
            .I(N__3113));
    Span4Mux_v I__393 (
            .O(N__3116),
            .I(N__3110));
    Sp12to4 I__392 (
            .O(N__3113),
            .I(N__3107));
    Sp12to4 I__391 (
            .O(N__3110),
            .I(N__3104));
    Span12Mux_h I__390 (
            .O(N__3107),
            .I(N__3101));
    Span12Mux_h I__389 (
            .O(N__3104),
            .I(N__3098));
    Span12Mux_v I__388 (
            .O(N__3101),
            .I(N__3095));
    Span12Mux_h I__387 (
            .O(N__3098),
            .I(N__3092));
    Span12Mux_h I__386 (
            .O(N__3095),
            .I(N__3089));
    Odrv12 I__385 (
            .O(N__3092),
            .I(D_LL_040_in_6));
    Odrv12 I__384 (
            .O(N__3089),
            .I(D_LL_040_in_6));
    InMux I__383 (
            .O(N__3084),
            .I(N__3081));
    LocalMux I__382 (
            .O(N__3081),
            .I(N__3078));
    Span12Mux_v I__381 (
            .O(N__3078),
            .I(N__3075));
    Span12Mux_h I__380 (
            .O(N__3075),
            .I(N__3072));
    Odrv12 I__379 (
            .O(N__3072),
            .I(D_UM_040_in_6));
    IoInMux I__378 (
            .O(N__3069),
            .I(N__3066));
    LocalMux I__377 (
            .O(N__3066),
            .I(N__3063));
    Span12Mux_s4_h I__376 (
            .O(N__3063),
            .I(N__3060));
    Span12Mux_v I__375 (
            .O(N__3060),
            .I(N__3057));
    Odrv12 I__374 (
            .O(N__3057),
            .I(un1_D_UM_040_6));
    InMux I__373 (
            .O(N__3054),
            .I(N__3051));
    LocalMux I__372 (
            .O(N__3051),
            .I(N__3048));
    Odrv12 I__371 (
            .O(N__3048),
            .I(D_LM_AMIGA_in_2));
    IoInMux I__370 (
            .O(N__3045),
            .I(N__3042));
    LocalMux I__369 (
            .O(N__3042),
            .I(N__3039));
    Span12Mux_s11_h I__368 (
            .O(N__3039),
            .I(N__3036));
    Span12Mux_v I__367 (
            .O(N__3036),
            .I(N__3033));
    Odrv12 I__366 (
            .O(N__3033),
            .I(N_120));
    IoInMux I__365 (
            .O(N__3030),
            .I(N__3027));
    LocalMux I__364 (
            .O(N__3027),
            .I(N__3024));
    IoSpan4Mux I__363 (
            .O(N__3024),
            .I(N__3020));
    InMux I__362 (
            .O(N__3023),
            .I(N__3017));
    IoSpan4Mux I__361 (
            .O(N__3020),
            .I(N__3014));
    LocalMux I__360 (
            .O(N__3017),
            .I(N__3011));
    Span4Mux_s2_h I__359 (
            .O(N__3014),
            .I(N__3008));
    Span12Mux_v I__358 (
            .O(N__3011),
            .I(N__3005));
    Sp12to4 I__357 (
            .O(N__3008),
            .I(N__3002));
    Span12Mux_v I__356 (
            .O(N__3005),
            .I(N__2999));
    Span12Mux_h I__355 (
            .O(N__3002),
            .I(N__2996));
    Span12Mux_h I__354 (
            .O(N__2999),
            .I(N__2993));
    Span12Mux_h I__353 (
            .O(N__2996),
            .I(N__2990));
    Odrv12 I__352 (
            .O(N__2993),
            .I(D_LM_040_in_0));
    Odrv12 I__351 (
            .O(N__2990),
            .I(D_LM_040_in_0));
    InMux I__350 (
            .O(N__2985),
            .I(N__2982));
    LocalMux I__349 (
            .O(N__2982),
            .I(N__2979));
    Span4Mux_v I__348 (
            .O(N__2979),
            .I(N__2976));
    Span4Mux_h I__347 (
            .O(N__2976),
            .I(N__2973));
    Sp12to4 I__346 (
            .O(N__2973),
            .I(N__2970));
    Span12Mux_h I__345 (
            .O(N__2970),
            .I(N__2967));
    Odrv12 I__344 (
            .O(N__2967),
            .I(D_UU_040_in_0));
    IoInMux I__343 (
            .O(N__2964),
            .I(N__2961));
    LocalMux I__342 (
            .O(N__2961),
            .I(N__2958));
    IoSpan4Mux I__341 (
            .O(N__2958),
            .I(N__2955));
    Span4Mux_s2_v I__340 (
            .O(N__2955),
            .I(N__2952));
    Span4Mux_v I__339 (
            .O(N__2952),
            .I(N__2949));
    Odrv4 I__338 (
            .O(N__2949),
            .I(un1_D_UU_040_0));
    InMux I__337 (
            .O(N__2946),
            .I(N__2943));
    LocalMux I__336 (
            .O(N__2943),
            .I(N__2940));
    Span4Mux_v I__335 (
            .O(N__2940),
            .I(N__2937));
    Span4Mux_h I__334 (
            .O(N__2937),
            .I(N__2934));
    Sp12to4 I__333 (
            .O(N__2934),
            .I(N__2931));
    Span12Mux_h I__332 (
            .O(N__2931),
            .I(N__2928));
    Odrv12 I__331 (
            .O(N__2928),
            .I(D_UU_040_in_4));
    IoInMux I__330 (
            .O(N__2925),
            .I(N__2922));
    LocalMux I__329 (
            .O(N__2922),
            .I(N__2919));
    Span4Mux_s1_h I__328 (
            .O(N__2919),
            .I(N__2916));
    Sp12to4 I__327 (
            .O(N__2916),
            .I(N__2912));
    InMux I__326 (
            .O(N__2915),
            .I(N__2909));
    Span12Mux_v I__325 (
            .O(N__2912),
            .I(N__2906));
    LocalMux I__324 (
            .O(N__2909),
            .I(N__2903));
    Span12Mux_h I__323 (
            .O(N__2906),
            .I(N__2900));
    Span12Mux_v I__322 (
            .O(N__2903),
            .I(N__2897));
    Span12Mux_h I__321 (
            .O(N__2900),
            .I(N__2894));
    Span12Mux_h I__320 (
            .O(N__2897),
            .I(N__2891));
    Odrv12 I__319 (
            .O(N__2894),
            .I(D_LM_040_in_4));
    Odrv12 I__318 (
            .O(N__2891),
            .I(D_LM_040_in_4));
    IoInMux I__317 (
            .O(N__2886),
            .I(N__2883));
    LocalMux I__316 (
            .O(N__2883),
            .I(N__2880));
    IoSpan4Mux I__315 (
            .O(N__2880),
            .I(N__2877));
    Span4Mux_s3_v I__314 (
            .O(N__2877),
            .I(N__2874));
    Odrv4 I__313 (
            .O(N__2874),
            .I(un1_D_UU_040_4));
    InMux I__312 (
            .O(N__2871),
            .I(N__2868));
    LocalMux I__311 (
            .O(N__2868),
            .I(N__2865));
    Span4Mux_v I__310 (
            .O(N__2865),
            .I(N__2862));
    Sp12to4 I__309 (
            .O(N__2862),
            .I(N__2859));
    Span12Mux_h I__308 (
            .O(N__2859),
            .I(N__2856));
    Span12Mux_h I__307 (
            .O(N__2856),
            .I(N__2853));
    Odrv12 I__306 (
            .O(N__2853),
            .I(D_UU_040_in_6));
    IoInMux I__305 (
            .O(N__2850),
            .I(N__2847));
    LocalMux I__304 (
            .O(N__2847),
            .I(N__2844));
    Span4Mux_s2_h I__303 (
            .O(N__2844),
            .I(N__2840));
    InMux I__302 (
            .O(N__2843),
            .I(N__2837));
    Span4Mux_h I__301 (
            .O(N__2840),
            .I(N__2834));
    LocalMux I__300 (
            .O(N__2837),
            .I(N__2831));
    Span4Mux_h I__299 (
            .O(N__2834),
            .I(N__2826));
    Span4Mux_v I__298 (
            .O(N__2831),
            .I(N__2826));
    Span4Mux_v I__297 (
            .O(N__2826),
            .I(N__2823));
    Sp12to4 I__296 (
            .O(N__2823),
            .I(N__2820));
    Span12Mux_h I__295 (
            .O(N__2820),
            .I(N__2817));
    Span12Mux_h I__294 (
            .O(N__2817),
            .I(N__2814));
    Odrv12 I__293 (
            .O(N__2814),
            .I(D_LM_040_in_6));
    IoInMux I__292 (
            .O(N__2811),
            .I(N__2808));
    LocalMux I__291 (
            .O(N__2808),
            .I(N__2805));
    Span4Mux_s2_v I__290 (
            .O(N__2805),
            .I(N__2802));
    Span4Mux_h I__289 (
            .O(N__2802),
            .I(N__2799));
    Span4Mux_v I__288 (
            .O(N__2799),
            .I(N__2796));
    Odrv4 I__287 (
            .O(N__2796),
            .I(un1_D_UU_040_6));
    IoInMux I__286 (
            .O(N__2793),
            .I(N__2790));
    LocalMux I__285 (
            .O(N__2790),
            .I(N__2787));
    Span4Mux_s0_v I__284 (
            .O(N__2787),
            .I(N__2784));
    Sp12to4 I__283 (
            .O(N__2784),
            .I(N__2781));
    Span12Mux_h I__282 (
            .O(N__2781),
            .I(N__2778));
    Span12Mux_v I__281 (
            .O(N__2778),
            .I(N__2775));
    Span12Mux_v I__280 (
            .O(N__2775),
            .I(N__2772));
    Odrv12 I__279 (
            .O(N__2772),
            .I(TAn_in));
    IoInMux I__278 (
            .O(N__2769),
            .I(N__2766));
    LocalMux I__277 (
            .O(N__2766),
            .I(N__2763));
    Odrv12 I__276 (
            .O(N__2763),
            .I(RESETn_c_i));
    IoInMux I__275 (
            .O(N__2760),
            .I(N__2757));
    LocalMux I__274 (
            .O(N__2757),
            .I(N__2754));
    Odrv12 I__273 (
            .O(N__2754),
            .I(U111_CYCLE_SM_A_AMIGA_0_i_1));
    InMux I__272 (
            .O(N__2751),
            .I(N__2748));
    LocalMux I__271 (
            .O(N__2748),
            .I(N__2745));
    Span4Mux_h I__270 (
            .O(N__2745),
            .I(N__2742));
    Span4Mux_v I__269 (
            .O(N__2742),
            .I(N__2739));
    Odrv4 I__268 (
            .O(N__2739),
            .I(A_040_c_0));
    IoInMux I__267 (
            .O(N__2736),
            .I(N__2733));
    LocalMux I__266 (
            .O(N__2733),
            .I(N__2730));
    Span4Mux_s2_v I__265 (
            .O(N__2730),
            .I(N__2727));
    Span4Mux_v I__264 (
            .O(N__2727),
            .I(N__2724));
    Odrv4 I__263 (
            .O(N__2724),
            .I(A_AMIGA_c_0));
    InMux I__262 (
            .O(N__2721),
            .I(N__2718));
    LocalMux I__261 (
            .O(N__2718),
            .I(N__2715));
    Span4Mux_v I__260 (
            .O(N__2715),
            .I(N__2712));
    Sp12to4 I__259 (
            .O(N__2712),
            .I(N__2709));
    Odrv12 I__258 (
            .O(N__2709),
            .I(D_LL_AMIGA_in_4));
    IoInMux I__257 (
            .O(N__2706),
            .I(N__2703));
    LocalMux I__256 (
            .O(N__2703),
            .I(N__2700));
    Span4Mux_s3_h I__255 (
            .O(N__2700),
            .I(N__2697));
    Sp12to4 I__254 (
            .O(N__2697),
            .I(N__2694));
    Span12Mux_s8_v I__253 (
            .O(N__2694),
            .I(N__2691));
    Span12Mux_h I__252 (
            .O(N__2691),
            .I(N__2688));
    Odrv12 I__251 (
            .O(N__2688),
            .I(un2_D_LL_AMIGA_4));
    InMux I__250 (
            .O(N__2685),
            .I(N__2682));
    LocalMux I__249 (
            .O(N__2682),
            .I(N__2679));
    Span12Mux_v I__248 (
            .O(N__2679),
            .I(N__2676));
    Odrv12 I__247 (
            .O(N__2676),
            .I(D_LL_AMIGA_in_1));
    IoInMux I__246 (
            .O(N__2673),
            .I(N__2670));
    LocalMux I__245 (
            .O(N__2670),
            .I(N__2667));
    IoSpan4Mux I__244 (
            .O(N__2667),
            .I(N__2664));
    Span4Mux_s1_h I__243 (
            .O(N__2664),
            .I(N__2661));
    Span4Mux_v I__242 (
            .O(N__2661),
            .I(N__2658));
    Sp12to4 I__241 (
            .O(N__2658),
            .I(N__2655));
    Span12Mux_s10_h I__240 (
            .O(N__2655),
            .I(N__2652));
    Odrv12 I__239 (
            .O(N__2652),
            .I(un2_D_LL_AMIGA_1));
    IoInMux I__238 (
            .O(N__2649),
            .I(N__2646));
    LocalMux I__237 (
            .O(N__2646),
            .I(N__2643));
    Span4Mux_s1_v I__236 (
            .O(N__2643),
            .I(N__2640));
    Span4Mux_v I__235 (
            .O(N__2640),
            .I(N__2637));
    Sp12to4 I__234 (
            .O(N__2637),
            .I(N__2634));
    Span12Mux_h I__233 (
            .O(N__2634),
            .I(N__2631));
    Span12Mux_v I__232 (
            .O(N__2631),
            .I(N__2628));
    Span12Mux_v I__231 (
            .O(N__2628),
            .I(N__2625));
    Odrv12 I__230 (
            .O(N__2625),
            .I(TSn_in));
    IoInMux I__229 (
            .O(N__2622),
            .I(N__2619));
    LocalMux I__228 (
            .O(N__2619),
            .I(N__2616));
    Span4Mux_s0_h I__227 (
            .O(N__2616),
            .I(N__2613));
    Span4Mux_h I__226 (
            .O(N__2613),
            .I(N__2610));
    Span4Mux_h I__225 (
            .O(N__2610),
            .I(N__2607));
    Sp12to4 I__224 (
            .O(N__2607),
            .I(N__2604));
    Span12Mux_s11_v I__223 (
            .O(N__2604),
            .I(N__2601));
    Span12Mux_v I__222 (
            .O(N__2601),
            .I(N__2598));
    Span12Mux_h I__221 (
            .O(N__2598),
            .I(N__2595));
    Odrv12 I__220 (
            .O(N__2595),
            .I(TCIn_c));
    INV \INVU111_CYCLE_SM.TS_OUTC  (
            .O(\INVU111_CYCLE_SM.TS_OUTC_net ),
            .I(N__6381));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__2769),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_1.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_1.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_1_10_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_1_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4645),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_0  (
            .in0(_gnd_net_),
            .in1(N__3461),
            .in2(_gnd_net_),
            .in3(N__3405),
            .lcout(U111_CYCLE_SM_A_AMIGA_0_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_6  (
            .in0(N__2751),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3404),
            .lcout(A_AMIGA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_6_3_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_6_3_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_6_3_1  (
            .in0(N__2721),
            .in1(N__7585),
            .in2(_gnd_net_),
            .in3(N__7894),
            .lcout(un2_D_LL_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_6_3_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_6_3_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_6_3_4  (
            .in0(N__7893),
            .in1(N__4399),
            .in2(_gnd_net_),
            .in3(N__2685),
            .lcout(un2_D_LL_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_6_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_6_10_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_6_10_1  (
            .in0(N__3282),
            .in1(N__3260),
            .in2(_gnd_net_),
            .in3(N__7751),
            .lcout(un1_D_UM_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_6_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_6_10_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_6_10_4  (
            .in0(N__7753),
            .in1(N__4229),
            .in2(_gnd_net_),
            .in3(N__3204),
            .lcout(N_119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_6_10_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_6_10_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_6_10_6  (
            .in0(N__7752),
            .in1(N__6299),
            .in2(_gnd_net_),
            .in3(N__3165),
            .lcout(N_121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_6_12_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_6_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_6_12_1  (
            .in0(N__7818),
            .in1(N__3131),
            .in2(_gnd_net_),
            .in3(N__3084),
            .lcout(un1_D_UM_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_6_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_6_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_6_12_5  (
            .in0(N__7817),
            .in1(N__3752),
            .in2(_gnd_net_),
            .in3(N__3054),
            .lcout(N_120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_6_20_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_6_20_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_6_20_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_6_20_1  (
            .in0(N__3023),
            .in1(N__2985),
            .in2(_gnd_net_),
            .in3(N__7895),
            .lcout(un1_D_UU_040_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_6_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_6_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_6_20_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_6_20_4  (
            .in0(N__7896),
            .in1(N__2946),
            .in2(_gnd_net_),
            .in3(N__2915),
            .lcout(un1_D_UU_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_6_20_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_6_20_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_6_20_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_6_20_7  (
            .in0(N__2871),
            .in1(N__2843),
            .in2(_gnd_net_),
            .in3(N__7897),
            .lcout(un1_D_UU_040_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_7_3_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_7_3_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_7_3_3  (
            .in0(N__3549),
            .in1(N__6720),
            .in2(_gnd_net_),
            .in3(N__7851),
            .lcout(un2_D_LL_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_7_3_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_7_3_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_7_3_6  (
            .in0(N__7852),
            .in1(N__6080),
            .in2(_gnd_net_),
            .in3(N__3510),
            .lcout(un2_D_LL_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_7_7_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_7_7_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_7_7_4  (
            .in0(N__4960),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3471),
            .lcout(\U111_CYCLE_SM.N_151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_7_7_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_7_7_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_7_7_6  (
            .in0(N__7805),
            .in1(N__6204),
            .in2(_gnd_net_),
            .in3(N__3444),
            .lcout(N_122),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.A2_EN_LC_7_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.A2_EN_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.A2_EN_LC_7_10_1 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \U111_CYCLE_SM.A2_EN_LC_7_10_1  (
            .in0(N__3389),
            .in1(N__3927),
            .in2(_gnd_net_),
            .in3(N__5121),
            .lcout(\U111_CYCLE_SM.A2_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6385),
            .ce(),
            .sr(N__6331));
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_7_10_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.PORT_MISMATCH_LC_7_10_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U111_CYCLE_SM.PORT_MISMATCH_LC_7_10_2  (
            .in0(N__3990),
            .in1(N__6417),
            .in2(N__4977),
            .in3(N__5089),
            .lcout(\U111_CYCLE_SM.PORT_MISMATCHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6385),
            .ce(),
            .sr(N__6331));
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_7_10_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.FLIP_WORD_LC_7_10_6 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_LC_7_10_6  (
            .in0(N__5122),
            .in1(N__7750),
            .in2(N__3378),
            .in3(N__5088),
            .lcout(\U111_CYCLE_SM.FLIP_WORDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6385),
            .ce(),
            .sr(N__6331));
    defparam \U111_CYCLE_SM.UU_LATCHED_2_LC_7_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_2_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_2_LC_7_11_1 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_2_LC_7_11_1  (
            .in0(N__3707),
            .in1(N__6606),
            .in2(N__3759),
            .in3(N__7191),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6382),
            .ce(),
            .sr(N__6332));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_7_15_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_7_15_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_7_15_1  (
            .in0(N__3366),
            .in1(N__3342),
            .in2(_gnd_net_),
            .in3(N__7806),
            .lcout(un1_D_UM_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_7_15_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_7_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_7_15_2  (
            .in0(N__7807),
            .in1(N__3882),
            .in2(_gnd_net_),
            .in3(N__3837),
            .lcout(un1_D_UM_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_7_15_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_7_15_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_7_15_4  (
            .in0(N__7808),
            .in1(N__5527),
            .in2(_gnd_net_),
            .in3(N__3795),
            .lcout(N_115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNINJKT_2_LC_7_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNINJKT_2_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNINJKT_2_LC_7_20_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNINJKT_2_LC_7_20_2  (
            .in0(N__8421),
            .in1(N__3751),
            .in2(_gnd_net_),
            .in3(N__3711),
            .lcout(N_129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_7_20_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_7_20_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_7_20_4  (
            .in0(N__3672),
            .in1(N__3650),
            .in2(_gnd_net_),
            .in3(N__7909),
            .lcout(un1_D_UU_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TSn_iobuf_RNO_LC_8_7_3.C_ON=1'b0;
    defparam TSn_iobuf_RNO_LC_8_7_3.SEQ_MODE=4'b0000;
    defparam TSn_iobuf_RNO_LC_8_7_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 TSn_iobuf_RNO_LC_8_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7230),
            .lcout(CPUBGn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_8_7_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_8_7_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_8_7_4  (
            .in0(N__7871),
            .in1(N__5049),
            .in2(_gnd_net_),
            .in3(N__3579),
            .lcout(un2_D_LL_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_8_9_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_8_9_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_8_9_0  (
            .in0(N__5350),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3914),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_112_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_8_9_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_5_LC_8_9_1 .LUT_INIT=16'b1100110000001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_5_LC_8_9_1  (
            .in0(N__4490),
            .in1(N__4641),
            .in2(N__3552),
            .in3(N__4124),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6386),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_8_9_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_EN_RNO_0_LC_8_9_6 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \U111_CYCLE_SM.TS_EN_RNO_0_LC_8_9_6  (
            .in0(N__5351),
            .in1(N__5114),
            .in2(N__4519),
            .in3(N__3913),
            .lcout(\U111_CYCLE_SM.N_132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_8_9_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_4_LC_8_9_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_4_LC_8_9_7  (
            .in0(N__5115),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4640),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6386),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_8_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_1_LC_8_10_0 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_1_LC_8_10_0  (
            .in0(N__4643),
            .in1(N__3926),
            .in2(N__6465),
            .in3(N__4045),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6383),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_8_10_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_8_10_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_8_10_1  (
            .in0(N__3988),
            .in1(N__4569),
            .in2(N__4547),
            .in3(N__3999),
            .lcout(),
            .ltout(\U111_CYCLE_SM.N_144_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_8_10_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_0_LC_8_10_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_0_LC_8_10_2  (
            .in0(N__4642),
            .in1(N__3933),
            .in2(N__3936),
            .in3(N__3888),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6383),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_8_10_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_8_10_3 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_8_10_3  (
            .in0(N__5381),
            .in1(N__4568),
            .in2(_gnd_net_),
            .in3(N__3912),
            .lcout(\U111_CYCLE_SM.N_142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_8_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_3_LC_8_10_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_3_LC_8_10_4  (
            .in0(N__4644),
            .in1(N__3989),
            .in2(_gnd_net_),
            .in3(N__4587),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6383),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_8_10_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_8_10_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_8_10_5  (
            .in0(N__4538),
            .in1(N__5380),
            .in2(_gnd_net_),
            .in3(N__3911),
            .lcout(\U111_CYCLE_SM.N_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_RNILNBJ_LC_8_10_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_RNILNBJ_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.BURST_RNILNBJ_LC_8_10_6 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \U111_CYCLE_SM.BURST_RNILNBJ_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3915),
            .in3(N__4044),
            .lcout(\U111_CYCLE_SM.N_195 ),
            .ltout(\U111_CYCLE_SM.N_195_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_8_10_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_8_10_7 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_8_10_7  (
            .in0(N__4542),
            .in1(N__6628),
            .in2(N__3891),
            .in3(N__5800),
            .lcout(\U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.BURST_LC_8_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_LC_8_11_0 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \U111_CYCLE_SM.BURST_LC_8_11_0  (
            .in0(N__6534),
            .in1(N__6498),
            .in2(N__6464),
            .in3(N__4047),
            .lcout(\U111_CYCLE_SM.BURSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6380),
            .ce(),
            .sr(N__6333));
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_8_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_COUNT_1_LC_8_11_1 .LUT_INIT=16'b0000110100000010;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_1_LC_8_11_1  (
            .in0(N__4027),
            .in1(N__4586),
            .in2(N__6463),
            .in3(N__4011),
            .lcout(\U111_CYCLE_SM.BURST_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6380),
            .ce(),
            .sr(N__6333));
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_8_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.BURST_COUNT_0_LC_8_11_2 .LUT_INIT=16'b0100010000010001;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_0_LC_8_11_2  (
            .in0(N__6453),
            .in1(N__4585),
            .in2(_gnd_net_),
            .in3(N__4028),
            .lcout(\U111_CYCLE_SM.BURST_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6380),
            .ce(),
            .sr(N__6333));
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_8_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_8_11_4 .LUT_INIT=16'b1111011101110111;
    LogicCell40 \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_8_11_4  (
            .in0(N__4080),
            .in1(N__4046),
            .in2(N__4029),
            .in3(N__4010),
            .lcout(\U111_CYCLE_SM.N_109 ),
            .ltout(\U111_CYCLE_SM.N_109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_2_LC_8_11_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_2_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_1_2_LC_8_11_5 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_1_2_LC_8_11_5  (
            .in0(N__4543),
            .in1(N__5087),
            .in2(N__3993),
            .in3(N__3987),
            .lcout(\U111_CYCLE_SM.N_140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_1_LC_8_12_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_1_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_1_LC_8_12_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_1_LC_8_12_0  (
            .in0(N__4358),
            .in1(N__6600),
            .in2(N__4407),
            .in3(N__7188),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6377),
            .ce(),
            .sr(N__6335));
    defparam \U111_CYCLE_SM.UM_LATCHED_4_LC_8_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_4_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_4_LC_8_12_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_4_LC_8_12_5  (
            .in0(N__7189),
            .in1(N__7601),
            .in2(N__7590),
            .in3(N__6602),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6377),
            .ce(),
            .sr(N__6335));
    defparam \U111_CYCLE_SM.UU_LATCHED_3_LC_8_12_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_3_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_3_LC_8_12_6 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_3_LC_8_12_6  (
            .in0(N__4169),
            .in1(N__6601),
            .in2(N__4230),
            .in3(N__7190),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6377),
            .ce(),
            .sr(N__6335));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_13_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_13_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_13_3  (
            .in0(N__7840),
            .in1(N__5618),
            .in2(_gnd_net_),
            .in3(N__3969),
            .lcout(N_117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_8_13_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_8_13_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_8_13_4  (
            .in0(N__4443),
            .in1(N__5444),
            .in2(_gnd_net_),
            .in3(N__7839),
            .lcout(N_118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_RNI51EL_1_LC_8_15_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNI51EL_1_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNI51EL_1_LC_8_15_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_RNI51EL_1_LC_8_15_5  (
            .in0(N__4400),
            .in1(N__4362),
            .in2(_gnd_net_),
            .in3(N__8397),
            .lcout(un1_D_UM_AMIGA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_15_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_15_6  (
            .in0(N__4326),
            .in1(N__5681),
            .in2(_gnd_net_),
            .in3(N__7883),
            .lcout(N_116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_BUFFERS.N_102_i_LC_8_20_0 .C_ON=1'b0;
    defparam \U111_BUFFERS.N_102_i_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \U111_BUFFERS.N_102_i_LC_8_20_0 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U111_BUFFERS.N_102_i_LC_8_20_0  (
            .in0(N__7258),
            .in1(N__4265),
            .in2(_gnd_net_),
            .in3(N__7449),
            .lcout(N_102_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_BUFFERS.un1_DMA_EN_0_0_LC_8_20_2 .C_ON=1'b0;
    defparam \U111_BUFFERS.un1_DMA_EN_0_0_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_BUFFERS.un1_DMA_EN_0_0_LC_8_20_2 .LUT_INIT=16'b0010001001100110;
    LogicCell40 \U111_BUFFERS.un1_DMA_EN_0_0_LC_8_20_2  (
            .in0(N__7067),
            .in1(N__7257),
            .in2(_gnd_net_),
            .in3(N__4266),
            .lcout(BUFDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_BUFFERS.DMA_EN_i_0_LC_8_20_4 .C_ON=1'b0;
    defparam \U111_BUFFERS.DMA_EN_i_0_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \U111_BUFFERS.DMA_EN_i_0_LC_8_20_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U111_BUFFERS.DMA_EN_i_0_LC_8_20_4  (
            .in0(_gnd_net_),
            .in1(N__7256),
            .in2(_gnd_net_),
            .in3(N__4264),
            .lcout(N_104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIPLKT_3_LC_8_20_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIPLKT_3_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIPLKT_3_LC_8_20_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNIPLKT_3_LC_8_20_6  (
            .in0(N__8423),
            .in1(N__4213),
            .in2(_gnd_net_),
            .in3(N__4179),
            .lcout(N_128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_EN_LC_9_9_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_EN_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TS_EN_LC_9_9_1 .LUT_INIT=16'b0000011100000100;
    LogicCell40 \U111_CYCLE_SM.TS_EN_LC_9_9_1  (
            .in0(N__4137),
            .in1(N__4131),
            .in2(N__4125),
            .in3(N__4110),
            .lcout(\U111_CYCLE_SM.TS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6384),
            .ce(),
            .sr(N__6336));
    defparam \U111_CYCLE_SM.TS_OUT_LC_9_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_OUT_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TS_OUT_LC_9_10_0 .LUT_INIT=16'b0111011101010111;
    LogicCell40 \U111_CYCLE_SM.TS_OUT_LC_9_10_0  (
            .in0(N__4646),
            .in1(N__4109),
            .in2(N__7438),
            .in3(N__5816),
            .lcout(TS_OUT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU111_CYCLE_SM.TS_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_9_10_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNO_0_LC_9_10_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNO_0_LC_9_10_7  (
            .in0(N__4973),
            .in1(N__5086),
            .in2(_gnd_net_),
            .in3(N__6413),
            .lcout(\U111_CYCLE_SM.N_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNINRNR_LC_9_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNINRNR_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNINRNR_LC_9_11_0 .LUT_INIT=16'b1010101011101010;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNINRNR_LC_9_11_0  (
            .in0(N__5784),
            .in1(N__7302),
            .in2(N__7088),
            .in3(N__7323),
            .lcout(U111_CYCLE_SM_OFFBOARD_EN_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_9_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_9_11_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_9_11_1  (
            .in0(N__6627),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7137),
            .lcout(\U111_CYCLE_SM.LATCH_EN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_9_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_9_11_2 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_9_11_2  (
            .in0(N__5384),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4566),
            .lcout(\U111_CYCLE_SM.N_106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_DELAY_RNIDR7G_LC_9_11_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_DELAY_RNIDR7G_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TS_DELAY_RNIDR7G_LC_9_11_3 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \U111_CYCLE_SM.TS_DELAY_RNIDR7G_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5817),
            .in3(N__7423),
            .lcout(\U111_CYCLE_SM.un4_TS_OUT_i_0 ),
            .ltout(\U111_CYCLE_SM.un4_TS_OUT_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI9UTM_0_LC_9_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI9UTM_0_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNI9UTM_0_LC_9_11_4 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNI9UTM_0_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4665),
            .in3(N__6626),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_9_11_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_2_LC_9_11_5 .LUT_INIT=16'b0000000010110000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_2_LC_9_11_5  (
            .in0(N__5093),
            .in1(N__4662),
            .in2(N__4656),
            .in3(N__4593),
            .lcout(\U111_CYCLE_SM.CYCLE_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6378),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_9_11_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_9_11_6 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_9_11_6  (
            .in0(N__5383),
            .in1(_gnd_net_),
            .in2(N__4537),
            .in3(N__4565),
            .lcout(\U111_CYCLE_SM.N_107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_0_2_LC_9_11_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_0_2_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_0_2_LC_9_11_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_0_2_LC_9_11_7  (
            .in0(N__4567),
            .in1(N__5382),
            .in2(_gnd_net_),
            .in3(N__4520),
            .lcout(\U111_CYCLE_SM.N_107_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_4_LC_9_12_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_4_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_4_LC_9_12_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_4_LC_9_12_0  (
            .in0(N__6593),
            .in1(N__5462),
            .in2(N__5451),
            .in3(N__7174),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6375),
            .ce(),
            .sr(N__6337));
    defparam \U111_CYCLE_SM.LATCH_EN_LC_9_12_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LATCH_EN_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LATCH_EN_LC_9_12_1 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \U111_CYCLE_SM.LATCH_EN_LC_9_12_1  (
            .in0(N__5133),
            .in1(N__5123),
            .in2(N__8363),
            .in3(N__6458),
            .lcout(\U111_CYCLE_SM.LATCH_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6375),
            .ce(),
            .sr(N__6337));
    defparam \U111_CYCLE_SM.UU_LATCHED_6_LC_9_12_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_6_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_6_LC_9_12_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_6_LC_9_12_2  (
            .in0(N__6595),
            .in1(N__5699),
            .in2(N__5688),
            .in3(N__7176),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6375),
            .ce(),
            .sr(N__6337));
    defparam \U111_CYCLE_SM.UM_LATCHED_7_LC_9_12_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_7_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_7_LC_9_12_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_7_LC_9_12_3  (
            .in0(N__7173),
            .in1(N__5045),
            .in2(N__5013),
            .in3(N__6592),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6375),
            .ce(),
            .sr(N__6337));
    defparam \U111_CYCLE_SM.TA_DIS_LC_9_12_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.TA_DIS_LC_9_12_4 .LUT_INIT=16'b0001000011111110;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_LC_9_12_4  (
            .in0(N__5124),
            .in1(N__5094),
            .in2(N__6130),
            .in3(N__5058),
            .lcout(\U111_CYCLE_SM.TA_DISZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6375),
            .ce(),
            .sr(N__6337));
    defparam \U111_CYCLE_SM.UM_LATCHED_3_LC_9_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_3_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_3_LC_9_12_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_3_LC_9_12_5  (
            .in0(N__7172),
            .in1(N__6026),
            .in2(N__6084),
            .in3(N__6591),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6375),
            .ce(),
            .sr(N__6337));
    defparam \U111_CYCLE_SM.UU_LATCHED_7_LC_9_12_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_7_LC_9_12_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_7_LC_9_12_6 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_7_LC_9_12_6  (
            .in0(N__6596),
            .in1(N__5541),
            .in2(N__5507),
            .in3(N__7177),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6375),
            .ce(),
            .sr(N__6337));
    defparam \U111_CYCLE_SM.UU_LATCHED_5_LC_9_12_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_5_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_5_LC_9_12_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_5_LC_9_12_7  (
            .in0(N__7175),
            .in1(N__5576),
            .in2(N__5625),
            .in3(N__6594),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6375),
            .ce(),
            .sr(N__6337));
    defparam \U111_CYCLE_SM.UM_LATCHED_RNIHDEL_7_LC_9_13_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNIHDEL_7_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNIHDEL_7_LC_9_13_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_RNIHDEL_7_LC_9_13_1  (
            .in0(N__8337),
            .in1(N__5044),
            .in2(_gnd_net_),
            .in3(N__5012),
            .lcout(un1_D_UM_AMIGA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_9_13_7.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_9_13_7.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_THRU_LUT4_0_LC_9_13_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_CLK40_THRU_LUT4_0_LC_9_13_7 (
            .in0(N__6390),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_CLK40_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIVRKT_6_LC_9_17_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIVRKT_6_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIVRKT_6_LC_9_17_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNIVRKT_6_LC_9_17_2  (
            .in0(N__5703),
            .in1(N__5668),
            .in2(_gnd_net_),
            .in3(N__8403),
            .lcout(N_124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNITPKT_5_LC_9_17_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNITPKT_5_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNITPKT_5_LC_9_17_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNITPKT_5_LC_9_17_5  (
            .in0(N__8402),
            .in1(N__5611),
            .in2(_gnd_net_),
            .in3(N__5580),
            .lcout(N_126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNI1UKT_7_LC_9_17_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNI1UKT_7_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNI1UKT_7_LC_9_17_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNI1UKT_7_LC_9_17_6  (
            .in0(N__5540),
            .in1(N__5508),
            .in2(_gnd_net_),
            .in3(N__8401),
            .lcout(N_123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIRNKT_4_LC_9_18_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIRNKT_4_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIRNKT_4_LC_9_18_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNIRNKT_4_LC_9_18_0  (
            .in0(N__5466),
            .in1(N__5440),
            .in2(_gnd_net_),
            .in3(N__8404),
            .lcout(N_127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_DIS_RNI576J_LC_9_18_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNI576J_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNI576J_LC_9_18_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNI576J_LC_9_18_1  (
            .in0(N__5388),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6137),
            .lcout(U111_CYCLE_SM_TEA_CPUn_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_9_18_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_9_18_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_9_18_3  (
            .in0(N__5298),
            .in1(N__5276),
            .in2(_gnd_net_),
            .in3(N__7903),
            .lcout(un1_D_UU_040_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_9_19_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_9_19_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_9_19_2  (
            .in0(N__5220),
            .in1(N__5198),
            .in2(_gnd_net_),
            .in3(N__7920),
            .lcout(un1_D_UM_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_RNI95EL_3_LC_9_19_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNI95EL_3_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNI95EL_3_LC_9_19_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_RNI95EL_3_LC_9_19_5  (
            .in0(N__6070),
            .in1(N__6033),
            .in2(_gnd_net_),
            .in3(N__8422),
            .lcout(un1_D_UM_AMIGA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_9_19_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_9_19_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_9_19_6  (
            .in0(N__6000),
            .in1(N__5958),
            .in2(_gnd_net_),
            .in3(N__7919),
            .lcout(un1_D_UM_040_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_10_6_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_10_6_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_10_6_3  (
            .in0(N__7902),
            .in1(N__8466),
            .in2(_gnd_net_),
            .in3(N__5919),
            .lcout(un2_D_LL_AMIGA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_10_6_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_10_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_10_6_6  (
            .in0(N__5877),
            .in1(N__7698),
            .in2(_gnd_net_),
            .in3(N__7901),
            .lcout(un2_D_LL_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TS_DELAY_LC_10_10_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TS_DELAY_LC_10_10_0 .SEQ_MODE=4'b1001;
    defparam \U111_CYCLE_SM.TS_DELAY_LC_10_10_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U111_CYCLE_SM.TS_DELAY_LC_10_10_0  (
            .in0(N__5838),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U111_CYCLE_SM.TS_DELAYZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6379),
            .ce(),
            .sr(N__6334));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_10_10_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_10_10_4 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_10_10_4  (
            .in0(N__7167),
            .in1(N__6635),
            .in2(N__7089),
            .in3(N__5802),
            .lcout(\U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6379),
            .ce(),
            .sr(N__6334));
    defparam \U111_CYCLE_SM.UM_LATCHED_2_LC_10_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_2_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_2_LC_10_11_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_2_LC_10_11_1  (
            .in0(N__6589),
            .in1(N__6674),
            .in2(N__6712),
            .in3(N__7139),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6376),
            .ce(),
            .sr(N__6338));
    defparam \U111_CYCLE_SM.UM_LATCHED_0_LC_10_11_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_0_LC_10_11_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_0_LC_10_11_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_0_LC_10_11_2  (
            .in0(N__7138),
            .in1(N__8555),
            .in2(N__8540),
            .in3(N__6588),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6376),
            .ce(),
            .sr(N__6338));
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_10_11_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_10_11_4 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_10_11_4 .LUT_INIT=16'b0010001000101110;
    LogicCell40 \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_10_11_4  (
            .in0(N__5783),
            .in1(N__6642),
            .in2(N__7087),
            .in3(N__5801),
            .lcout(\U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6376),
            .ce(),
            .sr(N__6338));
    defparam \U111_CYCLE_SM.CYCLE_EN_LC_10_11_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_EN_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.CYCLE_EN_LC_10_11_6 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \U111_CYCLE_SM.CYCLE_EN_LC_10_11_6  (
            .in0(N__7318),
            .in1(N__6641),
            .in2(_gnd_net_),
            .in3(N__6457),
            .lcout(\U111_CYCLE_SM.CYCLE_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6376),
            .ce(),
            .sr(N__6338));
    defparam \U111_CYCLE_SM.UM_LATCHED_6_LC_10_11_7 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_6_LC_10_11_7 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_6_LC_10_11_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_6_LC_10_11_7  (
            .in0(N__6590),
            .in1(N__8477),
            .in2(N__8465),
            .in3(N__7140),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6376),
            .ce(),
            .sr(N__6338));
    defparam \U111_CYCLE_SM.UU_LATCHED_1_LC_10_12_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_1_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_1_LC_10_12_1 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_1_LC_10_12_1  (
            .in0(N__6254),
            .in1(N__6604),
            .in2(N__6306),
            .in3(N__7171),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6374),
            .ce(),
            .sr(N__6339));
    defparam \U111_CYCLE_SM.UU_LATCHED_0_LC_10_12_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_0_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UU_LATCHED_0_LC_10_12_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_0_LC_10_12_2  (
            .in0(N__7170),
            .in1(N__6215),
            .in2(N__6200),
            .in3(N__6605),
            .lcout(\U111_CYCLE_SM.UU_LATCHEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6374),
            .ce(),
            .sr(N__6339));
    defparam \U111_CYCLE_SM.UM_LATCHED_5_LC_10_12_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_5_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.UM_LATCHED_5_LC_10_12_5 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_5_LC_10_12_5  (
            .in0(N__7646),
            .in1(N__6603),
            .in2(N__7694),
            .in3(N__7169),
            .lcout(\U111_CYCLE_SM.UM_LATCHEDZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6374),
            .ce(),
            .sr(N__6339));
    defparam \U111_CYCLE_SM.LW_TRANS_LC_10_12_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \U111_CYCLE_SM.LW_TRANS_LC_10_12_6 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \U111_CYCLE_SM.LW_TRANS_LC_10_12_6  (
            .in0(N__6533),
            .in1(N__6409),
            .in2(N__6497),
            .in3(N__6462),
            .lcout(\U111_CYCLE_SM.LW_TRANSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6374),
            .ce(),
            .sr(N__6339));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNILHKT_1_LC_10_18_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNILHKT_1_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNILHKT_1_LC_10_18_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNILHKT_1_LC_10_18_0  (
            .in0(N__8425),
            .in1(N__6292),
            .in2(_gnd_net_),
            .in3(N__6258),
            .lcout(N_130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIJFKT_0_LC_10_18_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIJFKT_0_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UU_LATCHED_RNIJFKT_0_LC_10_18_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UU_LATCHED_RNIJFKT_0_LC_10_18_1  (
            .in0(N__6219),
            .in1(N__6182),
            .in2(_gnd_net_),
            .in3(N__8424),
            .lcout(N_131),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_10_18_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_10_18_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_10_18_4  (
            .in0(N__6138),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7445),
            .lcout(N_66),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_RNID9EL_5_LC_10_19_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNID9EL_5_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNID9EL_5_LC_10_19_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_RNID9EL_5_LC_10_19_1  (
            .in0(N__7670),
            .in1(N__7653),
            .in2(_gnd_net_),
            .in3(N__8427),
            .lcout(un1_D_UM_AMIGA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_RNIB7EL_4_LC_10_19_3 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNIB7EL_4_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNIB7EL_4_LC_10_19_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_RNIB7EL_4_LC_10_19_3  (
            .in0(N__7611),
            .in1(N__7586),
            .in2(_gnd_net_),
            .in3(N__8426),
            .lcout(un1_D_UM_AMIGA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_10_19_4 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_10_19_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_10_19_4  (
            .in0(N__7918),
            .in1(N__7527),
            .in2(_gnd_net_),
            .in3(N__7493),
            .lcout(un1_D_UU_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LBENn_c_sbtinv_LC_11_1_1.C_ON=1'b0;
    defparam LBENn_c_sbtinv_LC_11_1_1.SEQ_MODE=4'b0000;
    defparam LBENn_c_sbtinv_LC_11_1_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 LBENn_c_sbtinv_LC_11_1_1 (
            .in0(N__7408),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(LBENn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_11_1_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_11_1_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_11_1_2  (
            .in0(N__7365),
            .in1(N__8544),
            .in2(_gnd_net_),
            .in3(N__7917),
            .lcout(un2_D_LL_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.CYCLE_EN_RNI26B3_LC_11_11_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.CYCLE_EN_RNI26B3_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.CYCLE_EN_RNI26B3_LC_11_11_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U111_CYCLE_SM.CYCLE_EN_RNI26B3_LC_11_11_0  (
            .in0(N__7319),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7301),
            .lcout(CPUBGn_c),
            .ltout(CPUBGn_c_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI8QUM_LC_11_11_1 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI8QUM_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI8QUM_LC_11_11_1 .LUT_INIT=16'b1010101011111010;
    LogicCell40 \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI8QUM_LC_11_11_1  (
            .in0(N__7168),
            .in1(_gnd_net_),
            .in2(N__7092),
            .in3(N__7068),
            .lcout(N_62_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_RNI73EL_2_LC_11_11_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNI73EL_2_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNI73EL_2_LC_11_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_RNI73EL_2_LC_11_11_5  (
            .in0(N__8396),
            .in1(N__6713),
            .in2(_gnd_net_),
            .in3(N__6675),
            .lcout(un1_D_UM_AMIGA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_RNI3VDL_0_LC_11_12_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNI3VDL_0_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNI3VDL_0_LC_11_12_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_RNI3VDL_0_LC_11_12_2  (
            .in0(N__8556),
            .in1(N__8519),
            .in2(_gnd_net_),
            .in3(N__8364),
            .lcout(un1_D_UM_AMIGA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.UM_LATCHED_RNIFBEL_6_LC_11_12_6 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNIFBEL_6_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.UM_LATCHED_RNIFBEL_6_LC_11_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.UM_LATCHED_RNIFBEL_6_LC_11_12_6  (
            .in0(N__8478),
            .in1(N__8452),
            .in2(_gnd_net_),
            .in3(N__8365),
            .lcout(N_125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_12_10_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_12_10_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_12_10_2  (
            .in0(N__7850),
            .in1(N__8279),
            .in2(_gnd_net_),
            .in3(N__8238),
            .lcout(un1_D_UM_040_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_10_7.C_ON=1'b0;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_10_7.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8205),
            .lcout(GB_BUFFER_CLK80_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_12_20_0 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_12_20_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_12_20_0  (
            .in0(N__7922),
            .in1(N__8160),
            .in2(_gnd_net_),
            .in3(N__8132),
            .lcout(un1_D_UU_040_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_12_20_2 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_12_20_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_12_20_2  (
            .in0(N__7923),
            .in1(N__8073),
            .in2(_gnd_net_),
            .in3(N__8048),
            .lcout(un1_D_UU_040_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_20_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_20_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_20_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_12_20_5 .C_ON=1'b0;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_12_20_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_12_20_5  (
            .in0(N__7976),
            .in1(N__7941),
            .in2(_gnd_net_),
            .in3(N__7921),
            .lcout(un1_D_UM_040_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U111_TOP

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 20 2025 20:31:24

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    TM,
    TT,
    A,
    CIACS1n,
    TICK50,
    RAMSPACEn,
    TICK60,
    CIACS0n,
    CLK6,
    CLK40_IN,
    CLK28_IN,
    REGSPACEn,
    CLK_CIA,
    BUFENn,
    TSn,
    RESETn,
    OVL,
    TACKn,
    ROMENn,
    PORTSIZE);

    input [1:0] TM;
    input [1:0] TT;
    input [31:1] A;
    output CIACS1n;
    output TICK50;
    output RAMSPACEn;
    output TICK60;
    output CIACS0n;
    input CLK6;
    input CLK40_IN;
    input CLK28_IN;
    output REGSPACEn;
    output CLK_CIA;
    output BUFENn;
    input TSn;
    input RESETn;
    input OVL;
    inout TACKn;
    output ROMENn;
    output PORTSIZE;

    wire N__7109;
    wire N__7108;
    wire N__7107;
    wire N__7099;
    wire N__7098;
    wire N__7097;
    wire N__7088;
    wire N__7087;
    wire N__7086;
    wire N__7079;
    wire N__7078;
    wire N__7077;
    wire N__7070;
    wire N__7069;
    wire N__7068;
    wire N__7061;
    wire N__7060;
    wire N__7059;
    wire N__7052;
    wire N__7051;
    wire N__7050;
    wire N__7043;
    wire N__7042;
    wire N__7041;
    wire N__7034;
    wire N__7033;
    wire N__7032;
    wire N__7025;
    wire N__7024;
    wire N__7023;
    wire N__7016;
    wire N__7015;
    wire N__7014;
    wire N__7007;
    wire N__7006;
    wire N__7005;
    wire N__6998;
    wire N__6997;
    wire N__6996;
    wire N__6989;
    wire N__6988;
    wire N__6987;
    wire N__6980;
    wire N__6979;
    wire N__6978;
    wire N__6971;
    wire N__6970;
    wire N__6969;
    wire N__6962;
    wire N__6961;
    wire N__6960;
    wire N__6953;
    wire N__6952;
    wire N__6951;
    wire N__6944;
    wire N__6943;
    wire N__6942;
    wire N__6935;
    wire N__6934;
    wire N__6933;
    wire N__6926;
    wire N__6925;
    wire N__6924;
    wire N__6917;
    wire N__6916;
    wire N__6915;
    wire N__6908;
    wire N__6907;
    wire N__6906;
    wire N__6899;
    wire N__6898;
    wire N__6897;
    wire N__6890;
    wire N__6889;
    wire N__6888;
    wire N__6881;
    wire N__6880;
    wire N__6879;
    wire N__6872;
    wire N__6871;
    wire N__6870;
    wire N__6863;
    wire N__6862;
    wire N__6861;
    wire N__6854;
    wire N__6853;
    wire N__6852;
    wire N__6845;
    wire N__6844;
    wire N__6843;
    wire N__6836;
    wire N__6835;
    wire N__6834;
    wire N__6827;
    wire N__6826;
    wire N__6825;
    wire N__6818;
    wire N__6817;
    wire N__6816;
    wire N__6809;
    wire N__6808;
    wire N__6807;
    wire N__6800;
    wire N__6799;
    wire N__6798;
    wire N__6791;
    wire N__6790;
    wire N__6789;
    wire N__6782;
    wire N__6781;
    wire N__6780;
    wire N__6773;
    wire N__6772;
    wire N__6771;
    wire N__6764;
    wire N__6763;
    wire N__6762;
    wire N__6745;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6733;
    wire N__6730;
    wire N__6727;
    wire N__6724;
    wire N__6721;
    wire N__6720;
    wire N__6717;
    wire N__6714;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6696;
    wire N__6693;
    wire N__6690;
    wire N__6685;
    wire N__6684;
    wire N__6683;
    wire N__6682;
    wire N__6681;
    wire N__6680;
    wire N__6679;
    wire N__6678;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6621;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6591;
    wire N__6588;
    wire N__6585;
    wire N__6580;
    wire N__6577;
    wire N__6576;
    wire N__6573;
    wire N__6570;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6558;
    wire N__6555;
    wire N__6552;
    wire N__6547;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6531;
    wire N__6528;
    wire N__6525;
    wire N__6520;
    wire N__6517;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6505;
    wire N__6502;
    wire N__6499;
    wire N__6496;
    wire N__6493;
    wire N__6490;
    wire N__6489;
    wire N__6486;
    wire N__6483;
    wire N__6478;
    wire N__6475;
    wire N__6474;
    wire N__6471;
    wire N__6468;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6439;
    wire N__6436;
    wire N__6435;
    wire N__6432;
    wire N__6429;
    wire N__6424;
    wire N__6421;
    wire N__6420;
    wire N__6417;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6403;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6391;
    wire N__6390;
    wire N__6389;
    wire N__6388;
    wire N__6387;
    wire N__6386;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6372;
    wire N__6365;
    wire N__6362;
    wire N__6355;
    wire N__6352;
    wire N__6351;
    wire N__6350;
    wire N__6349;
    wire N__6348;
    wire N__6347;
    wire N__6346;
    wire N__6343;
    wire N__6340;
    wire N__6337;
    wire N__6328;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6312;
    wire N__6311;
    wire N__6308;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6283;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6271;
    wire N__6270;
    wire N__6267;
    wire N__6264;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6252;
    wire N__6249;
    wire N__6246;
    wire N__6241;
    wire N__6240;
    wire N__6237;
    wire N__6234;
    wire N__6229;
    wire N__6228;
    wire N__6227;
    wire N__6226;
    wire N__6225;
    wire N__6224;
    wire N__6223;
    wire N__6222;
    wire N__6219;
    wire N__6212;
    wire N__6203;
    wire N__6200;
    wire N__6193;
    wire N__6192;
    wire N__6189;
    wire N__6188;
    wire N__6183;
    wire N__6180;
    wire N__6175;
    wire N__6174;
    wire N__6171;
    wire N__6170;
    wire N__6169;
    wire N__6166;
    wire N__6161;
    wire N__6158;
    wire N__6155;
    wire N__6148;
    wire N__6147;
    wire N__6144;
    wire N__6141;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6129;
    wire N__6126;
    wire N__6123;
    wire N__6118;
    wire N__6115;
    wire N__6112;
    wire N__6111;
    wire N__6108;
    wire N__6105;
    wire N__6100;
    wire N__6097;
    wire N__6096;
    wire N__6093;
    wire N__6090;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6075;
    wire N__6072;
    wire N__6069;
    wire N__6064;
    wire N__6063;
    wire N__6060;
    wire N__6057;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6042;
    wire N__6039;
    wire N__6036;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6010;
    wire N__6009;
    wire N__6008;
    wire N__6007;
    wire N__6006;
    wire N__6005;
    wire N__6004;
    wire N__6003;
    wire N__5998;
    wire N__5993;
    wire N__5984;
    wire N__5977;
    wire N__5976;
    wire N__5973;
    wire N__5972;
    wire N__5971;
    wire N__5970;
    wire N__5969;
    wire N__5968;
    wire N__5967;
    wire N__5964;
    wire N__5961;
    wire N__5958;
    wire N__5947;
    wire N__5938;
    wire N__5937;
    wire N__5936;
    wire N__5935;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5927;
    wire N__5926;
    wire N__5925;
    wire N__5920;
    wire N__5909;
    wire N__5906;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire N__5886;
    wire N__5883;
    wire N__5880;
    wire N__5875;
    wire N__5872;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5848;
    wire N__5845;
    wire N__5842;
    wire N__5839;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5827;
    wire N__5826;
    wire N__5823;
    wire N__5820;
    wire N__5815;
    wire N__5814;
    wire N__5811;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5794;
    wire N__5793;
    wire N__5790;
    wire N__5787;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5769;
    wire N__5768;
    wire N__5765;
    wire N__5760;
    wire N__5755;
    wire N__5752;
    wire N__5751;
    wire N__5750;
    wire N__5747;
    wire N__5742;
    wire N__5737;
    wire N__5734;
    wire N__5733;
    wire N__5732;
    wire N__5731;
    wire N__5730;
    wire N__5727;
    wire N__5724;
    wire N__5717;
    wire N__5710;
    wire N__5707;
    wire N__5706;
    wire N__5701;
    wire N__5698;
    wire N__5697;
    wire N__5696;
    wire N__5693;
    wire N__5688;
    wire N__5683;
    wire N__5680;
    wire N__5679;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5655;
    wire N__5652;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5635;
    wire N__5634;
    wire N__5633;
    wire N__5632;
    wire N__5631;
    wire N__5628;
    wire N__5627;
    wire N__5622;
    wire N__5619;
    wire N__5612;
    wire N__5605;
    wire N__5604;
    wire N__5603;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5565;
    wire N__5564;
    wire N__5563;
    wire N__5562;
    wire N__5559;
    wire N__5552;
    wire N__5549;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5476;
    wire N__5473;
    wire N__5472;
    wire N__5469;
    wire N__5466;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5440;
    wire N__5437;
    wire N__5434;
    wire N__5431;
    wire N__5428;
    wire N__5427;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5419;
    wire N__5416;
    wire N__5411;
    wire N__5406;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5394;
    wire N__5393;
    wire N__5392;
    wire N__5391;
    wire N__5388;
    wire N__5385;
    wire N__5378;
    wire N__5371;
    wire N__5368;
    wire N__5367;
    wire N__5366;
    wire N__5365;
    wire N__5364;
    wire N__5363;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5349;
    wire N__5348;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5334;
    wire N__5329;
    wire N__5326;
    wire N__5319;
    wire N__5316;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5302;
    wire N__5301;
    wire N__5298;
    wire N__5297;
    wire N__5290;
    wire N__5287;
    wire N__5282;
    wire N__5281;
    wire N__5280;
    wire N__5277;
    wire N__5274;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5244;
    wire N__5243;
    wire N__5240;
    wire N__5239;
    wire N__5238;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5230;
    wire N__5227;
    wire N__5224;
    wire N__5221;
    wire N__5218;
    wire N__5215;
    wire N__5212;
    wire N__5209;
    wire N__5204;
    wire N__5201;
    wire N__5196;
    wire N__5193;
    wire N__5188;
    wire N__5183;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5157;
    wire N__5154;
    wire N__5151;
    wire N__5150;
    wire N__5145;
    wire N__5142;
    wire N__5137;
    wire N__5134;
    wire N__5133;
    wire N__5132;
    wire N__5131;
    wire N__5130;
    wire N__5129;
    wire N__5124;
    wire N__5117;
    wire N__5114;
    wire N__5107;
    wire N__5106;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5098;
    wire N__5095;
    wire N__5094;
    wire N__5093;
    wire N__5092;
    wire N__5085;
    wire N__5078;
    wire N__5075;
    wire N__5068;
    wire N__5065;
    wire N__5064;
    wire N__5063;
    wire N__5062;
    wire N__5061;
    wire N__5060;
    wire N__5059;
    wire N__5056;
    wire N__5049;
    wire N__5044;
    wire N__5041;
    wire N__5032;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5020;
    wire N__5017;
    wire N__5014;
    wire N__5011;
    wire N__5008;
    wire N__5005;
    wire N__5002;
    wire N__4999;
    wire N__4996;
    wire N__4993;
    wire N__4990;
    wire N__4987;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4963;
    wire N__4960;
    wire N__4957;
    wire N__4954;
    wire N__4951;
    wire N__4948;
    wire N__4945;
    wire N__4942;
    wire N__4939;
    wire N__4936;
    wire N__4933;
    wire N__4930;
    wire N__4927;
    wire N__4926;
    wire N__4925;
    wire N__4922;
    wire N__4917;
    wire N__4912;
    wire N__4909;
    wire N__4908;
    wire N__4903;
    wire N__4900;
    wire N__4899;
    wire N__4898;
    wire N__4897;
    wire N__4894;
    wire N__4891;
    wire N__4884;
    wire N__4879;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4866;
    wire N__4861;
    wire N__4858;
    wire N__4857;
    wire N__4856;
    wire N__4853;
    wire N__4848;
    wire N__4843;
    wire N__4840;
    wire N__4837;
    wire N__4836;
    wire N__4835;
    wire N__4834;
    wire N__4833;
    wire N__4830;
    wire N__4821;
    wire N__4816;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4806;
    wire N__4805;
    wire N__4804;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4778;
    wire N__4775;
    wire N__4774;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4764;
    wire N__4761;
    wire N__4758;
    wire N__4755;
    wire N__4752;
    wire N__4749;
    wire N__4744;
    wire N__4737;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4723;
    wire N__4720;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4687;
    wire N__4686;
    wire N__4685;
    wire N__4682;
    wire N__4681;
    wire N__4680;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4664;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4650;
    wire N__4647;
    wire N__4644;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4618;
    wire N__4615;
    wire N__4612;
    wire N__4609;
    wire N__4606;
    wire N__4605;
    wire N__4604;
    wire N__4601;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4582;
    wire N__4575;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4558;
    wire N__4555;
    wire N__4552;
    wire N__4549;
    wire N__4546;
    wire N__4543;
    wire N__4542;
    wire N__4539;
    wire N__4536;
    wire N__4531;
    wire N__4530;
    wire N__4527;
    wire N__4524;
    wire N__4521;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4509;
    wire N__4508;
    wire N__4505;
    wire N__4504;
    wire N__4503;
    wire N__4502;
    wire N__4499;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4483;
    wire N__4478;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4459;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4447;
    wire N__4444;
    wire N__4443;
    wire N__4440;
    wire N__4439;
    wire N__4438;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4399;
    wire N__4396;
    wire N__4393;
    wire N__4392;
    wire N__4389;
    wire N__4388;
    wire N__4387;
    wire N__4384;
    wire N__4381;
    wire N__4376;
    wire N__4373;
    wire N__4372;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4354;
    wire N__4353;
    wire N__4352;
    wire N__4351;
    wire N__4348;
    wire N__4343;
    wire N__4338;
    wire N__4337;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4329;
    wire N__4328;
    wire N__4323;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4309;
    wire N__4308;
    wire N__4305;
    wire N__4300;
    wire N__4297;
    wire N__4294;
    wire N__4285;
    wire N__4282;
    wire N__4281;
    wire N__4280;
    wire N__4277;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4213;
    wire N__4212;
    wire N__4211;
    wire N__4210;
    wire N__4209;
    wire N__4206;
    wire N__4197;
    wire N__4192;
    wire N__4191;
    wire N__4190;
    wire N__4189;
    wire N__4188;
    wire N__4185;
    wire N__4176;
    wire N__4171;
    wire N__4170;
    wire N__4169;
    wire N__4166;
    wire N__4161;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4144;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4122;
    wire N__4117;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4107;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4095;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4078;
    wire N__4077;
    wire N__4076;
    wire N__4075;
    wire N__4072;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4045;
    wire N__4042;
    wire N__4039;
    wire N__4038;
    wire N__4037;
    wire N__4036;
    wire N__4035;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4025;
    wire N__4022;
    wire N__4017;
    wire N__4006;
    wire N__4003;
    wire N__4000;
    wire N__3997;
    wire N__3994;
    wire N__3991;
    wire N__3988;
    wire N__3985;
    wire N__3982;
    wire N__3979;
    wire N__3978;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3961;
    wire N__3960;
    wire N__3959;
    wire N__3958;
    wire N__3955;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3940;
    wire N__3931;
    wire N__3928;
    wire N__3927;
    wire N__3926;
    wire N__3925;
    wire N__3924;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3910;
    wire N__3901;
    wire N__3900;
    wire N__3899;
    wire N__3896;
    wire N__3895;
    wire N__3894;
    wire N__3893;
    wire N__3892;
    wire N__3891;
    wire N__3888;
    wire N__3885;
    wire N__3882;
    wire N__3879;
    wire N__3876;
    wire N__3869;
    wire N__3856;
    wire N__3853;
    wire N__3852;
    wire N__3851;
    wire N__3850;
    wire N__3847;
    wire N__3846;
    wire N__3843;
    wire N__3838;
    wire N__3835;
    wire N__3830;
    wire N__3823;
    wire N__3820;
    wire N__3817;
    wire N__3814;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3802;
    wire N__3799;
    wire N__3796;
    wire N__3795;
    wire N__3792;
    wire N__3791;
    wire N__3790;
    wire N__3787;
    wire N__3786;
    wire N__3781;
    wire N__3778;
    wire N__3775;
    wire N__3772;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3760;
    wire N__3757;
    wire N__3754;
    wire N__3749;
    wire N__3746;
    wire N__3743;
    wire N__3736;
    wire N__3733;
    wire N__3730;
    wire N__3727;
    wire N__3726;
    wire N__3723;
    wire N__3720;
    wire N__3715;
    wire N__3712;
    wire N__3709;
    wire N__3706;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3694;
    wire N__3691;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3679;
    wire N__3678;
    wire N__3675;
    wire N__3672;
    wire N__3667;
    wire N__3664;
    wire N__3661;
    wire N__3658;
    wire N__3655;
    wire N__3652;
    wire N__3649;
    wire N__3646;
    wire N__3643;
    wire N__3642;
    wire N__3641;
    wire N__3638;
    wire N__3633;
    wire N__3628;
    wire N__3627;
    wire N__3624;
    wire N__3621;
    wire N__3618;
    wire N__3613;
    wire N__3610;
    wire N__3607;
    wire N__3606;
    wire N__3605;
    wire N__3604;
    wire N__3603;
    wire N__3600;
    wire N__3597;
    wire N__3594;
    wire N__3591;
    wire N__3588;
    wire N__3577;
    wire N__3576;
    wire N__3575;
    wire N__3572;
    wire N__3571;
    wire N__3568;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3550;
    wire N__3547;
    wire N__3544;
    wire N__3541;
    wire N__3538;
    wire N__3537;
    wire N__3534;
    wire N__3531;
    wire N__3526;
    wire N__3525;
    wire N__3522;
    wire N__3519;
    wire N__3516;
    wire N__3511;
    wire N__3508;
    wire N__3505;
    wire N__3504;
    wire N__3503;
    wire N__3502;
    wire N__3497;
    wire N__3494;
    wire N__3493;
    wire N__3490;
    wire N__3487;
    wire N__3484;
    wire N__3479;
    wire N__3476;
    wire N__3475;
    wire N__3474;
    wire N__3471;
    wire N__3468;
    wire N__3465;
    wire N__3460;
    wire N__3455;
    wire N__3452;
    wire N__3449;
    wire N__3446;
    wire N__3443;
    wire N__3440;
    wire N__3437;
    wire N__3432;
    wire N__3429;
    wire N__3424;
    wire N__3421;
    wire N__3418;
    wire N__3417;
    wire N__3414;
    wire N__3411;
    wire N__3408;
    wire N__3405;
    wire N__3400;
    wire N__3397;
    wire N__3394;
    wire N__3391;
    wire N__3388;
    wire N__3385;
    wire N__3382;
    wire N__3379;
    wire N__3376;
    wire N__3373;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3361;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3345;
    wire N__3344;
    wire N__3339;
    wire N__3336;
    wire N__3331;
    wire N__3328;
    wire N__3325;
    wire N__3322;
    wire N__3321;
    wire N__3316;
    wire N__3315;
    wire N__3312;
    wire N__3309;
    wire N__3304;
    wire N__3301;
    wire N__3298;
    wire N__3295;
    wire N__3292;
    wire N__3289;
    wire N__3286;
    wire N__3283;
    wire N__3280;
    wire N__3277;
    wire N__3274;
    wire N__3271;
    wire N__3268;
    wire N__3265;
    wire N__3262;
    wire N__3259;
    wire N__3256;
    wire N__3253;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3241;
    wire N__3240;
    wire N__3235;
    wire N__3234;
    wire N__3231;
    wire N__3228;
    wire N__3225;
    wire N__3222;
    wire N__3217;
    wire N__3214;
    wire N__3213;
    wire N__3212;
    wire N__3209;
    wire N__3206;
    wire N__3203;
    wire N__3202;
    wire N__3199;
    wire N__3194;
    wire N__3191;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3177;
    wire N__3172;
    wire N__3169;
    wire N__3166;
    wire N__3165;
    wire N__3162;
    wire N__3161;
    wire N__3158;
    wire N__3155;
    wire N__3152;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3123;
    wire N__3120;
    wire N__3117;
    wire N__3112;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3099;
    wire N__3094;
    wire N__3093;
    wire N__3090;
    wire N__3087;
    wire N__3082;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3070;
    wire N__3069;
    wire N__3064;
    wire N__3061;
    wire N__3058;
    wire N__3055;
    wire N__3052;
    wire N__3049;
    wire N__3046;
    wire N__3043;
    wire N__3040;
    wire N__3037;
    wire N__3036;
    wire N__3033;
    wire N__3030;
    wire N__3025;
    wire N__3024;
    wire N__3021;
    wire N__3018;
    wire N__3015;
    wire N__3010;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__2998;
    wire N__2997;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2982;
    wire N__2979;
    wire N__2974;
    wire N__2971;
    wire N__2968;
    wire N__2965;
    wire N__2964;
    wire N__2961;
    wire N__2958;
    wire N__2953;
    wire N__2950;
    wire N__2947;
    wire N__2944;
    wire N__2943;
    wire N__2940;
    wire N__2937;
    wire N__2934;
    wire N__2931;
    wire N__2926;
    wire N__2923;
    wire N__2920;
    wire N__2917;
    wire N__2914;
    wire N__2913;
    wire N__2910;
    wire N__2907;
    wire N__2902;
    wire N__2899;
    wire N__2896;
    wire N__2893;
    wire N__2890;
    wire N__2887;
    wire N__2884;
    wire N__2883;
    wire N__2880;
    wire N__2877;
    wire N__2872;
    wire N__2869;
    wire N__2866;
    wire N__2863;
    wire N__2860;
    wire N__2859;
    wire N__2854;
    wire N__2851;
    wire N__2848;
    wire N__2845;
    wire N__2842;
    wire N__2839;
    wire N__2838;
    wire N__2833;
    wire N__2830;
    wire N__2827;
    wire N__2824;
    wire N__2821;
    wire N__2820;
    wire N__2817;
    wire N__2814;
    wire N__2811;
    wire N__2806;
    wire N__2803;
    wire N__2800;
    wire N__2797;
    wire N__2794;
    wire N__2793;
    wire N__2790;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2776;
    wire N__2773;
    wire N__2770;
    wire N__2767;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2755;
    wire N__2752;
    wire N__2749;
    wire N__2746;
    wire N__2743;
    wire N__2740;
    wire N__2737;
    wire N__2734;
    wire N__2731;
    wire N__2728;
    wire N__2725;
    wire N__2724;
    wire N__2723;
    wire N__2722;
    wire N__2721;
    wire N__2720;
    wire N__2719;
    wire N__2718;
    wire N__2717;
    wire N__2716;
    wire N__2715;
    wire N__2714;
    wire N__2713;
    wire N__2712;
    wire N__2711;
    wire N__2710;
    wire N__2677;
    wire CLK80_OUT;
    wire GNDG0;
    wire VCCG0;
    wire A_c_16;
    wire A_c_17;
    wire A_c_31;
    wire A_c_24;
    wire A_c_25;
    wire \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_3 ;
    wire A_c_30;
    wire A_c_28;
    wire A_c_29;
    wire A_c_27;
    wire \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4 ;
    wire A_c_20;
    wire \U409_TRANSFER_ACK.N_41_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3Z0Z_2 ;
    wire U409_CIA_PORTSIZE_i_a2_0_3;
    wire A_c_19;
    wire A_c_18;
    wire TT_c_0;
    wire A_c_26;
    wire TT_c_1;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_11_cascade_ ;
    wire \U409_TRANSFER_ACK.N_17 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_4 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_11 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_14 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_10 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_17 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_16 ;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ;
    wire TM_c_0;
    wire TM_c_1;
    wire PORTSIZE_i_a2;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_12 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ;
    wire \U409_CIA.N_89 ;
    wire A_c_22;
    wire OVL_c;
    wire \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3Z0Z_4_cascade_ ;
    wire N_53_i;
    wire \U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ;
    wire \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ;
    wire TACK_OUTn;
    wire \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.N_54_4_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_5_cascade_ ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a3_0_1_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a3_0_1_0_cascade_ ;
    wire \U409_TRANSFER_ACK.N_54_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0Z0Z_0 ;
    wire A_c_23;
    wire \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3Z0Z_4 ;
    wire \U409_ADDRESS_DECODE.N_16_i ;
    wire un1_RAMSPACEn_i_i_a3_cascade_;
    wire N_11_i;
    wire un1_RAMSPACEn_i_i_a3;
    wire TACKn_in;
    wire un1_REGSPACEn_i_i_a3_0_a2_cascade_;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire N_90;
    wire A_c_21;
    wire N_80;
    wire N_52_i;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6 ;
    wire \INVU409_TRANSFER_ACK.TACK_EN_iC_net ;
    wire \U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en ;
    wire ROMENn_c;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.ROMENnC_net ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_0 ;
    wire TSn_c;
    wire N_76;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_EN_e_1 ;
    wire \U409_TRANSFER_ACK.N_28_4 ;
    wire \U409_TRANSFER_ACK.N_28_3 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.N_64 ;
    wire \U409_TRANSFER_ACK.N_63_cascade_ ;
    wire \U409_TRANSFER_ACK.m9_i_1_cascade_ ;
    wire \U409_TRANSFER_ACK.N_45 ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire \U409_TRANSFER_ACK.N_73 ;
    wire \U409_TRANSFER_ACK.N_60 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_ ;
    wire \U409_TRANSFER_ACK.N_65 ;
    wire CLK40_IN_c;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_68 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_23 ;
    wire CONSTANT_ONE_NET;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_CIACS1n_i;
    wire CIA_ENABLE;
    wire CIA_ENABLE_cascade_;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_CIACS0n_i;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_1C_net ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_0C_net ;
    wire RESETn_c;
    wire RESETn_c_i;
    wire \U409_CIA.N_93_cascade_ ;
    wire \U409_CIA.VMA_RNOZ0Z_1_cascade_ ;
    wire \U409_CIA.VMA_3_0_a2_2 ;
    wire \U409_CIA.VMAZ0 ;
    wire \U409_CIA.N_91_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a2_2 ;
    wire \U409_CIA.N_91 ;
    wire \U409_CIA.un1_CIA_CLK_COUNT_2_1 ;
    wire \U409_CIA.CLK_CIA_r_1_cascade_ ;
    wire \U409_CIA.CLK_CIA6_1_0 ;
    wire CLK_CIA_c;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire TICK50_c;
    wire bfn_13_2_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire bfn_13_3_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire \U409_CIA.CLK_CIA6_1 ;
    wire bfn_13_12_0_;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.CIA_CLK_COUNT11 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_6 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_5 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_6 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_7 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire CLK28_IN_c_g;
    wire \U409_TICK.TICK503_11 ;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.TICK603_11 ;
    wire \U409_TICK.TICK603_8_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_9 ;
    wire TICK60_c;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire bfn_15_1_0_;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire bfn_15_2_0_;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire CLK6_c_g;
    wire TACK_EN_i;
    wire N_525_i;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__4804),
            .RESETB(N__5026),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__7107),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__7109),
            .DIN(N__7108),
            .DOUT(N__7107),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__7109),
            .PADOUT(N__7108),
            .PADIN(N__7107),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__7097),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__7099),
            .DIN(N__7098),
            .DOUT(N__7097),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__7099),
            .PADOUT(N__7098),
            .PADIN(N__7097),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__7088),
            .DIN(N__7087),
            .DOUT(N__7086),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__7088),
            .PADOUT(N__7087),
            .PADIN(N__7086),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__7079),
            .DIN(N__7078),
            .DOUT(N__7077),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__7079),
            .PADOUT(N__7078),
            .PADIN(N__7077),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__7070),
            .DIN(N__7069),
            .DOUT(N__7068),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__7070),
            .PADOUT(N__7069),
            .PADIN(N__7068),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS1n_obuf_iopad (
            .OE(N__7061),
            .DIN(N__7060),
            .DOUT(N__7059),
            .PACKAGEPIN(CIACS1n));
    defparam CIACS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS1n_obuf_preio (
            .PADOEN(N__7061),
            .PADOUT(N__7060),
            .PADIN(N__7059),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4993),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_obuf_iopad (
            .OE(N__7052),
            .DIN(N__7051),
            .DOUT(N__7050),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGSPACEn_obuf_preio (
            .PADOEN(N__7052),
            .PADOUT(N__7051),
            .PADIN(N__7050),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4249),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_1_iopad (
            .OE(N__7043),
            .DIN(N__7042),
            .DOUT(N__7041),
            .PACKAGEPIN(TM[1]));
    defparam TM_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_1_preio (
            .PADOEN(N__7043),
            .PADOUT(N__7042),
            .PADIN(N__7041),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__7034),
            .DIN(N__7033),
            .DOUT(N__7032),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__7034),
            .PADOUT(N__7033),
            .PADIN(N__7032),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_CIA_obuf_iopad (
            .OE(N__7025),
            .DIN(N__7024),
            .DOUT(N__7023),
            .PACKAGEPIN(CLK_CIA));
    defparam CLK_CIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_CIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_CIA_obuf_preio (
            .PADOEN(N__7025),
            .PADOUT(N__7024),
            .PADIN(N__7023),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5440),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__7016),
            .DIN(N__7015),
            .DOUT(N__7014),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__7016),
            .PADOUT(N__7015),
            .PADIN(N__7014),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_obuf_iopad (
            .OE(N__7007),
            .DIN(N__7006),
            .DOUT(N__7005),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMSPACEn_obuf_preio (
            .PADOEN(N__7007),
            .PADOUT(N__7006),
            .PADIN(N__7005),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3388),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__6998),
            .DIN(N__6997),
            .DOUT(N__6996),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__6998),
            .PADOUT(N__6997),
            .PADIN(N__6996),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6643),
            .DIN0(TACKn_in),
            .DOUT0(N__3661),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__6989),
            .DIN(N__6988),
            .DOUT(N__6987),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__6989),
            .PADOUT(N__6988),
            .PADIN(N__6987),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ROMENn_obuf_iopad (
            .OE(N__6980),
            .DIN(N__6979),
            .DOUT(N__6978),
            .PACKAGEPIN(ROMENn));
    defparam ROMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ROMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ROMENn_obuf_preio (
            .PADOEN(N__6980),
            .PADOUT(N__6979),
            .PADIN(N__6978),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4150),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__6971),
            .DIN(N__6970),
            .DOUT(N__6969),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__6971),
            .PADOUT(N__6970),
            .PADIN(N__6969),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__6962),
            .DIN(N__6961),
            .DOUT(N__6960),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__6962),
            .PADOUT(N__6961),
            .PADIN(N__6960),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__6953),
            .DIN(N__6952),
            .DOUT(N__6951),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__6953),
            .PADOUT(N__6952),
            .PADIN(N__6951),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3712),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__6944),
            .DIN(N__6943),
            .DOUT(N__6942),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__6944),
            .PADOUT(N__6943),
            .PADIN(N__6942),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3295),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__6935),
            .DIN(N__6934),
            .DOUT(N__6933),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__6935),
            .PADOUT(N__6934),
            .PADIN(N__6933),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__6926),
            .DIN(N__6925),
            .DOUT(N__6924),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__6926),
            .PADOUT(N__6925),
            .PADIN(N__6924),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__6917),
            .DIN(N__6916),
            .DOUT(N__6915),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__6917),
            .PADOUT(N__6916),
            .PADIN(N__6915),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__6908),
            .DIN(N__6907),
            .DOUT(N__6906),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__6908),
            .PADOUT(N__6907),
            .PADIN(N__6906),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__6899),
            .DIN(N__6898),
            .DOUT(N__6897),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__6899),
            .PADOUT(N__6898),
            .PADIN(N__6897),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__6890),
            .DIN(N__6889),
            .DOUT(N__6888),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__6890),
            .PADOUT(N__6889),
            .PADIN(N__6888),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_0_iopad (
            .OE(N__6881),
            .DIN(N__6880),
            .DOUT(N__6879),
            .PACKAGEPIN(TM[0]));
    defparam TM_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_0_preio (
            .PADOEN(N__6881),
            .PADOUT(N__6880),
            .PADIN(N__6879),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__6872),
            .DIN(N__6871),
            .DOUT(N__6870),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__6872),
            .PADOUT(N__6871),
            .PADIN(N__6870),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__6863),
            .DIN(N__6862),
            .DOUT(N__6861),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__6863),
            .PADOUT(N__6862),
            .PADIN(N__6861),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__6854),
            .DIN(N__6853),
            .DOUT(N__6852),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__6854),
            .PADOUT(N__6853),
            .PADIN(N__6852),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS0n_obuf_iopad (
            .OE(N__6845),
            .DIN(N__6844),
            .DOUT(N__6843),
            .PACKAGEPIN(CIACS0n));
    defparam CIACS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS0n_obuf_preio (
            .PADOEN(N__6845),
            .PADOUT(N__6844),
            .PADIN(N__6843),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4948),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__6836),
            .DIN(N__6835),
            .DOUT(N__6834),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__6836),
            .PADOUT(N__6835),
            .PADIN(N__6834),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5533),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__6827),
            .DIN(N__6826),
            .DOUT(N__6825),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__6827),
            .PADOUT(N__6826),
            .PADIN(N__6825),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__6818),
            .DIN(N__6817),
            .DOUT(N__6816),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__6818),
            .PADOUT(N__6817),
            .PADIN(N__6816),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__6809),
            .DIN(N__6808),
            .DOUT(N__6807),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__6809),
            .PADOUT(N__6808),
            .PADIN(N__6807),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__6800),
            .DIN(N__6799),
            .DOUT(N__6798),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__6800),
            .PADOUT(N__6799),
            .PADIN(N__6798),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__6791),
            .DIN(N__6790),
            .DOUT(N__6789),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__6791),
            .PADOUT(N__6790),
            .PADIN(N__6789),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__6782),
            .DIN(N__6781),
            .DOUT(N__6780),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__6782),
            .PADOUT(N__6781),
            .PADIN(N__6780),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5899),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__6773),
            .DIN(N__6772),
            .DOUT(N__6771),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__6773),
            .PADOUT(N__6772),
            .PADIN(N__6771),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__6764),
            .DIN(N__6763),
            .DOUT(N__6762),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__6764),
            .PADOUT(N__6763),
            .PADIN(N__6762),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1592 (
            .O(N__6745),
            .I(N__6741));
    InMux I__1591 (
            .O(N__6744),
            .I(N__6738));
    LocalMux I__1590 (
            .O(N__6741),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__1589 (
            .O(N__6738),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    CascadeMux I__1588 (
            .O(N__6733),
            .I(N__6730));
    InMux I__1587 (
            .O(N__6730),
            .I(N__6727));
    LocalMux I__1586 (
            .O(N__6727),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__1585 (
            .O(N__6724),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__1584 (
            .O(N__6721),
            .I(N__6717));
    InMux I__1583 (
            .O(N__6720),
            .I(N__6714));
    LocalMux I__1582 (
            .O(N__6717),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__1581 (
            .O(N__6714),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    InMux I__1580 (
            .O(N__6709),
            .I(N__6706));
    LocalMux I__1579 (
            .O(N__6706),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__1578 (
            .O(N__6703),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__1577 (
            .O(N__6700),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__1576 (
            .O(N__6697),
            .I(N__6693));
    InMux I__1575 (
            .O(N__6696),
            .I(N__6690));
    LocalMux I__1574 (
            .O(N__6693),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__1573 (
            .O(N__6690),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    ClkMux I__1572 (
            .O(N__6685),
            .I(N__6661));
    ClkMux I__1571 (
            .O(N__6684),
            .I(N__6661));
    ClkMux I__1570 (
            .O(N__6683),
            .I(N__6661));
    ClkMux I__1569 (
            .O(N__6682),
            .I(N__6661));
    ClkMux I__1568 (
            .O(N__6681),
            .I(N__6661));
    ClkMux I__1567 (
            .O(N__6680),
            .I(N__6661));
    ClkMux I__1566 (
            .O(N__6679),
            .I(N__6661));
    ClkMux I__1565 (
            .O(N__6678),
            .I(N__6661));
    GlobalMux I__1564 (
            .O(N__6661),
            .I(N__6658));
    gio2CtrlBuf I__1563 (
            .O(N__6658),
            .I(CLK6_c_g));
    InMux I__1562 (
            .O(N__6655),
            .I(N__6652));
    LocalMux I__1561 (
            .O(N__6652),
            .I(N__6649));
    Span12Mux_v I__1560 (
            .O(N__6649),
            .I(N__6646));
    Odrv12 I__1559 (
            .O(N__6646),
            .I(TACK_EN_i));
    IoInMux I__1558 (
            .O(N__6643),
            .I(N__6640));
    LocalMux I__1557 (
            .O(N__6640),
            .I(N__6637));
    IoSpan4Mux I__1556 (
            .O(N__6637),
            .I(N__6634));
    Span4Mux_s3_v I__1555 (
            .O(N__6634),
            .I(N__6631));
    Span4Mux_v I__1554 (
            .O(N__6631),
            .I(N__6628));
    Span4Mux_v I__1553 (
            .O(N__6628),
            .I(N__6625));
    Odrv4 I__1552 (
            .O(N__6625),
            .I(N_525_i));
    CascadeMux I__1551 (
            .O(N__6622),
            .I(N__6618));
    InMux I__1550 (
            .O(N__6621),
            .I(N__6615));
    InMux I__1549 (
            .O(N__6618),
            .I(N__6612));
    LocalMux I__1548 (
            .O(N__6615),
            .I(N__6609));
    LocalMux I__1547 (
            .O(N__6612),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    Odrv4 I__1546 (
            .O(N__6609),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    InMux I__1545 (
            .O(N__6604),
            .I(N__6601));
    LocalMux I__1544 (
            .O(N__6601),
            .I(N__6598));
    Odrv4 I__1543 (
            .O(N__6598),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__1542 (
            .O(N__6595),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__1541 (
            .O(N__6592),
            .I(N__6588));
    InMux I__1540 (
            .O(N__6591),
            .I(N__6585));
    LocalMux I__1539 (
            .O(N__6588),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__1538 (
            .O(N__6585),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    InMux I__1537 (
            .O(N__6580),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__1536 (
            .O(N__6577),
            .I(N__6573));
    InMux I__1535 (
            .O(N__6576),
            .I(N__6570));
    LocalMux I__1534 (
            .O(N__6573),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__1533 (
            .O(N__6570),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__1532 (
            .O(N__6565),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__1531 (
            .O(N__6562),
            .I(N__6559));
    LocalMux I__1530 (
            .O(N__6559),
            .I(N__6555));
    InMux I__1529 (
            .O(N__6558),
            .I(N__6552));
    Odrv4 I__1528 (
            .O(N__6555),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__1527 (
            .O(N__6552),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    InMux I__1526 (
            .O(N__6547),
            .I(N__6544));
    LocalMux I__1525 (
            .O(N__6544),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__1524 (
            .O(N__6541),
            .I(bfn_15_2_0_));
    InMux I__1523 (
            .O(N__6538),
            .I(N__6535));
    LocalMux I__1522 (
            .O(N__6535),
            .I(N__6532));
    Span4Mux_v I__1521 (
            .O(N__6532),
            .I(N__6528));
    InMux I__1520 (
            .O(N__6531),
            .I(N__6525));
    Odrv4 I__1519 (
            .O(N__6528),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__1518 (
            .O(N__6525),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    InMux I__1517 (
            .O(N__6520),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__1516 (
            .O(N__6517),
            .I(N__6513));
    InMux I__1515 (
            .O(N__6516),
            .I(N__6510));
    LocalMux I__1514 (
            .O(N__6513),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__1513 (
            .O(N__6510),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__1512 (
            .O(N__6505),
            .I(N__6502));
    LocalMux I__1511 (
            .O(N__6502),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__1510 (
            .O(N__6499),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__1509 (
            .O(N__6496),
            .I(N__6493));
    LocalMux I__1508 (
            .O(N__6493),
            .I(N__6490));
    Span4Mux_h I__1507 (
            .O(N__6490),
            .I(N__6486));
    InMux I__1506 (
            .O(N__6489),
            .I(N__6483));
    Odrv4 I__1505 (
            .O(N__6486),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__1504 (
            .O(N__6483),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    InMux I__1503 (
            .O(N__6478),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__1502 (
            .O(N__6475),
            .I(N__6471));
    InMux I__1501 (
            .O(N__6474),
            .I(N__6468));
    LocalMux I__1500 (
            .O(N__6471),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__1499 (
            .O(N__6468),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    CascadeMux I__1498 (
            .O(N__6463),
            .I(N__6460));
    InMux I__1497 (
            .O(N__6460),
            .I(N__6457));
    LocalMux I__1496 (
            .O(N__6457),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__1495 (
            .O(N__6454),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__1494 (
            .O(N__6451),
            .I(N__6447));
    InMux I__1493 (
            .O(N__6450),
            .I(N__6444));
    LocalMux I__1492 (
            .O(N__6447),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__1491 (
            .O(N__6444),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    InMux I__1490 (
            .O(N__6439),
            .I(N__6436));
    LocalMux I__1489 (
            .O(N__6436),
            .I(N__6432));
    InMux I__1488 (
            .O(N__6435),
            .I(N__6429));
    Odrv4 I__1487 (
            .O(N__6432),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__1486 (
            .O(N__6429),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    CascadeMux I__1485 (
            .O(N__6424),
            .I(N__6421));
    InMux I__1484 (
            .O(N__6421),
            .I(N__6417));
    CascadeMux I__1483 (
            .O(N__6420),
            .I(N__6414));
    LocalMux I__1482 (
            .O(N__6417),
            .I(N__6411));
    InMux I__1481 (
            .O(N__6414),
            .I(N__6408));
    Odrv4 I__1480 (
            .O(N__6411),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__1479 (
            .O(N__6408),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    InMux I__1478 (
            .O(N__6403),
            .I(N__6399));
    InMux I__1477 (
            .O(N__6402),
            .I(N__6396));
    LocalMux I__1476 (
            .O(N__6399),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__1475 (
            .O(N__6396),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    CascadeMux I__1474 (
            .O(N__6391),
            .I(N__6382));
    InMux I__1473 (
            .O(N__6390),
            .I(N__6379));
    InMux I__1472 (
            .O(N__6389),
            .I(N__6372));
    InMux I__1471 (
            .O(N__6388),
            .I(N__6372));
    InMux I__1470 (
            .O(N__6387),
            .I(N__6372));
    InMux I__1469 (
            .O(N__6386),
            .I(N__6365));
    InMux I__1468 (
            .O(N__6385),
            .I(N__6365));
    InMux I__1467 (
            .O(N__6382),
            .I(N__6365));
    LocalMux I__1466 (
            .O(N__6379),
            .I(N__6362));
    LocalMux I__1465 (
            .O(N__6372),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__1464 (
            .O(N__6365),
            .I(\U409_TICK.TICK603_9 ));
    Odrv4 I__1463 (
            .O(N__6362),
            .I(\U409_TICK.TICK603_9 ));
    CascadeMux I__1462 (
            .O(N__6355),
            .I(N__6352));
    InMux I__1461 (
            .O(N__6352),
            .I(N__6343));
    InMux I__1460 (
            .O(N__6351),
            .I(N__6340));
    InMux I__1459 (
            .O(N__6350),
            .I(N__6337));
    InMux I__1458 (
            .O(N__6349),
            .I(N__6328));
    InMux I__1457 (
            .O(N__6348),
            .I(N__6328));
    InMux I__1456 (
            .O(N__6347),
            .I(N__6328));
    InMux I__1455 (
            .O(N__6346),
            .I(N__6328));
    LocalMux I__1454 (
            .O(N__6343),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__1453 (
            .O(N__6340),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__1452 (
            .O(N__6337),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__1451 (
            .O(N__6328),
            .I(\U409_TICK.TICK603_14 ));
    CascadeMux I__1450 (
            .O(N__6319),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    InMux I__1449 (
            .O(N__6316),
            .I(N__6313));
    LocalMux I__1448 (
            .O(N__6313),
            .I(N__6308));
    CascadeMux I__1447 (
            .O(N__6312),
            .I(N__6304));
    InMux I__1446 (
            .O(N__6311),
            .I(N__6301));
    Span4Mux_h I__1445 (
            .O(N__6308),
            .I(N__6298));
    InMux I__1444 (
            .O(N__6307),
            .I(N__6295));
    InMux I__1443 (
            .O(N__6304),
            .I(N__6292));
    LocalMux I__1442 (
            .O(N__6301),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    Odrv4 I__1441 (
            .O(N__6298),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__1440 (
            .O(N__6295),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__1439 (
            .O(N__6292),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__1438 (
            .O(N__6283),
            .I(N__6279));
    InMux I__1437 (
            .O(N__6282),
            .I(N__6276));
    LocalMux I__1436 (
            .O(N__6279),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__1435 (
            .O(N__6276),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__1434 (
            .O(N__6271),
            .I(N__6267));
    InMux I__1433 (
            .O(N__6270),
            .I(N__6264));
    LocalMux I__1432 (
            .O(N__6267),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__1431 (
            .O(N__6264),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    CascadeMux I__1430 (
            .O(N__6259),
            .I(N__6256));
    InMux I__1429 (
            .O(N__6256),
            .I(N__6253));
    LocalMux I__1428 (
            .O(N__6253),
            .I(N__6249));
    InMux I__1427 (
            .O(N__6252),
            .I(N__6246));
    Odrv4 I__1426 (
            .O(N__6249),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__1425 (
            .O(N__6246),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__1424 (
            .O(N__6241),
            .I(N__6237));
    InMux I__1423 (
            .O(N__6240),
            .I(N__6234));
    LocalMux I__1422 (
            .O(N__6237),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__1421 (
            .O(N__6234),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__1420 (
            .O(N__6229),
            .I(N__6219));
    InMux I__1419 (
            .O(N__6228),
            .I(N__6212));
    InMux I__1418 (
            .O(N__6227),
            .I(N__6212));
    InMux I__1417 (
            .O(N__6226),
            .I(N__6212));
    InMux I__1416 (
            .O(N__6225),
            .I(N__6203));
    InMux I__1415 (
            .O(N__6224),
            .I(N__6203));
    InMux I__1414 (
            .O(N__6223),
            .I(N__6203));
    InMux I__1413 (
            .O(N__6222),
            .I(N__6203));
    LocalMux I__1412 (
            .O(N__6219),
            .I(N__6200));
    LocalMux I__1411 (
            .O(N__6212),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__1410 (
            .O(N__6203),
            .I(\U409_TICK.TICK603_10 ));
    Odrv4 I__1409 (
            .O(N__6200),
            .I(\U409_TICK.TICK603_10 ));
    CascadeMux I__1408 (
            .O(N__6193),
            .I(N__6189));
    InMux I__1407 (
            .O(N__6192),
            .I(N__6183));
    InMux I__1406 (
            .O(N__6189),
            .I(N__6183));
    InMux I__1405 (
            .O(N__6188),
            .I(N__6180));
    LocalMux I__1404 (
            .O(N__6183),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__1403 (
            .O(N__6180),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    CascadeMux I__1402 (
            .O(N__6175),
            .I(N__6171));
    CascadeMux I__1401 (
            .O(N__6174),
            .I(N__6166));
    InMux I__1400 (
            .O(N__6171),
            .I(N__6161));
    InMux I__1399 (
            .O(N__6170),
            .I(N__6161));
    InMux I__1398 (
            .O(N__6169),
            .I(N__6158));
    InMux I__1397 (
            .O(N__6166),
            .I(N__6155));
    LocalMux I__1396 (
            .O(N__6161),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__1395 (
            .O(N__6158),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__1394 (
            .O(N__6155),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__1393 (
            .O(N__6148),
            .I(N__6144));
    InMux I__1392 (
            .O(N__6147),
            .I(N__6141));
    LocalMux I__1391 (
            .O(N__6144),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__1390 (
            .O(N__6141),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__1389 (
            .O(N__6136),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__1388 (
            .O(N__6133),
            .I(N__6130));
    LocalMux I__1387 (
            .O(N__6130),
            .I(N__6126));
    InMux I__1386 (
            .O(N__6129),
            .I(N__6123));
    Odrv4 I__1385 (
            .O(N__6126),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__1384 (
            .O(N__6123),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__1383 (
            .O(N__6118),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    CascadeMux I__1382 (
            .O(N__6115),
            .I(N__6112));
    InMux I__1381 (
            .O(N__6112),
            .I(N__6108));
    InMux I__1380 (
            .O(N__6111),
            .I(N__6105));
    LocalMux I__1379 (
            .O(N__6108),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__1378 (
            .O(N__6105),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    InMux I__1377 (
            .O(N__6100),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__1376 (
            .O(N__6097),
            .I(N__6093));
    InMux I__1375 (
            .O(N__6096),
            .I(N__6090));
    LocalMux I__1374 (
            .O(N__6093),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__1373 (
            .O(N__6090),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__1372 (
            .O(N__6085),
            .I(N__6082));
    LocalMux I__1371 (
            .O(N__6082),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__1370 (
            .O(N__6079),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    InMux I__1369 (
            .O(N__6076),
            .I(N__6072));
    InMux I__1368 (
            .O(N__6075),
            .I(N__6069));
    LocalMux I__1367 (
            .O(N__6072),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__1366 (
            .O(N__6069),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__1365 (
            .O(N__6064),
            .I(N__6060));
    InMux I__1364 (
            .O(N__6063),
            .I(N__6057));
    LocalMux I__1363 (
            .O(N__6060),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__1362 (
            .O(N__6057),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    InMux I__1361 (
            .O(N__6052),
            .I(N__6049));
    LocalMux I__1360 (
            .O(N__6049),
            .I(\U409_TICK.TICK603_11 ));
    CascadeMux I__1359 (
            .O(N__6046),
            .I(\U409_TICK.TICK603_8_cascade_ ));
    InMux I__1358 (
            .O(N__6043),
            .I(N__6039));
    InMux I__1357 (
            .O(N__6042),
            .I(N__6036));
    LocalMux I__1356 (
            .O(N__6039),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__1355 (
            .O(N__6036),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    CascadeMux I__1354 (
            .O(N__6031),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    InMux I__1353 (
            .O(N__6028),
            .I(N__6025));
    LocalMux I__1352 (
            .O(N__6025),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__1351 (
            .O(N__6022),
            .I(N__6018));
    InMux I__1350 (
            .O(N__6021),
            .I(N__6015));
    LocalMux I__1349 (
            .O(N__6018),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__1348 (
            .O(N__6015),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__1347 (
            .O(N__6010),
            .I(N__5998));
    InMux I__1346 (
            .O(N__6009),
            .I(N__5998));
    InMux I__1345 (
            .O(N__6008),
            .I(N__5993));
    InMux I__1344 (
            .O(N__6007),
            .I(N__5993));
    InMux I__1343 (
            .O(N__6006),
            .I(N__5984));
    InMux I__1342 (
            .O(N__6005),
            .I(N__5984));
    InMux I__1341 (
            .O(N__6004),
            .I(N__5984));
    InMux I__1340 (
            .O(N__6003),
            .I(N__5984));
    LocalMux I__1339 (
            .O(N__5998),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__1338 (
            .O(N__5993),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__1337 (
            .O(N__5984),
            .I(\U409_TICK.TICK503_10 ));
    CascadeMux I__1336 (
            .O(N__5977),
            .I(N__5973));
    InMux I__1335 (
            .O(N__5976),
            .I(N__5964));
    InMux I__1334 (
            .O(N__5973),
            .I(N__5961));
    InMux I__1333 (
            .O(N__5972),
            .I(N__5958));
    InMux I__1332 (
            .O(N__5971),
            .I(N__5947));
    InMux I__1331 (
            .O(N__5970),
            .I(N__5947));
    InMux I__1330 (
            .O(N__5969),
            .I(N__5947));
    InMux I__1329 (
            .O(N__5968),
            .I(N__5947));
    InMux I__1328 (
            .O(N__5967),
            .I(N__5947));
    LocalMux I__1327 (
            .O(N__5964),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__1326 (
            .O(N__5961),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__1325 (
            .O(N__5958),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__1324 (
            .O(N__5947),
            .I(\U409_TICK.TICK503_14 ));
    CascadeMux I__1323 (
            .O(N__5938),
            .I(N__5931));
    CascadeMux I__1322 (
            .O(N__5937),
            .I(N__5928));
    InMux I__1321 (
            .O(N__5936),
            .I(N__5920));
    InMux I__1320 (
            .O(N__5935),
            .I(N__5920));
    InMux I__1319 (
            .O(N__5934),
            .I(N__5909));
    InMux I__1318 (
            .O(N__5931),
            .I(N__5909));
    InMux I__1317 (
            .O(N__5928),
            .I(N__5909));
    InMux I__1316 (
            .O(N__5927),
            .I(N__5909));
    InMux I__1315 (
            .O(N__5926),
            .I(N__5909));
    InMux I__1314 (
            .O(N__5925),
            .I(N__5906));
    LocalMux I__1313 (
            .O(N__5920),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1312 (
            .O(N__5909),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1311 (
            .O(N__5906),
            .I(\U409_TICK.TICK503_9 ));
    IoInMux I__1310 (
            .O(N__5899),
            .I(N__5896));
    LocalMux I__1309 (
            .O(N__5896),
            .I(N__5893));
    IoSpan4Mux I__1308 (
            .O(N__5893),
            .I(N__5890));
    Span4Mux_s3_v I__1307 (
            .O(N__5890),
            .I(N__5887));
    Span4Mux_v I__1306 (
            .O(N__5887),
            .I(N__5883));
    InMux I__1305 (
            .O(N__5886),
            .I(N__5880));
    Odrv4 I__1304 (
            .O(N__5883),
            .I(TICK60_c));
    LocalMux I__1303 (
            .O(N__5880),
            .I(TICK60_c));
    CascadeMux I__1302 (
            .O(N__5875),
            .I(N__5872));
    InMux I__1301 (
            .O(N__5872),
            .I(N__5869));
    LocalMux I__1300 (
            .O(N__5869),
            .I(N__5866));
    Odrv4 I__1299 (
            .O(N__5866),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__1298 (
            .O(N__5863),
            .I(N__5860));
    LocalMux I__1297 (
            .O(N__5860),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    CascadeMux I__1296 (
            .O(N__5857),
            .I(N__5854));
    InMux I__1295 (
            .O(N__5854),
            .I(N__5851));
    LocalMux I__1294 (
            .O(N__5851),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__1293 (
            .O(N__5848),
            .I(N__5845));
    LocalMux I__1292 (
            .O(N__5845),
            .I(\U409_TICK.TICK503_11 ));
    CascadeMux I__1291 (
            .O(N__5842),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    InMux I__1290 (
            .O(N__5839),
            .I(N__5835));
    InMux I__1289 (
            .O(N__5838),
            .I(N__5832));
    LocalMux I__1288 (
            .O(N__5835),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__1287 (
            .O(N__5832),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__1286 (
            .O(N__5827),
            .I(N__5823));
    InMux I__1285 (
            .O(N__5826),
            .I(N__5820));
    LocalMux I__1284 (
            .O(N__5823),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__1283 (
            .O(N__5820),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    CascadeMux I__1282 (
            .O(N__5815),
            .I(N__5811));
    InMux I__1281 (
            .O(N__5814),
            .I(N__5807));
    InMux I__1280 (
            .O(N__5811),
            .I(N__5804));
    InMux I__1279 (
            .O(N__5810),
            .I(N__5801));
    LocalMux I__1278 (
            .O(N__5807),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__1277 (
            .O(N__5804),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__1276 (
            .O(N__5801),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    InMux I__1275 (
            .O(N__5794),
            .I(N__5790));
    InMux I__1274 (
            .O(N__5793),
            .I(N__5787));
    LocalMux I__1273 (
            .O(N__5790),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__1272 (
            .O(N__5787),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    CascadeMux I__1271 (
            .O(N__5782),
            .I(N__5779));
    InMux I__1270 (
            .O(N__5779),
            .I(N__5776));
    LocalMux I__1269 (
            .O(N__5776),
            .I(N__5773));
    Odrv4 I__1268 (
            .O(N__5773),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__1267 (
            .O(N__5770),
            .I(N__5765));
    InMux I__1266 (
            .O(N__5769),
            .I(N__5760));
    InMux I__1265 (
            .O(N__5768),
            .I(N__5760));
    LocalMux I__1264 (
            .O(N__5765),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1263 (
            .O(N__5760),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    InMux I__1262 (
            .O(N__5755),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__1261 (
            .O(N__5752),
            .I(N__5747));
    InMux I__1260 (
            .O(N__5751),
            .I(N__5742));
    InMux I__1259 (
            .O(N__5750),
            .I(N__5742));
    LocalMux I__1258 (
            .O(N__5747),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1257 (
            .O(N__5742),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    InMux I__1256 (
            .O(N__5737),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__1255 (
            .O(N__5734),
            .I(N__5727));
    InMux I__1254 (
            .O(N__5733),
            .I(N__5724));
    InMux I__1253 (
            .O(N__5732),
            .I(N__5717));
    InMux I__1252 (
            .O(N__5731),
            .I(N__5717));
    InMux I__1251 (
            .O(N__5730),
            .I(N__5717));
    LocalMux I__1250 (
            .O(N__5727),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1249 (
            .O(N__5724),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1248 (
            .O(N__5717),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    InMux I__1247 (
            .O(N__5710),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__1246 (
            .O(N__5707),
            .I(N__5701));
    InMux I__1245 (
            .O(N__5706),
            .I(N__5701));
    LocalMux I__1244 (
            .O(N__5701),
            .I(\U409_CIA.CIA_CLK_COUNT11 ));
    InMux I__1243 (
            .O(N__5698),
            .I(N__5693));
    InMux I__1242 (
            .O(N__5697),
            .I(N__5688));
    InMux I__1241 (
            .O(N__5696),
            .I(N__5688));
    LocalMux I__1240 (
            .O(N__5693),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1239 (
            .O(N__5688),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    InMux I__1238 (
            .O(N__5683),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    InMux I__1237 (
            .O(N__5680),
            .I(N__5675));
    InMux I__1236 (
            .O(N__5679),
            .I(N__5672));
    InMux I__1235 (
            .O(N__5678),
            .I(N__5669));
    LocalMux I__1234 (
            .O(N__5675),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__1233 (
            .O(N__5672),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__1232 (
            .O(N__5669),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    InMux I__1231 (
            .O(N__5662),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ));
    InMux I__1230 (
            .O(N__5659),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ));
    CascadeMux I__1229 (
            .O(N__5656),
            .I(N__5652));
    InMux I__1228 (
            .O(N__5655),
            .I(N__5648));
    InMux I__1227 (
            .O(N__5652),
            .I(N__5645));
    InMux I__1226 (
            .O(N__5651),
            .I(N__5642));
    LocalMux I__1225 (
            .O(N__5648),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__1224 (
            .O(N__5645),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__1223 (
            .O(N__5642),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    CascadeMux I__1222 (
            .O(N__5635),
            .I(N__5628));
    InMux I__1221 (
            .O(N__5634),
            .I(N__5622));
    InMux I__1220 (
            .O(N__5633),
            .I(N__5622));
    InMux I__1219 (
            .O(N__5632),
            .I(N__5619));
    InMux I__1218 (
            .O(N__5631),
            .I(N__5612));
    InMux I__1217 (
            .O(N__5628),
            .I(N__5612));
    InMux I__1216 (
            .O(N__5627),
            .I(N__5612));
    LocalMux I__1215 (
            .O(N__5622),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1214 (
            .O(N__5619),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1213 (
            .O(N__5612),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    ClkMux I__1212 (
            .O(N__5605),
            .I(N__5596));
    ClkMux I__1211 (
            .O(N__5604),
            .I(N__5596));
    ClkMux I__1210 (
            .O(N__5603),
            .I(N__5596));
    GlobalMux I__1209 (
            .O(N__5596),
            .I(N__5593));
    gio2CtrlBuf I__1208 (
            .O(N__5593),
            .I(CLK28_IN_c_g));
    InMux I__1207 (
            .O(N__5590),
            .I(bfn_13_3_0_));
    InMux I__1206 (
            .O(N__5587),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__1205 (
            .O(N__5584),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__1204 (
            .O(N__5581),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__1203 (
            .O(N__5578),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__1202 (
            .O(N__5575),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__1201 (
            .O(N__5572),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__1200 (
            .O(N__5569),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__1199 (
            .O(N__5566),
            .I(N__5559));
    InMux I__1198 (
            .O(N__5565),
            .I(N__5552));
    InMux I__1197 (
            .O(N__5564),
            .I(N__5552));
    InMux I__1196 (
            .O(N__5563),
            .I(N__5552));
    InMux I__1195 (
            .O(N__5562),
            .I(N__5549));
    LocalMux I__1194 (
            .O(N__5559),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1193 (
            .O(N__5552),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1192 (
            .O(N__5549),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    InMux I__1191 (
            .O(N__5542),
            .I(N__5539));
    LocalMux I__1190 (
            .O(N__5539),
            .I(\U409_CIA.CLK_CIA6_1 ));
    CascadeMux I__1189 (
            .O(N__5536),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    IoInMux I__1188 (
            .O(N__5533),
            .I(N__5530));
    LocalMux I__1187 (
            .O(N__5530),
            .I(N__5527));
    Span4Mux_s2_v I__1186 (
            .O(N__5527),
            .I(N__5524));
    Span4Mux_v I__1185 (
            .O(N__5524),
            .I(N__5521));
    Span4Mux_h I__1184 (
            .O(N__5521),
            .I(N__5517));
    InMux I__1183 (
            .O(N__5520),
            .I(N__5514));
    Odrv4 I__1182 (
            .O(N__5517),
            .I(TICK50_c));
    LocalMux I__1181 (
            .O(N__5514),
            .I(TICK50_c));
    InMux I__1180 (
            .O(N__5509),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__1179 (
            .O(N__5506),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__1178 (
            .O(N__5503),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__1177 (
            .O(N__5500),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    InMux I__1176 (
            .O(N__5497),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__1175 (
            .O(N__5494),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    CascadeMux I__1174 (
            .O(N__5491),
            .I(N__5488));
    InMux I__1173 (
            .O(N__5488),
            .I(N__5485));
    LocalMux I__1172 (
            .O(N__5485),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__1171 (
            .O(N__5482),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__1170 (
            .O(N__5479),
            .I(N__5476));
    LocalMux I__1169 (
            .O(N__5476),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ));
    InMux I__1168 (
            .O(N__5473),
            .I(N__5469));
    InMux I__1167 (
            .O(N__5472),
            .I(N__5466));
    LocalMux I__1166 (
            .O(N__5469),
            .I(\U409_CIA.N_91 ));
    LocalMux I__1165 (
            .O(N__5466),
            .I(\U409_CIA.N_91 ));
    InMux I__1164 (
            .O(N__5461),
            .I(N__5458));
    LocalMux I__1163 (
            .O(N__5458),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_2_1 ));
    CascadeMux I__1162 (
            .O(N__5455),
            .I(\U409_CIA.CLK_CIA_r_1_cascade_ ));
    InMux I__1161 (
            .O(N__5452),
            .I(N__5448));
    InMux I__1160 (
            .O(N__5451),
            .I(N__5445));
    LocalMux I__1159 (
            .O(N__5448),
            .I(\U409_CIA.CLK_CIA6_1_0 ));
    LocalMux I__1158 (
            .O(N__5445),
            .I(\U409_CIA.CLK_CIA6_1_0 ));
    IoInMux I__1157 (
            .O(N__5440),
            .I(N__5437));
    LocalMux I__1156 (
            .O(N__5437),
            .I(N__5434));
    Span4Mux_s2_v I__1155 (
            .O(N__5434),
            .I(N__5431));
    Span4Mux_h I__1154 (
            .O(N__5431),
            .I(N__5428));
    Span4Mux_v I__1153 (
            .O(N__5428),
            .I(N__5423));
    InMux I__1152 (
            .O(N__5427),
            .I(N__5420));
    CascadeMux I__1151 (
            .O(N__5426),
            .I(N__5416));
    Sp12to4 I__1150 (
            .O(N__5423),
            .I(N__5411));
    LocalMux I__1149 (
            .O(N__5420),
            .I(N__5411));
    InMux I__1148 (
            .O(N__5419),
            .I(N__5406));
    InMux I__1147 (
            .O(N__5416),
            .I(N__5406));
    Odrv12 I__1146 (
            .O(N__5411),
            .I(CLK_CIA_c));
    LocalMux I__1145 (
            .O(N__5406),
            .I(CLK_CIA_c));
    CascadeMux I__1144 (
            .O(N__5401),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    CascadeMux I__1143 (
            .O(N__5398),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    InMux I__1142 (
            .O(N__5395),
            .I(N__5388));
    InMux I__1141 (
            .O(N__5394),
            .I(N__5385));
    InMux I__1140 (
            .O(N__5393),
            .I(N__5378));
    InMux I__1139 (
            .O(N__5392),
            .I(N__5378));
    InMux I__1138 (
            .O(N__5391),
            .I(N__5378));
    LocalMux I__1137 (
            .O(N__5388),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__1136 (
            .O(N__5385),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__1135 (
            .O(N__5378),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__1134 (
            .O(N__5371),
            .I(N__5368));
    LocalMux I__1133 (
            .O(N__5368),
            .I(N__5359));
    InMux I__1132 (
            .O(N__5367),
            .I(N__5356));
    InMux I__1131 (
            .O(N__5366),
            .I(N__5353));
    InMux I__1130 (
            .O(N__5365),
            .I(N__5350));
    CascadeMux I__1129 (
            .O(N__5364),
            .I(N__5345));
    CascadeMux I__1128 (
            .O(N__5363),
            .I(N__5342));
    CascadeMux I__1127 (
            .O(N__5362),
            .I(N__5339));
    Span4Mux_h I__1126 (
            .O(N__5359),
            .I(N__5334));
    LocalMux I__1125 (
            .O(N__5356),
            .I(N__5334));
    LocalMux I__1124 (
            .O(N__5353),
            .I(N__5329));
    LocalMux I__1123 (
            .O(N__5350),
            .I(N__5329));
    InMux I__1122 (
            .O(N__5349),
            .I(N__5326));
    InMux I__1121 (
            .O(N__5348),
            .I(N__5319));
    InMux I__1120 (
            .O(N__5345),
            .I(N__5319));
    InMux I__1119 (
            .O(N__5342),
            .I(N__5319));
    InMux I__1118 (
            .O(N__5339),
            .I(N__5316));
    Span4Mux_v I__1117 (
            .O(N__5334),
            .I(N__5312));
    Span4Mux_h I__1116 (
            .O(N__5329),
            .I(N__5309));
    LocalMux I__1115 (
            .O(N__5326),
            .I(N__5302));
    LocalMux I__1114 (
            .O(N__5319),
            .I(N__5302));
    LocalMux I__1113 (
            .O(N__5316),
            .I(N__5302));
    CascadeMux I__1112 (
            .O(N__5315),
            .I(N__5298));
    Span4Mux_h I__1111 (
            .O(N__5312),
            .I(N__5290));
    Span4Mux_v I__1110 (
            .O(N__5309),
            .I(N__5290));
    Span4Mux_h I__1109 (
            .O(N__5302),
            .I(N__5290));
    InMux I__1108 (
            .O(N__5301),
            .I(N__5287));
    InMux I__1107 (
            .O(N__5298),
            .I(N__5282));
    InMux I__1106 (
            .O(N__5297),
            .I(N__5282));
    Span4Mux_v I__1105 (
            .O(N__5290),
            .I(N__5277));
    LocalMux I__1104 (
            .O(N__5287),
            .I(N__5274));
    LocalMux I__1103 (
            .O(N__5282),
            .I(N__5271));
    InMux I__1102 (
            .O(N__5281),
            .I(N__5268));
    InMux I__1101 (
            .O(N__5280),
            .I(N__5265));
    Sp12to4 I__1100 (
            .O(N__5277),
            .I(N__5254));
    Span12Mux_v I__1099 (
            .O(N__5274),
            .I(N__5254));
    Sp12to4 I__1098 (
            .O(N__5271),
            .I(N__5254));
    LocalMux I__1097 (
            .O(N__5268),
            .I(N__5254));
    LocalMux I__1096 (
            .O(N__5265),
            .I(N__5254));
    Span12Mux_v I__1095 (
            .O(N__5254),
            .I(N__5251));
    Span12Mux_h I__1094 (
            .O(N__5251),
            .I(N__5248));
    Odrv12 I__1093 (
            .O(N__5248),
            .I(RESETn_c));
    SRMux I__1092 (
            .O(N__5245),
            .I(N__5240));
    SRMux I__1091 (
            .O(N__5244),
            .I(N__5234));
    SRMux I__1090 (
            .O(N__5243),
            .I(N__5231));
    LocalMux I__1089 (
            .O(N__5240),
            .I(N__5227));
    SRMux I__1088 (
            .O(N__5239),
            .I(N__5224));
    SRMux I__1087 (
            .O(N__5238),
            .I(N__5221));
    SRMux I__1086 (
            .O(N__5237),
            .I(N__5218));
    LocalMux I__1085 (
            .O(N__5234),
            .I(N__5215));
    LocalMux I__1084 (
            .O(N__5231),
            .I(N__5212));
    SRMux I__1083 (
            .O(N__5230),
            .I(N__5209));
    Span4Mux_h I__1082 (
            .O(N__5227),
            .I(N__5204));
    LocalMux I__1081 (
            .O(N__5224),
            .I(N__5204));
    LocalMux I__1080 (
            .O(N__5221),
            .I(N__5201));
    LocalMux I__1079 (
            .O(N__5218),
            .I(N__5196));
    Span4Mux_h I__1078 (
            .O(N__5215),
            .I(N__5196));
    Span4Mux_v I__1077 (
            .O(N__5212),
            .I(N__5193));
    LocalMux I__1076 (
            .O(N__5209),
            .I(N__5188));
    Sp12to4 I__1075 (
            .O(N__5204),
            .I(N__5188));
    Span4Mux_v I__1074 (
            .O(N__5201),
            .I(N__5183));
    Span4Mux_v I__1073 (
            .O(N__5196),
            .I(N__5183));
    Odrv4 I__1072 (
            .O(N__5193),
            .I(RESETn_c_i));
    Odrv12 I__1071 (
            .O(N__5188),
            .I(RESETn_c_i));
    Odrv4 I__1070 (
            .O(N__5183),
            .I(RESETn_c_i));
    CascadeMux I__1069 (
            .O(N__5176),
            .I(\U409_CIA.N_93_cascade_ ));
    CascadeMux I__1068 (
            .O(N__5173),
            .I(\U409_CIA.VMA_RNOZ0Z_1_cascade_ ));
    InMux I__1067 (
            .O(N__5170),
            .I(N__5167));
    LocalMux I__1066 (
            .O(N__5167),
            .I(N__5164));
    Span4Mux_v I__1065 (
            .O(N__5164),
            .I(N__5161));
    Odrv4 I__1064 (
            .O(N__5161),
            .I(\U409_CIA.VMA_3_0_a2_2 ));
    InMux I__1063 (
            .O(N__5158),
            .I(N__5154));
    InMux I__1062 (
            .O(N__5157),
            .I(N__5151));
    LocalMux I__1061 (
            .O(N__5154),
            .I(N__5145));
    LocalMux I__1060 (
            .O(N__5151),
            .I(N__5145));
    InMux I__1059 (
            .O(N__5150),
            .I(N__5142));
    Odrv12 I__1058 (
            .O(N__5145),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__1057 (
            .O(N__5142),
            .I(\U409_CIA.VMAZ0 ));
    CascadeMux I__1056 (
            .O(N__5137),
            .I(\U409_CIA.N_91_cascade_ ));
    InMux I__1055 (
            .O(N__5134),
            .I(N__5124));
    InMux I__1054 (
            .O(N__5133),
            .I(N__5124));
    InMux I__1053 (
            .O(N__5132),
            .I(N__5117));
    InMux I__1052 (
            .O(N__5131),
            .I(N__5117));
    InMux I__1051 (
            .O(N__5130),
            .I(N__5117));
    InMux I__1050 (
            .O(N__5129),
            .I(N__5114));
    LocalMux I__1049 (
            .O(N__5124),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1048 (
            .O(N__5117),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1047 (
            .O(N__5114),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__1046 (
            .O(N__5107),
            .I(N__5102));
    CascadeMux I__1045 (
            .O(N__5106),
            .I(N__5099));
    CascadeMux I__1044 (
            .O(N__5105),
            .I(N__5095));
    InMux I__1043 (
            .O(N__5102),
            .I(N__5085));
    InMux I__1042 (
            .O(N__5099),
            .I(N__5085));
    InMux I__1041 (
            .O(N__5098),
            .I(N__5085));
    InMux I__1040 (
            .O(N__5095),
            .I(N__5078));
    InMux I__1039 (
            .O(N__5094),
            .I(N__5078));
    InMux I__1038 (
            .O(N__5093),
            .I(N__5078));
    InMux I__1037 (
            .O(N__5092),
            .I(N__5075));
    LocalMux I__1036 (
            .O(N__5085),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1035 (
            .O(N__5078),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1034 (
            .O(N__5075),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    InMux I__1033 (
            .O(N__5068),
            .I(N__5065));
    LocalMux I__1032 (
            .O(N__5065),
            .I(N__5056));
    InMux I__1031 (
            .O(N__5064),
            .I(N__5049));
    InMux I__1030 (
            .O(N__5063),
            .I(N__5049));
    InMux I__1029 (
            .O(N__5062),
            .I(N__5049));
    InMux I__1028 (
            .O(N__5061),
            .I(N__5044));
    InMux I__1027 (
            .O(N__5060),
            .I(N__5044));
    InMux I__1026 (
            .O(N__5059),
            .I(N__5041));
    Odrv4 I__1025 (
            .O(N__5056),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1024 (
            .O(N__5049),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1023 (
            .O(N__5044),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1022 (
            .O(N__5041),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__1021 (
            .O(N__5032),
            .I(N__5029));
    LocalMux I__1020 (
            .O(N__5029),
            .I(\U409_TRANSFER_ACK.N_23 ));
    IoInMux I__1019 (
            .O(N__5026),
            .I(N__5023));
    LocalMux I__1018 (
            .O(N__5023),
            .I(N__5020));
    Span4Mux_s2_v I__1017 (
            .O(N__5020),
            .I(N__5017));
    Span4Mux_v I__1016 (
            .O(N__5017),
            .I(N__5014));
    Odrv4 I__1015 (
            .O(N__5014),
            .I(CONSTANT_ONE_NET));
    InMux I__1014 (
            .O(N__5011),
            .I(N__5008));
    LocalMux I__1013 (
            .O(N__5008),
            .I(N__5005));
    Span4Mux_v I__1012 (
            .O(N__5005),
            .I(N__5002));
    Sp12to4 I__1011 (
            .O(N__5002),
            .I(N__4999));
    Span12Mux_h I__1010 (
            .O(N__4999),
            .I(N__4996));
    Odrv12 I__1009 (
            .O(N__4996),
            .I(A_c_13));
    IoInMux I__1008 (
            .O(N__4993),
            .I(N__4990));
    LocalMux I__1007 (
            .O(N__4990),
            .I(N__4987));
    IoSpan4Mux I__1006 (
            .O(N__4987),
            .I(N__4984));
    Span4Mux_s2_h I__1005 (
            .O(N__4984),
            .I(N__4981));
    Sp12to4 I__1004 (
            .O(N__4981),
            .I(N__4978));
    Span12Mux_h I__1003 (
            .O(N__4978),
            .I(N__4975));
    Odrv12 I__1002 (
            .O(N__4975),
            .I(U409_ADDRESS_DECODE_un1_CIACS1n_i));
    InMux I__1001 (
            .O(N__4972),
            .I(N__4969));
    LocalMux I__1000 (
            .O(N__4969),
            .I(CIA_ENABLE));
    CascadeMux I__999 (
            .O(N__4966),
            .I(CIA_ENABLE_cascade_));
    InMux I__998 (
            .O(N__4963),
            .I(N__4960));
    LocalMux I__997 (
            .O(N__4960),
            .I(N__4957));
    Span12Mux_s10_v I__996 (
            .O(N__4957),
            .I(N__4954));
    Span12Mux_h I__995 (
            .O(N__4954),
            .I(N__4951));
    Odrv12 I__994 (
            .O(N__4951),
            .I(A_c_12));
    IoInMux I__993 (
            .O(N__4948),
            .I(N__4945));
    LocalMux I__992 (
            .O(N__4945),
            .I(N__4942));
    IoSpan4Mux I__991 (
            .O(N__4942),
            .I(N__4939));
    IoSpan4Mux I__990 (
            .O(N__4939),
            .I(N__4936));
    Sp12to4 I__989 (
            .O(N__4936),
            .I(N__4933));
    Span12Mux_s7_h I__988 (
            .O(N__4933),
            .I(N__4930));
    Odrv12 I__987 (
            .O(N__4930),
            .I(U409_ADDRESS_DECODE_un1_CIACS0n_i));
    InMux I__986 (
            .O(N__4927),
            .I(N__4922));
    InMux I__985 (
            .O(N__4926),
            .I(N__4917));
    InMux I__984 (
            .O(N__4925),
            .I(N__4917));
    LocalMux I__983 (
            .O(N__4922),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__982 (
            .O(N__4917),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    CascadeMux I__981 (
            .O(N__4912),
            .I(N__4909));
    InMux I__980 (
            .O(N__4909),
            .I(N__4903));
    InMux I__979 (
            .O(N__4908),
            .I(N__4903));
    LocalMux I__978 (
            .O(N__4903),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    CascadeMux I__977 (
            .O(N__4900),
            .I(N__4894));
    InMux I__976 (
            .O(N__4899),
            .I(N__4891));
    InMux I__975 (
            .O(N__4898),
            .I(N__4884));
    InMux I__974 (
            .O(N__4897),
            .I(N__4884));
    InMux I__973 (
            .O(N__4894),
            .I(N__4884));
    LocalMux I__972 (
            .O(N__4891),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    LocalMux I__971 (
            .O(N__4884),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    InMux I__970 (
            .O(N__4879),
            .I(N__4876));
    LocalMux I__969 (
            .O(N__4876),
            .I(\U409_TRANSFER_ACK.N_64 ));
    CascadeMux I__968 (
            .O(N__4873),
            .I(\U409_TRANSFER_ACK.N_63_cascade_ ));
    CascadeMux I__967 (
            .O(N__4870),
            .I(\U409_TRANSFER_ACK.m9_i_1_cascade_ ));
    InMux I__966 (
            .O(N__4867),
            .I(N__4861));
    InMux I__965 (
            .O(N__4866),
            .I(N__4861));
    LocalMux I__964 (
            .O(N__4861),
            .I(\U409_TRANSFER_ACK.N_45 ));
    InMux I__963 (
            .O(N__4858),
            .I(N__4853));
    InMux I__962 (
            .O(N__4857),
            .I(N__4848));
    InMux I__961 (
            .O(N__4856),
            .I(N__4848));
    LocalMux I__960 (
            .O(N__4853),
            .I(\U409_TRANSFER_ACK.N_73 ));
    LocalMux I__959 (
            .O(N__4848),
            .I(\U409_TRANSFER_ACK.N_73 ));
    InMux I__958 (
            .O(N__4843),
            .I(N__4840));
    LocalMux I__957 (
            .O(N__4840),
            .I(\U409_TRANSFER_ACK.N_60 ));
    InMux I__956 (
            .O(N__4837),
            .I(N__4830));
    InMux I__955 (
            .O(N__4836),
            .I(N__4821));
    InMux I__954 (
            .O(N__4835),
            .I(N__4821));
    InMux I__953 (
            .O(N__4834),
            .I(N__4821));
    InMux I__952 (
            .O(N__4833),
            .I(N__4821));
    LocalMux I__951 (
            .O(N__4830),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__950 (
            .O(N__4821),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    CascadeMux I__949 (
            .O(N__4816),
            .I(\U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_ ));
    InMux I__948 (
            .O(N__4813),
            .I(N__4810));
    LocalMux I__947 (
            .O(N__4810),
            .I(\U409_TRANSFER_ACK.N_65 ));
    CascadeMux I__946 (
            .O(N__4807),
            .I(N__4800));
    CascadeMux I__945 (
            .O(N__4806),
            .I(N__4797));
    CascadeMux I__944 (
            .O(N__4805),
            .I(N__4794));
    IoInMux I__943 (
            .O(N__4804),
            .I(N__4791));
    InMux I__942 (
            .O(N__4803),
            .I(N__4788));
    InMux I__941 (
            .O(N__4800),
            .I(N__4785));
    InMux I__940 (
            .O(N__4797),
            .I(N__4782));
    InMux I__939 (
            .O(N__4794),
            .I(N__4779));
    LocalMux I__938 (
            .O(N__4791),
            .I(N__4775));
    LocalMux I__937 (
            .O(N__4788),
            .I(N__4770));
    LocalMux I__936 (
            .O(N__4785),
            .I(N__4767));
    LocalMux I__935 (
            .O(N__4782),
            .I(N__4764));
    LocalMux I__934 (
            .O(N__4779),
            .I(N__4761));
    InMux I__933 (
            .O(N__4778),
            .I(N__4758));
    IoSpan4Mux I__932 (
            .O(N__4775),
            .I(N__4755));
    InMux I__931 (
            .O(N__4774),
            .I(N__4752));
    InMux I__930 (
            .O(N__4773),
            .I(N__4749));
    Span4Mux_v I__929 (
            .O(N__4770),
            .I(N__4744));
    Span4Mux_h I__928 (
            .O(N__4767),
            .I(N__4744));
    Span4Mux_v I__927 (
            .O(N__4764),
            .I(N__4737));
    Span4Mux_h I__926 (
            .O(N__4761),
            .I(N__4737));
    LocalMux I__925 (
            .O(N__4758),
            .I(N__4737));
    Span4Mux_s0_v I__924 (
            .O(N__4755),
            .I(N__4734));
    LocalMux I__923 (
            .O(N__4752),
            .I(N__4731));
    LocalMux I__922 (
            .O(N__4749),
            .I(N__4728));
    Span4Mux_v I__921 (
            .O(N__4744),
            .I(N__4723));
    Span4Mux_h I__920 (
            .O(N__4737),
            .I(N__4723));
    Sp12to4 I__919 (
            .O(N__4734),
            .I(N__4720));
    Span4Mux_h I__918 (
            .O(N__4731),
            .I(N__4715));
    Span4Mux_h I__917 (
            .O(N__4728),
            .I(N__4715));
    Span4Mux_v I__916 (
            .O(N__4723),
            .I(N__4712));
    Span12Mux_v I__915 (
            .O(N__4720),
            .I(N__4709));
    Sp12to4 I__914 (
            .O(N__4715),
            .I(N__4706));
    Span4Mux_v I__913 (
            .O(N__4712),
            .I(N__4703));
    Span12Mux_v I__912 (
            .O(N__4709),
            .I(N__4700));
    Span12Mux_v I__911 (
            .O(N__4706),
            .I(N__4697));
    Span4Mux_v I__910 (
            .O(N__4703),
            .I(N__4694));
    Odrv12 I__909 (
            .O(N__4700),
            .I(CLK40_IN_c));
    Odrv12 I__908 (
            .O(N__4697),
            .I(CLK40_IN_c));
    Odrv4 I__907 (
            .O(N__4694),
            .I(CLK40_IN_c));
    CascadeMux I__906 (
            .O(N__4687),
            .I(N__4682));
    InMux I__905 (
            .O(N__4686),
            .I(N__4676));
    InMux I__904 (
            .O(N__4685),
            .I(N__4673));
    InMux I__903 (
            .O(N__4682),
            .I(N__4664));
    InMux I__902 (
            .O(N__4681),
            .I(N__4664));
    InMux I__901 (
            .O(N__4680),
            .I(N__4664));
    InMux I__900 (
            .O(N__4679),
            .I(N__4664));
    LocalMux I__899 (
            .O(N__4676),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__898 (
            .O(N__4673),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__897 (
            .O(N__4664),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    InMux I__896 (
            .O(N__4657),
            .I(N__4654));
    LocalMux I__895 (
            .O(N__4654),
            .I(\U409_TRANSFER_ACK.N_68 ));
    CascadeMux I__894 (
            .O(N__4651),
            .I(N__4647));
    InMux I__893 (
            .O(N__4650),
            .I(N__4644));
    InMux I__892 (
            .O(N__4647),
            .I(N__4641));
    LocalMux I__891 (
            .O(N__4644),
            .I(N__4638));
    LocalMux I__890 (
            .O(N__4641),
            .I(N__4635));
    Span4Mux_v I__889 (
            .O(N__4638),
            .I(N__4631));
    Span4Mux_v I__888 (
            .O(N__4635),
            .I(N__4628));
    InMux I__887 (
            .O(N__4634),
            .I(N__4625));
    Sp12to4 I__886 (
            .O(N__4631),
            .I(N__4618));
    Sp12to4 I__885 (
            .O(N__4628),
            .I(N__4618));
    LocalMux I__884 (
            .O(N__4625),
            .I(N__4618));
    Span12Mux_h I__883 (
            .O(N__4618),
            .I(N__4615));
    Span12Mux_v I__882 (
            .O(N__4615),
            .I(N__4612));
    Odrv12 I__881 (
            .O(N__4612),
            .I(TSn_c));
    CascadeMux I__880 (
            .O(N__4609),
            .I(N__4606));
    InMux I__879 (
            .O(N__4606),
            .I(N__4601));
    CascadeMux I__878 (
            .O(N__4605),
            .I(N__4597));
    CascadeMux I__877 (
            .O(N__4604),
            .I(N__4594));
    LocalMux I__876 (
            .O(N__4601),
            .I(N__4591));
    InMux I__875 (
            .O(N__4600),
            .I(N__4588));
    InMux I__874 (
            .O(N__4597),
            .I(N__4585));
    InMux I__873 (
            .O(N__4594),
            .I(N__4582));
    Span4Mux_h I__872 (
            .O(N__4591),
            .I(N__4575));
    LocalMux I__871 (
            .O(N__4588),
            .I(N__4575));
    LocalMux I__870 (
            .O(N__4585),
            .I(N__4575));
    LocalMux I__869 (
            .O(N__4582),
            .I(N__4572));
    Span4Mux_v I__868 (
            .O(N__4575),
            .I(N__4569));
    Span12Mux_v I__867 (
            .O(N__4572),
            .I(N__4566));
    Span4Mux_h I__866 (
            .O(N__4569),
            .I(N__4563));
    Odrv12 I__865 (
            .O(N__4566),
            .I(N_76));
    Odrv4 I__864 (
            .O(N__4563),
            .I(N_76));
    InMux I__863 (
            .O(N__4558),
            .I(N__4555));
    LocalMux I__862 (
            .O(N__4555),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ));
    CascadeMux I__861 (
            .O(N__4552),
            .I(N__4549));
    InMux I__860 (
            .O(N__4549),
            .I(N__4546));
    LocalMux I__859 (
            .O(N__4546),
            .I(\U409_TRANSFER_ACK.ROM_TACK_EN_e_1 ));
    InMux I__858 (
            .O(N__4543),
            .I(N__4539));
    InMux I__857 (
            .O(N__4542),
            .I(N__4536));
    LocalMux I__856 (
            .O(N__4539),
            .I(\U409_TRANSFER_ACK.N_28_4 ));
    LocalMux I__855 (
            .O(N__4536),
            .I(\U409_TRANSFER_ACK.N_28_4 ));
    CascadeMux I__854 (
            .O(N__4531),
            .I(N__4527));
    InMux I__853 (
            .O(N__4530),
            .I(N__4524));
    InMux I__852 (
            .O(N__4527),
            .I(N__4521));
    LocalMux I__851 (
            .O(N__4524),
            .I(N__4516));
    LocalMux I__850 (
            .O(N__4521),
            .I(N__4516));
    Span4Mux_v I__849 (
            .O(N__4516),
            .I(N__4513));
    Odrv4 I__848 (
            .O(N__4513),
            .I(\U409_TRANSFER_ACK.N_28_3 ));
    InMux I__847 (
            .O(N__4510),
            .I(N__4505));
    CascadeMux I__846 (
            .O(N__4509),
            .I(N__4499));
    CascadeMux I__845 (
            .O(N__4508),
            .I(N__4495));
    LocalMux I__844 (
            .O(N__4505),
            .I(N__4492));
    InMux I__843 (
            .O(N__4504),
            .I(N__4483));
    InMux I__842 (
            .O(N__4503),
            .I(N__4483));
    InMux I__841 (
            .O(N__4502),
            .I(N__4483));
    InMux I__840 (
            .O(N__4499),
            .I(N__4483));
    InMux I__839 (
            .O(N__4498),
            .I(N__4478));
    InMux I__838 (
            .O(N__4495),
            .I(N__4478));
    Odrv4 I__837 (
            .O(N__4492),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__836 (
            .O(N__4483),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__835 (
            .O(N__4478),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    InMux I__834 (
            .O(N__4471),
            .I(N__4468));
    LocalMux I__833 (
            .O(N__4468),
            .I(un1_RAMSPACEn_i_i_a3));
    InMux I__832 (
            .O(N__4465),
            .I(N__4462));
    LocalMux I__831 (
            .O(N__4462),
            .I(N__4459));
    Span12Mux_h I__830 (
            .O(N__4459),
            .I(N__4456));
    Span12Mux_h I__829 (
            .O(N__4456),
            .I(N__4453));
    Span12Mux_v I__828 (
            .O(N__4453),
            .I(N__4450));
    Odrv12 I__827 (
            .O(N__4450),
            .I(TACKn_in));
    CascadeMux I__826 (
            .O(N__4447),
            .I(un1_REGSPACEn_i_i_a3_0_a2_cascade_));
    SRMux I__825 (
            .O(N__4444),
            .I(N__4440));
    SRMux I__824 (
            .O(N__4443),
            .I(N__4435));
    LocalMux I__823 (
            .O(N__4440),
            .I(N__4432));
    SRMux I__822 (
            .O(N__4439),
            .I(N__4429));
    SRMux I__821 (
            .O(N__4438),
            .I(N__4426));
    LocalMux I__820 (
            .O(N__4435),
            .I(N__4422));
    Span4Mux_v I__819 (
            .O(N__4432),
            .I(N__4419));
    LocalMux I__818 (
            .O(N__4429),
            .I(N__4416));
    LocalMux I__817 (
            .O(N__4426),
            .I(N__4413));
    SRMux I__816 (
            .O(N__4425),
            .I(N__4410));
    Span4Mux_v I__815 (
            .O(N__4422),
            .I(N__4399));
    Span4Mux_v I__814 (
            .O(N__4419),
            .I(N__4399));
    Span4Mux_h I__813 (
            .O(N__4416),
            .I(N__4399));
    Span4Mux_v I__812 (
            .O(N__4413),
            .I(N__4399));
    LocalMux I__811 (
            .O(N__4410),
            .I(N__4399));
    Span4Mux_h I__810 (
            .O(N__4399),
            .I(N__4396));
    Odrv4 I__809 (
            .O(N__4396),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__808 (
            .O(N__4393),
            .I(N__4389));
    CascadeMux I__807 (
            .O(N__4392),
            .I(N__4384));
    LocalMux I__806 (
            .O(N__4389),
            .I(N__4381));
    InMux I__805 (
            .O(N__4388),
            .I(N__4376));
    InMux I__804 (
            .O(N__4387),
            .I(N__4376));
    InMux I__803 (
            .O(N__4384),
            .I(N__4373));
    Span4Mux_v I__802 (
            .O(N__4381),
            .I(N__4367));
    LocalMux I__801 (
            .O(N__4376),
            .I(N__4367));
    LocalMux I__800 (
            .O(N__4373),
            .I(N__4364));
    InMux I__799 (
            .O(N__4372),
            .I(N__4361));
    Odrv4 I__798 (
            .O(N__4367),
            .I(N_90));
    Odrv4 I__797 (
            .O(N__4364),
            .I(N_90));
    LocalMux I__796 (
            .O(N__4361),
            .I(N_90));
    CascadeMux I__795 (
            .O(N__4354),
            .I(N__4348));
    InMux I__794 (
            .O(N__4353),
            .I(N__4343));
    InMux I__793 (
            .O(N__4352),
            .I(N__4343));
    InMux I__792 (
            .O(N__4351),
            .I(N__4338));
    InMux I__791 (
            .O(N__4348),
            .I(N__4338));
    LocalMux I__790 (
            .O(N__4343),
            .I(N__4333));
    LocalMux I__789 (
            .O(N__4338),
            .I(N__4330));
    InMux I__788 (
            .O(N__4337),
            .I(N__4323));
    InMux I__787 (
            .O(N__4336),
            .I(N__4323));
    Span4Mux_v I__786 (
            .O(N__4333),
            .I(N__4318));
    Span4Mux_v I__785 (
            .O(N__4330),
            .I(N__4318));
    InMux I__784 (
            .O(N__4329),
            .I(N__4315));
    InMux I__783 (
            .O(N__4328),
            .I(N__4312));
    LocalMux I__782 (
            .O(N__4323),
            .I(N__4309));
    Span4Mux_h I__781 (
            .O(N__4318),
            .I(N__4305));
    LocalMux I__780 (
            .O(N__4315),
            .I(N__4300));
    LocalMux I__779 (
            .O(N__4312),
            .I(N__4300));
    Span4Mux_v I__778 (
            .O(N__4309),
            .I(N__4297));
    InMux I__777 (
            .O(N__4308),
            .I(N__4294));
    Sp12to4 I__776 (
            .O(N__4305),
            .I(N__4285));
    Span12Mux_h I__775 (
            .O(N__4300),
            .I(N__4285));
    Sp12to4 I__774 (
            .O(N__4297),
            .I(N__4285));
    LocalMux I__773 (
            .O(N__4294),
            .I(N__4285));
    Odrv12 I__772 (
            .O(N__4285),
            .I(A_c_21));
    InMux I__771 (
            .O(N__4282),
            .I(N__4277));
    InMux I__770 (
            .O(N__4281),
            .I(N__4272));
    InMux I__769 (
            .O(N__4280),
            .I(N__4272));
    LocalMux I__768 (
            .O(N__4277),
            .I(N__4269));
    LocalMux I__767 (
            .O(N__4272),
            .I(N__4266));
    Span4Mux_h I__766 (
            .O(N__4269),
            .I(N__4262));
    Span4Mux_h I__765 (
            .O(N__4266),
            .I(N__4259));
    InMux I__764 (
            .O(N__4265),
            .I(N__4256));
    Odrv4 I__763 (
            .O(N__4262),
            .I(N_80));
    Odrv4 I__762 (
            .O(N__4259),
            .I(N_80));
    LocalMux I__761 (
            .O(N__4256),
            .I(N_80));
    IoInMux I__760 (
            .O(N__4249),
            .I(N__4246));
    LocalMux I__759 (
            .O(N__4246),
            .I(N__4243));
    IoSpan4Mux I__758 (
            .O(N__4243),
            .I(N__4240));
    IoSpan4Mux I__757 (
            .O(N__4240),
            .I(N__4237));
    Span4Mux_s0_v I__756 (
            .O(N__4237),
            .I(N__4234));
    Sp12to4 I__755 (
            .O(N__4234),
            .I(N__4231));
    Span12Mux_v I__754 (
            .O(N__4231),
            .I(N__4228));
    Odrv12 I__753 (
            .O(N__4228),
            .I(N_52_i));
    InMux I__752 (
            .O(N__4225),
            .I(N__4221));
    InMux I__751 (
            .O(N__4224),
            .I(N__4218));
    LocalMux I__750 (
            .O(N__4221),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__749 (
            .O(N__4218),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    InMux I__748 (
            .O(N__4213),
            .I(N__4206));
    InMux I__747 (
            .O(N__4212),
            .I(N__4197));
    InMux I__746 (
            .O(N__4211),
            .I(N__4197));
    InMux I__745 (
            .O(N__4210),
            .I(N__4197));
    InMux I__744 (
            .O(N__4209),
            .I(N__4197));
    LocalMux I__743 (
            .O(N__4206),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__742 (
            .O(N__4197),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    InMux I__741 (
            .O(N__4192),
            .I(N__4185));
    InMux I__740 (
            .O(N__4191),
            .I(N__4176));
    InMux I__739 (
            .O(N__4190),
            .I(N__4176));
    InMux I__738 (
            .O(N__4189),
            .I(N__4176));
    InMux I__737 (
            .O(N__4188),
            .I(N__4176));
    LocalMux I__736 (
            .O(N__4185),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__735 (
            .O(N__4176),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    InMux I__734 (
            .O(N__4171),
            .I(N__4166));
    InMux I__733 (
            .O(N__4170),
            .I(N__4161));
    InMux I__732 (
            .O(N__4169),
            .I(N__4161));
    LocalMux I__731 (
            .O(N__4166),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    LocalMux I__730 (
            .O(N__4161),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    CEMux I__729 (
            .O(N__4156),
            .I(N__4153));
    LocalMux I__728 (
            .O(N__4153),
            .I(\U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en ));
    IoInMux I__727 (
            .O(N__4150),
            .I(N__4147));
    LocalMux I__726 (
            .O(N__4147),
            .I(N__4144));
    IoSpan4Mux I__725 (
            .O(N__4144),
            .I(N__4141));
    Span4Mux_s2_v I__724 (
            .O(N__4141),
            .I(N__4138));
    Span4Mux_v I__723 (
            .O(N__4138),
            .I(N__4135));
    Sp12to4 I__722 (
            .O(N__4135),
            .I(N__4131));
    CascadeMux I__721 (
            .O(N__4134),
            .I(N__4128));
    Span12Mux_v I__720 (
            .O(N__4131),
            .I(N__4125));
    InMux I__719 (
            .O(N__4128),
            .I(N__4122));
    Odrv12 I__718 (
            .O(N__4125),
            .I(ROMENn_c));
    LocalMux I__717 (
            .O(N__4122),
            .I(ROMENn_c));
    CascadeMux I__716 (
            .O(N__4117),
            .I(N__4113));
    InMux I__715 (
            .O(N__4116),
            .I(N__4110));
    InMux I__714 (
            .O(N__4113),
            .I(N__4107));
    LocalMux I__713 (
            .O(N__4110),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__712 (
            .O(N__4107),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__711 (
            .O(N__4102),
            .I(N__4099));
    LocalMux I__710 (
            .O(N__4099),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_0 ));
    InMux I__709 (
            .O(N__4096),
            .I(N__4091));
    InMux I__708 (
            .O(N__4095),
            .I(N__4088));
    InMux I__707 (
            .O(N__4094),
            .I(N__4085));
    LocalMux I__706 (
            .O(N__4091),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__705 (
            .O(N__4088),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__704 (
            .O(N__4085),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    InMux I__703 (
            .O(N__4078),
            .I(N__4072));
    InMux I__702 (
            .O(N__4077),
            .I(N__4068));
    InMux I__701 (
            .O(N__4076),
            .I(N__4065));
    InMux I__700 (
            .O(N__4075),
            .I(N__4062));
    LocalMux I__699 (
            .O(N__4072),
            .I(N__4059));
    InMux I__698 (
            .O(N__4071),
            .I(N__4056));
    LocalMux I__697 (
            .O(N__4068),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__696 (
            .O(N__4065),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__695 (
            .O(N__4062),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    Odrv4 I__694 (
            .O(N__4059),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__693 (
            .O(N__4056),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    CascadeMux I__692 (
            .O(N__4045),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_ ));
    CascadeMux I__691 (
            .O(N__4042),
            .I(N__4039));
    InMux I__690 (
            .O(N__4039),
            .I(N__4031));
    InMux I__689 (
            .O(N__4038),
            .I(N__4028));
    InMux I__688 (
            .O(N__4037),
            .I(N__4025));
    InMux I__687 (
            .O(N__4036),
            .I(N__4022));
    InMux I__686 (
            .O(N__4035),
            .I(N__4017));
    InMux I__685 (
            .O(N__4034),
            .I(N__4017));
    LocalMux I__684 (
            .O(N__4031),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__683 (
            .O(N__4028),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__682 (
            .O(N__4025),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__681 (
            .O(N__4022),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__680 (
            .O(N__4017),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__679 (
            .O(N__4006),
            .I(\U409_TRANSFER_ACK.N_54_4_cascade_ ));
    InMux I__678 (
            .O(N__4003),
            .I(N__4000));
    LocalMux I__677 (
            .O(N__4000),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_5 ));
    CascadeMux I__676 (
            .O(N__3997),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_5_cascade_ ));
    InMux I__675 (
            .O(N__3994),
            .I(N__3991));
    LocalMux I__674 (
            .O(N__3991),
            .I(N__3988));
    Odrv4 I__673 (
            .O(N__3988),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out ));
    CascadeMux I__672 (
            .O(N__3985),
            .I(N__3982));
    InMux I__671 (
            .O(N__3982),
            .I(N__3979));
    LocalMux I__670 (
            .O(N__3979),
            .I(N__3974));
    InMux I__669 (
            .O(N__3978),
            .I(N__3971));
    InMux I__668 (
            .O(N__3977),
            .I(N__3968));
    Odrv4 I__667 (
            .O(N__3974),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    LocalMux I__666 (
            .O(N__3971),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    LocalMux I__665 (
            .O(N__3968),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    CascadeMux I__664 (
            .O(N__3961),
            .I(N__3955));
    InMux I__663 (
            .O(N__3960),
            .I(N__3951));
    InMux I__662 (
            .O(N__3959),
            .I(N__3948));
    InMux I__661 (
            .O(N__3958),
            .I(N__3945));
    InMux I__660 (
            .O(N__3955),
            .I(N__3940));
    InMux I__659 (
            .O(N__3954),
            .I(N__3940));
    LocalMux I__658 (
            .O(N__3951),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__657 (
            .O(N__3948),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__656 (
            .O(N__3945),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__655 (
            .O(N__3940),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    CascadeMux I__654 (
            .O(N__3931),
            .I(N__3928));
    InMux I__653 (
            .O(N__3928),
            .I(N__3921));
    InMux I__652 (
            .O(N__3927),
            .I(N__3918));
    InMux I__651 (
            .O(N__3926),
            .I(N__3915));
    InMux I__650 (
            .O(N__3925),
            .I(N__3910));
    InMux I__649 (
            .O(N__3924),
            .I(N__3910));
    LocalMux I__648 (
            .O(N__3921),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__647 (
            .O(N__3918),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__646 (
            .O(N__3915),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__645 (
            .O(N__3910),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    InMux I__644 (
            .O(N__3901),
            .I(N__3896));
    InMux I__643 (
            .O(N__3900),
            .I(N__3888));
    InMux I__642 (
            .O(N__3899),
            .I(N__3885));
    LocalMux I__641 (
            .O(N__3896),
            .I(N__3882));
    InMux I__640 (
            .O(N__3895),
            .I(N__3879));
    InMux I__639 (
            .O(N__3894),
            .I(N__3876));
    InMux I__638 (
            .O(N__3893),
            .I(N__3869));
    InMux I__637 (
            .O(N__3892),
            .I(N__3869));
    InMux I__636 (
            .O(N__3891),
            .I(N__3869));
    LocalMux I__635 (
            .O(N__3888),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__634 (
            .O(N__3885),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    Odrv4 I__633 (
            .O(N__3882),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__632 (
            .O(N__3879),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__631 (
            .O(N__3876),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__630 (
            .O(N__3869),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    CascadeMux I__629 (
            .O(N__3856),
            .I(N__3853));
    InMux I__628 (
            .O(N__3853),
            .I(N__3847));
    CascadeMux I__627 (
            .O(N__3852),
            .I(N__3843));
    InMux I__626 (
            .O(N__3851),
            .I(N__3838));
    InMux I__625 (
            .O(N__3850),
            .I(N__3838));
    LocalMux I__624 (
            .O(N__3847),
            .I(N__3835));
    InMux I__623 (
            .O(N__3846),
            .I(N__3830));
    InMux I__622 (
            .O(N__3843),
            .I(N__3830));
    LocalMux I__621 (
            .O(N__3838),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    Odrv4 I__620 (
            .O(N__3835),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__619 (
            .O(N__3830),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    InMux I__618 (
            .O(N__3823),
            .I(N__3820));
    LocalMux I__617 (
            .O(N__3820),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a3_0_1_0 ));
    CascadeMux I__616 (
            .O(N__3817),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a3_0_1_0_cascade_ ));
    InMux I__615 (
            .O(N__3814),
            .I(N__3810));
    InMux I__614 (
            .O(N__3813),
            .I(N__3807));
    LocalMux I__613 (
            .O(N__3810),
            .I(\U409_TRANSFER_ACK.N_54_4 ));
    LocalMux I__612 (
            .O(N__3807),
            .I(\U409_TRANSFER_ACK.N_54_4 ));
    InMux I__611 (
            .O(N__3802),
            .I(N__3799));
    LocalMux I__610 (
            .O(N__3799),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0Z0Z_0 ));
    CascadeMux I__609 (
            .O(N__3796),
            .I(N__3792));
    InMux I__608 (
            .O(N__3795),
            .I(N__3787));
    InMux I__607 (
            .O(N__3792),
            .I(N__3781));
    InMux I__606 (
            .O(N__3791),
            .I(N__3781));
    InMux I__605 (
            .O(N__3790),
            .I(N__3778));
    LocalMux I__604 (
            .O(N__3787),
            .I(N__3775));
    InMux I__603 (
            .O(N__3786),
            .I(N__3772));
    LocalMux I__602 (
            .O(N__3781),
            .I(N__3769));
    LocalMux I__601 (
            .O(N__3778),
            .I(N__3766));
    Span4Mux_v I__600 (
            .O(N__3775),
            .I(N__3763));
    LocalMux I__599 (
            .O(N__3772),
            .I(N__3760));
    Span4Mux_v I__598 (
            .O(N__3769),
            .I(N__3757));
    Span4Mux_v I__597 (
            .O(N__3766),
            .I(N__3754));
    Sp12to4 I__596 (
            .O(N__3763),
            .I(N__3749));
    Span12Mux_v I__595 (
            .O(N__3760),
            .I(N__3749));
    Span4Mux_h I__594 (
            .O(N__3757),
            .I(N__3746));
    Span4Mux_h I__593 (
            .O(N__3754),
            .I(N__3743));
    Odrv12 I__592 (
            .O(N__3749),
            .I(A_c_23));
    Odrv4 I__591 (
            .O(N__3746),
            .I(A_c_23));
    Odrv4 I__590 (
            .O(N__3743),
            .I(A_c_23));
    InMux I__589 (
            .O(N__3736),
            .I(N__3733));
    LocalMux I__588 (
            .O(N__3733),
            .I(\U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3Z0Z_4 ));
    InMux I__587 (
            .O(N__3730),
            .I(N__3727));
    LocalMux I__586 (
            .O(N__3727),
            .I(N__3723));
    InMux I__585 (
            .O(N__3726),
            .I(N__3720));
    Odrv4 I__584 (
            .O(N__3723),
            .I(\U409_ADDRESS_DECODE.N_16_i ));
    LocalMux I__583 (
            .O(N__3720),
            .I(\U409_ADDRESS_DECODE.N_16_i ));
    CascadeMux I__582 (
            .O(N__3715),
            .I(un1_RAMSPACEn_i_i_a3_cascade_));
    IoInMux I__581 (
            .O(N__3712),
            .I(N__3709));
    LocalMux I__580 (
            .O(N__3709),
            .I(N__3706));
    Span4Mux_s1_v I__579 (
            .O(N__3706),
            .I(N__3703));
    Sp12to4 I__578 (
            .O(N__3703),
            .I(N__3700));
    Span12Mux_h I__577 (
            .O(N__3700),
            .I(N__3697));
    Span12Mux_v I__576 (
            .O(N__3697),
            .I(N__3694));
    Odrv12 I__575 (
            .O(N__3694),
            .I(N_11_i));
    InMux I__574 (
            .O(N__3691),
            .I(N__3687));
    InMux I__573 (
            .O(N__3690),
            .I(N__3684));
    LocalMux I__572 (
            .O(N__3687),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    LocalMux I__571 (
            .O(N__3684),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    InMux I__570 (
            .O(N__3679),
            .I(N__3675));
    InMux I__569 (
            .O(N__3678),
            .I(N__3672));
    LocalMux I__568 (
            .O(N__3675),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    LocalMux I__567 (
            .O(N__3672),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    CascadeMux I__566 (
            .O(N__3667),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ));
    CascadeMux I__565 (
            .O(N__3664),
            .I(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ));
    IoInMux I__564 (
            .O(N__3661),
            .I(N__3658));
    LocalMux I__563 (
            .O(N__3658),
            .I(N__3655));
    Span4Mux_s1_v I__562 (
            .O(N__3655),
            .I(N__3652));
    Span4Mux_v I__561 (
            .O(N__3652),
            .I(N__3649));
    Sp12to4 I__560 (
            .O(N__3649),
            .I(N__3646));
    Span12Mux_s10_h I__559 (
            .O(N__3646),
            .I(N__3643));
    Span12Mux_v I__558 (
            .O(N__3643),
            .I(N__3638));
    InMux I__557 (
            .O(N__3642),
            .I(N__3633));
    InMux I__556 (
            .O(N__3641),
            .I(N__3633));
    Odrv12 I__555 (
            .O(N__3638),
            .I(TACK_OUTn));
    LocalMux I__554 (
            .O(N__3633),
            .I(TACK_OUTn));
    CascadeMux I__553 (
            .O(N__3628),
            .I(N__3624));
    InMux I__552 (
            .O(N__3627),
            .I(N__3621));
    InMux I__551 (
            .O(N__3624),
            .I(N__3618));
    LocalMux I__550 (
            .O(N__3621),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_6 ));
    LocalMux I__549 (
            .O(N__3618),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_6 ));
    InMux I__548 (
            .O(N__3613),
            .I(N__3610));
    LocalMux I__547 (
            .O(N__3610),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3 ));
    InMux I__546 (
            .O(N__3607),
            .I(N__3600));
    InMux I__545 (
            .O(N__3606),
            .I(N__3597));
    InMux I__544 (
            .O(N__3605),
            .I(N__3594));
    InMux I__543 (
            .O(N__3604),
            .I(N__3591));
    InMux I__542 (
            .O(N__3603),
            .I(N__3588));
    LocalMux I__541 (
            .O(N__3600),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__540 (
            .O(N__3597),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__539 (
            .O(N__3594),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__538 (
            .O(N__3591),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__537 (
            .O(N__3588),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    InMux I__536 (
            .O(N__3577),
            .I(N__3572));
    InMux I__535 (
            .O(N__3576),
            .I(N__3568));
    InMux I__534 (
            .O(N__3575),
            .I(N__3565));
    LocalMux I__533 (
            .O(N__3572),
            .I(N__3562));
    InMux I__532 (
            .O(N__3571),
            .I(N__3559));
    LocalMux I__531 (
            .O(N__3568),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__530 (
            .O(N__3565),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    Odrv4 I__529 (
            .O(N__3562),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__528 (
            .O(N__3559),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    CascadeMux I__527 (
            .O(N__3550),
            .I(N__3547));
    InMux I__526 (
            .O(N__3547),
            .I(N__3544));
    LocalMux I__525 (
            .O(N__3544),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    CascadeMux I__524 (
            .O(N__3541),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    InMux I__523 (
            .O(N__3538),
            .I(N__3534));
    InMux I__522 (
            .O(N__3537),
            .I(N__3531));
    LocalMux I__521 (
            .O(N__3534),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    LocalMux I__520 (
            .O(N__3531),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    CascadeMux I__519 (
            .O(N__3526),
            .I(N__3522));
    InMux I__518 (
            .O(N__3525),
            .I(N__3519));
    InMux I__517 (
            .O(N__3522),
            .I(N__3516));
    LocalMux I__516 (
            .O(N__3519),
            .I(N__3511));
    LocalMux I__515 (
            .O(N__3516),
            .I(N__3511));
    Span4Mux_v I__514 (
            .O(N__3511),
            .I(N__3508));
    Odrv4 I__513 (
            .O(N__3508),
            .I(\U409_CIA.N_89 ));
    InMux I__512 (
            .O(N__3505),
            .I(N__3497));
    InMux I__511 (
            .O(N__3504),
            .I(N__3497));
    InMux I__510 (
            .O(N__3503),
            .I(N__3494));
    CascadeMux I__509 (
            .O(N__3502),
            .I(N__3490));
    LocalMux I__508 (
            .O(N__3497),
            .I(N__3487));
    LocalMux I__507 (
            .O(N__3494),
            .I(N__3484));
    InMux I__506 (
            .O(N__3493),
            .I(N__3479));
    InMux I__505 (
            .O(N__3490),
            .I(N__3479));
    Span4Mux_v I__504 (
            .O(N__3487),
            .I(N__3476));
    Span4Mux_h I__503 (
            .O(N__3484),
            .I(N__3471));
    LocalMux I__502 (
            .O(N__3479),
            .I(N__3468));
    Span4Mux_v I__501 (
            .O(N__3476),
            .I(N__3465));
    InMux I__500 (
            .O(N__3475),
            .I(N__3460));
    InMux I__499 (
            .O(N__3474),
            .I(N__3460));
    Span4Mux_h I__498 (
            .O(N__3471),
            .I(N__3455));
    Span4Mux_v I__497 (
            .O(N__3468),
            .I(N__3455));
    Span4Mux_v I__496 (
            .O(N__3465),
            .I(N__3452));
    LocalMux I__495 (
            .O(N__3460),
            .I(N__3449));
    Span4Mux_v I__494 (
            .O(N__3455),
            .I(N__3446));
    Span4Mux_h I__493 (
            .O(N__3452),
            .I(N__3443));
    Sp12to4 I__492 (
            .O(N__3449),
            .I(N__3440));
    Span4Mux_v I__491 (
            .O(N__3446),
            .I(N__3437));
    Sp12to4 I__490 (
            .O(N__3443),
            .I(N__3432));
    Span12Mux_v I__489 (
            .O(N__3440),
            .I(N__3432));
    Span4Mux_h I__488 (
            .O(N__3437),
            .I(N__3429));
    Odrv12 I__487 (
            .O(N__3432),
            .I(A_c_22));
    Odrv4 I__486 (
            .O(N__3429),
            .I(A_c_22));
    InMux I__485 (
            .O(N__3424),
            .I(N__3421));
    LocalMux I__484 (
            .O(N__3421),
            .I(N__3418));
    Span4Mux_v I__483 (
            .O(N__3418),
            .I(N__3414));
    InMux I__482 (
            .O(N__3417),
            .I(N__3411));
    Span4Mux_h I__481 (
            .O(N__3414),
            .I(N__3408));
    LocalMux I__480 (
            .O(N__3411),
            .I(N__3405));
    Sp12to4 I__479 (
            .O(N__3408),
            .I(N__3400));
    Span12Mux_v I__478 (
            .O(N__3405),
            .I(N__3400));
    Span12Mux_v I__477 (
            .O(N__3400),
            .I(N__3397));
    Span12Mux_h I__476 (
            .O(N__3397),
            .I(N__3394));
    Odrv12 I__475 (
            .O(N__3394),
            .I(OVL_c));
    CascadeMux I__474 (
            .O(N__3391),
            .I(\U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3Z0Z_4_cascade_ ));
    IoInMux I__473 (
            .O(N__3388),
            .I(N__3385));
    LocalMux I__472 (
            .O(N__3385),
            .I(N__3382));
    Span4Mux_s2_v I__471 (
            .O(N__3382),
            .I(N__3379));
    Span4Mux_h I__470 (
            .O(N__3379),
            .I(N__3376));
    Sp12to4 I__469 (
            .O(N__3376),
            .I(N__3373));
    Span12Mux_v I__468 (
            .O(N__3373),
            .I(N__3370));
    Odrv12 I__467 (
            .O(N__3370),
            .I(N_53_i));
    InMux I__466 (
            .O(N__3367),
            .I(N__3364));
    LocalMux I__465 (
            .O(N__3364),
            .I(N__3361));
    Odrv4 I__464 (
            .O(N__3361),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_17 ));
    InMux I__463 (
            .O(N__3358),
            .I(N__3355));
    LocalMux I__462 (
            .O(N__3355),
            .I(N__3352));
    Span4Mux_v I__461 (
            .O(N__3352),
            .I(N__3349));
    Odrv4 I__460 (
            .O(N__3349),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_16 ));
    InMux I__459 (
            .O(N__3346),
            .I(N__3339));
    InMux I__458 (
            .O(N__3345),
            .I(N__3339));
    InMux I__457 (
            .O(N__3344),
            .I(N__3336));
    LocalMux I__456 (
            .O(N__3339),
            .I(N__3331));
    LocalMux I__455 (
            .O(N__3336),
            .I(N__3331));
    Span12Mux_h I__454 (
            .O(N__3331),
            .I(N__3328));
    Span12Mux_v I__453 (
            .O(N__3328),
            .I(N__3325));
    Odrv12 I__452 (
            .O(N__3325),
            .I(TM_c_0));
    InMux I__451 (
            .O(N__3322),
            .I(N__3316));
    InMux I__450 (
            .O(N__3321),
            .I(N__3316));
    LocalMux I__449 (
            .O(N__3316),
            .I(N__3312));
    InMux I__448 (
            .O(N__3315),
            .I(N__3309));
    Span4Mux_h I__447 (
            .O(N__3312),
            .I(N__3304));
    LocalMux I__446 (
            .O(N__3309),
            .I(N__3304));
    Span4Mux_h I__445 (
            .O(N__3304),
            .I(N__3301));
    Sp12to4 I__444 (
            .O(N__3301),
            .I(N__3298));
    Odrv12 I__443 (
            .O(N__3298),
            .I(TM_c_1));
    IoInMux I__442 (
            .O(N__3295),
            .I(N__3292));
    LocalMux I__441 (
            .O(N__3292),
            .I(N__3289));
    IoSpan4Mux I__440 (
            .O(N__3289),
            .I(N__3286));
    Span4Mux_s0_v I__439 (
            .O(N__3286),
            .I(N__3283));
    Sp12to4 I__438 (
            .O(N__3283),
            .I(N__3280));
    Span12Mux_v I__437 (
            .O(N__3280),
            .I(N__3277));
    Odrv12 I__436 (
            .O(N__3277),
            .I(PORTSIZE_i_a2));
    InMux I__435 (
            .O(N__3274),
            .I(N__3271));
    LocalMux I__434 (
            .O(N__3271),
            .I(N__3268));
    Span4Mux_v I__433 (
            .O(N__3268),
            .I(N__3265));
    Span4Mux_v I__432 (
            .O(N__3265),
            .I(N__3262));
    Odrv4 I__431 (
            .O(N__3262),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_12 ));
    InMux I__430 (
            .O(N__3259),
            .I(N__3256));
    LocalMux I__429 (
            .O(N__3256),
            .I(N__3253));
    Span4Mux_h I__428 (
            .O(N__3253),
            .I(N__3249));
    InMux I__427 (
            .O(N__3252),
            .I(N__3246));
    Odrv4 I__426 (
            .O(N__3249),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    LocalMux I__425 (
            .O(N__3246),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    InMux I__424 (
            .O(N__3241),
            .I(N__3235));
    InMux I__423 (
            .O(N__3240),
            .I(N__3235));
    LocalMux I__422 (
            .O(N__3235),
            .I(N__3231));
    InMux I__421 (
            .O(N__3234),
            .I(N__3228));
    Span4Mux_v I__420 (
            .O(N__3231),
            .I(N__3225));
    LocalMux I__419 (
            .O(N__3228),
            .I(N__3222));
    Odrv4 I__418 (
            .O(N__3225),
            .I(U409_CIA_PORTSIZE_i_a2_0_3));
    Odrv12 I__417 (
            .O(N__3222),
            .I(U409_CIA_PORTSIZE_i_a2_0_3));
    CascadeMux I__416 (
            .O(N__3217),
            .I(N__3214));
    InMux I__415 (
            .O(N__3214),
            .I(N__3209));
    InMux I__414 (
            .O(N__3213),
            .I(N__3206));
    InMux I__413 (
            .O(N__3212),
            .I(N__3203));
    LocalMux I__412 (
            .O(N__3209),
            .I(N__3199));
    LocalMux I__411 (
            .O(N__3206),
            .I(N__3194));
    LocalMux I__410 (
            .O(N__3203),
            .I(N__3194));
    InMux I__409 (
            .O(N__3202),
            .I(N__3191));
    Span4Mux_v I__408 (
            .O(N__3199),
            .I(N__3186));
    Span4Mux_v I__407 (
            .O(N__3194),
            .I(N__3186));
    LocalMux I__406 (
            .O(N__3191),
            .I(N__3183));
    Sp12to4 I__405 (
            .O(N__3186),
            .I(N__3180));
    Span4Mux_h I__404 (
            .O(N__3183),
            .I(N__3177));
    Span12Mux_h I__403 (
            .O(N__3180),
            .I(N__3172));
    Sp12to4 I__402 (
            .O(N__3177),
            .I(N__3172));
    Span12Mux_v I__401 (
            .O(N__3172),
            .I(N__3169));
    Odrv12 I__400 (
            .O(N__3169),
            .I(A_c_19));
    CascadeMux I__399 (
            .O(N__3166),
            .I(N__3162));
    InMux I__398 (
            .O(N__3165),
            .I(N__3158));
    InMux I__397 (
            .O(N__3162),
            .I(N__3155));
    InMux I__396 (
            .O(N__3161),
            .I(N__3152));
    LocalMux I__395 (
            .O(N__3158),
            .I(N__3145));
    LocalMux I__394 (
            .O(N__3155),
            .I(N__3145));
    LocalMux I__393 (
            .O(N__3152),
            .I(N__3145));
    Span4Mux_v I__392 (
            .O(N__3145),
            .I(N__3142));
    Sp12to4 I__391 (
            .O(N__3142),
            .I(N__3139));
    Span12Mux_h I__390 (
            .O(N__3139),
            .I(N__3136));
    Span12Mux_v I__389 (
            .O(N__3136),
            .I(N__3133));
    Odrv12 I__388 (
            .O(N__3133),
            .I(A_c_18));
    CascadeMux I__387 (
            .O(N__3130),
            .I(N__3127));
    InMux I__386 (
            .O(N__3127),
            .I(N__3124));
    LocalMux I__385 (
            .O(N__3124),
            .I(N__3120));
    InMux I__384 (
            .O(N__3123),
            .I(N__3117));
    Span4Mux_h I__383 (
            .O(N__3120),
            .I(N__3112));
    LocalMux I__382 (
            .O(N__3117),
            .I(N__3112));
    Span4Mux_v I__381 (
            .O(N__3112),
            .I(N__3109));
    Span4Mux_h I__380 (
            .O(N__3109),
            .I(N__3106));
    Sp12to4 I__379 (
            .O(N__3106),
            .I(N__3103));
    Odrv12 I__378 (
            .O(N__3103),
            .I(TT_c_0));
    InMux I__377 (
            .O(N__3100),
            .I(N__3094));
    InMux I__376 (
            .O(N__3099),
            .I(N__3094));
    LocalMux I__375 (
            .O(N__3094),
            .I(N__3090));
    InMux I__374 (
            .O(N__3093),
            .I(N__3087));
    Span4Mux_h I__373 (
            .O(N__3090),
            .I(N__3082));
    LocalMux I__372 (
            .O(N__3087),
            .I(N__3082));
    Span4Mux_v I__371 (
            .O(N__3082),
            .I(N__3079));
    Span4Mux_v I__370 (
            .O(N__3079),
            .I(N__3076));
    Span4Mux_h I__369 (
            .O(N__3076),
            .I(N__3073));
    Odrv4 I__368 (
            .O(N__3073),
            .I(A_c_26));
    InMux I__367 (
            .O(N__3070),
            .I(N__3064));
    InMux I__366 (
            .O(N__3069),
            .I(N__3064));
    LocalMux I__365 (
            .O(N__3064),
            .I(N__3061));
    Span4Mux_v I__364 (
            .O(N__3061),
            .I(N__3058));
    Span4Mux_h I__363 (
            .O(N__3058),
            .I(N__3055));
    Sp12to4 I__362 (
            .O(N__3055),
            .I(N__3052));
    Odrv12 I__361 (
            .O(N__3052),
            .I(TT_c_1));
    CascadeMux I__360 (
            .O(N__3049),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_11_cascade_ ));
    InMux I__359 (
            .O(N__3046),
            .I(N__3043));
    LocalMux I__358 (
            .O(N__3043),
            .I(N__3040));
    Odrv4 I__357 (
            .O(N__3040),
            .I(\U409_TRANSFER_ACK.N_17 ));
    InMux I__356 (
            .O(N__3037),
            .I(N__3033));
    InMux I__355 (
            .O(N__3036),
            .I(N__3030));
    LocalMux I__354 (
            .O(N__3033),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_4 ));
    LocalMux I__353 (
            .O(N__3030),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_4 ));
    CascadeMux I__352 (
            .O(N__3025),
            .I(N__3021));
    InMux I__351 (
            .O(N__3024),
            .I(N__3018));
    InMux I__350 (
            .O(N__3021),
            .I(N__3015));
    LocalMux I__349 (
            .O(N__3018),
            .I(N__3010));
    LocalMux I__348 (
            .O(N__3015),
            .I(N__3010));
    Odrv12 I__347 (
            .O(N__3010),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_11 ));
    InMux I__346 (
            .O(N__3007),
            .I(N__3004));
    LocalMux I__345 (
            .O(N__3004),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_14 ));
    InMux I__344 (
            .O(N__3001),
            .I(N__2998));
    LocalMux I__343 (
            .O(N__2998),
            .I(N__2994));
    InMux I__342 (
            .O(N__2997),
            .I(N__2991));
    Span4Mux_v I__341 (
            .O(N__2994),
            .I(N__2988));
    LocalMux I__340 (
            .O(N__2991),
            .I(N__2985));
    Span4Mux_h I__339 (
            .O(N__2988),
            .I(N__2982));
    Span4Mux_v I__338 (
            .O(N__2985),
            .I(N__2979));
    Odrv4 I__337 (
            .O(N__2982),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_10 ));
    Odrv4 I__336 (
            .O(N__2979),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_10 ));
    InMux I__335 (
            .O(N__2974),
            .I(N__2971));
    LocalMux I__334 (
            .O(N__2971),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1 ));
    InMux I__333 (
            .O(N__2968),
            .I(N__2965));
    LocalMux I__332 (
            .O(N__2965),
            .I(N__2961));
    InMux I__331 (
            .O(N__2964),
            .I(N__2958));
    Span4Mux_v I__330 (
            .O(N__2961),
            .I(N__2953));
    LocalMux I__329 (
            .O(N__2958),
            .I(N__2953));
    Span4Mux_h I__328 (
            .O(N__2953),
            .I(N__2950));
    Span4Mux_v I__327 (
            .O(N__2950),
            .I(N__2947));
    Odrv4 I__326 (
            .O(N__2947),
            .I(A_c_31));
    CascadeMux I__325 (
            .O(N__2944),
            .I(N__2940));
    CascadeMux I__324 (
            .O(N__2943),
            .I(N__2937));
    InMux I__323 (
            .O(N__2940),
            .I(N__2934));
    InMux I__322 (
            .O(N__2937),
            .I(N__2931));
    LocalMux I__321 (
            .O(N__2934),
            .I(N__2926));
    LocalMux I__320 (
            .O(N__2931),
            .I(N__2926));
    Span4Mux_v I__319 (
            .O(N__2926),
            .I(N__2923));
    Span4Mux_v I__318 (
            .O(N__2923),
            .I(N__2920));
    Span4Mux_h I__317 (
            .O(N__2920),
            .I(N__2917));
    Odrv4 I__316 (
            .O(N__2917),
            .I(A_c_24));
    InMux I__315 (
            .O(N__2914),
            .I(N__2910));
    InMux I__314 (
            .O(N__2913),
            .I(N__2907));
    LocalMux I__313 (
            .O(N__2910),
            .I(N__2902));
    LocalMux I__312 (
            .O(N__2907),
            .I(N__2902));
    Span4Mux_v I__311 (
            .O(N__2902),
            .I(N__2899));
    Span4Mux_h I__310 (
            .O(N__2899),
            .I(N__2896));
    Odrv4 I__309 (
            .O(N__2896),
            .I(A_c_25));
    InMux I__308 (
            .O(N__2893),
            .I(N__2890));
    LocalMux I__307 (
            .O(N__2890),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_3 ));
    InMux I__306 (
            .O(N__2887),
            .I(N__2884));
    LocalMux I__305 (
            .O(N__2884),
            .I(N__2880));
    InMux I__304 (
            .O(N__2883),
            .I(N__2877));
    Span4Mux_h I__303 (
            .O(N__2880),
            .I(N__2872));
    LocalMux I__302 (
            .O(N__2877),
            .I(N__2872));
    Span4Mux_v I__301 (
            .O(N__2872),
            .I(N__2869));
    Span4Mux_h I__300 (
            .O(N__2869),
            .I(N__2866));
    Odrv4 I__299 (
            .O(N__2866),
            .I(A_c_30));
    CascadeMux I__298 (
            .O(N__2863),
            .I(N__2860));
    InMux I__297 (
            .O(N__2860),
            .I(N__2854));
    InMux I__296 (
            .O(N__2859),
            .I(N__2854));
    LocalMux I__295 (
            .O(N__2854),
            .I(N__2851));
    Span4Mux_h I__294 (
            .O(N__2851),
            .I(N__2848));
    Span4Mux_v I__293 (
            .O(N__2848),
            .I(N__2845));
    Span4Mux_v I__292 (
            .O(N__2845),
            .I(N__2842));
    Odrv4 I__291 (
            .O(N__2842),
            .I(A_c_28));
    InMux I__290 (
            .O(N__2839),
            .I(N__2833));
    InMux I__289 (
            .O(N__2838),
            .I(N__2833));
    LocalMux I__288 (
            .O(N__2833),
            .I(N__2830));
    Sp12to4 I__287 (
            .O(N__2830),
            .I(N__2827));
    Span12Mux_v I__286 (
            .O(N__2827),
            .I(N__2824));
    Odrv12 I__285 (
            .O(N__2824),
            .I(A_c_29));
    CascadeMux I__284 (
            .O(N__2821),
            .I(N__2817));
    InMux I__283 (
            .O(N__2820),
            .I(N__2814));
    InMux I__282 (
            .O(N__2817),
            .I(N__2811));
    LocalMux I__281 (
            .O(N__2814),
            .I(N__2806));
    LocalMux I__280 (
            .O(N__2811),
            .I(N__2806));
    Odrv12 I__279 (
            .O(N__2806),
            .I(A_c_27));
    InMux I__278 (
            .O(N__2803),
            .I(N__2800));
    LocalMux I__277 (
            .O(N__2800),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4 ));
    InMux I__276 (
            .O(N__2797),
            .I(N__2794));
    LocalMux I__275 (
            .O(N__2794),
            .I(N__2790));
    CascadeMux I__274 (
            .O(N__2793),
            .I(N__2787));
    Span4Mux_v I__273 (
            .O(N__2790),
            .I(N__2784));
    InMux I__272 (
            .O(N__2787),
            .I(N__2781));
    Sp12to4 I__271 (
            .O(N__2784),
            .I(N__2776));
    LocalMux I__270 (
            .O(N__2781),
            .I(N__2776));
    Odrv12 I__269 (
            .O(N__2776),
            .I(A_c_20));
    CascadeMux I__268 (
            .O(N__2773),
            .I(\U409_TRANSFER_ACK.N_41_cascade_ ));
    InMux I__267 (
            .O(N__2770),
            .I(N__2767));
    LocalMux I__266 (
            .O(N__2767),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3Z0Z_2 ));
    InMux I__265 (
            .O(N__2764),
            .I(N__2761));
    LocalMux I__264 (
            .O(N__2761),
            .I(N__2758));
    Span4Mux_v I__263 (
            .O(N__2758),
            .I(N__2755));
    Sp12to4 I__262 (
            .O(N__2755),
            .I(N__2752));
    Span12Mux_s3_h I__261 (
            .O(N__2752),
            .I(N__2749));
    Span12Mux_v I__260 (
            .O(N__2749),
            .I(N__2746));
    Odrv12 I__259 (
            .O(N__2746),
            .I(A_c_16));
    InMux I__258 (
            .O(N__2743),
            .I(N__2740));
    LocalMux I__257 (
            .O(N__2740),
            .I(N__2737));
    Span4Mux_v I__256 (
            .O(N__2737),
            .I(N__2734));
    Sp12to4 I__255 (
            .O(N__2734),
            .I(N__2731));
    Span12Mux_v I__254 (
            .O(N__2731),
            .I(N__2728));
    Odrv12 I__253 (
            .O(N__2728),
            .I(A_c_17));
    ClkMux I__252 (
            .O(N__2725),
            .I(N__2677));
    ClkMux I__251 (
            .O(N__2724),
            .I(N__2677));
    ClkMux I__250 (
            .O(N__2723),
            .I(N__2677));
    ClkMux I__249 (
            .O(N__2722),
            .I(N__2677));
    ClkMux I__248 (
            .O(N__2721),
            .I(N__2677));
    ClkMux I__247 (
            .O(N__2720),
            .I(N__2677));
    ClkMux I__246 (
            .O(N__2719),
            .I(N__2677));
    ClkMux I__245 (
            .O(N__2718),
            .I(N__2677));
    ClkMux I__244 (
            .O(N__2717),
            .I(N__2677));
    ClkMux I__243 (
            .O(N__2716),
            .I(N__2677));
    ClkMux I__242 (
            .O(N__2715),
            .I(N__2677));
    ClkMux I__241 (
            .O(N__2714),
            .I(N__2677));
    ClkMux I__240 (
            .O(N__2713),
            .I(N__2677));
    ClkMux I__239 (
            .O(N__2712),
            .I(N__2677));
    ClkMux I__238 (
            .O(N__2711),
            .I(N__2677));
    ClkMux I__237 (
            .O(N__2710),
            .I(N__2677));
    GlobalMux I__236 (
            .O(N__2677),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.LASTCLK_0C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .I(N__2712));
    INV \INVU409_TRANSFER_ACK.LASTCLK_1C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .I(N__2711));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .I(N__2710));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__2713));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .I(N__2721));
    INV \INVU409_TRANSFER_ACK.ROMENnC  (
            .O(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .I(N__2717));
    INV \INVU409_TRANSFER_ACK.TACK_EN_iC  (
            .O(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .I(N__2715));
    INV \INVU409_TRANSFER_ACK.CIA_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .I(N__2714));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .I(N__2723));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .I(N__2720));
    INV \INVU409_TRANSFER_ACK.TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .I(N__2716));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .I(N__2724));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .I(N__2722));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .I(N__2719));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net ),
            .I(N__2718));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .I(N__2725));
    defparam IN_MUX_bfv_13_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_2_0_));
    defparam IN_MUX_bfv_13_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_3_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_13_3_0_));
    defparam IN_MUX_bfv_15_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_1_0_));
    defparam IN_MUX_bfv_15_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_2_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_15_2_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_12_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_CIA.PORTSIZE_i_a2_0_3_LC_1_12_5 .C_ON=1'b0;
    defparam \U409_CIA.PORTSIZE_i_a2_0_3_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.PORTSIZE_i_a2_0_3_LC_1_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.PORTSIZE_i_a2_0_3_LC_1_12_5  (
            .in0(N__2764),
            .in1(N__3790),
            .in2(N__2793),
            .in3(N__2743),
            .lcout(U409_CIA_PORTSIZE_i_a2_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_11_LC_1_14_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_11_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_11_LC_1_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_11_LC_1_14_5  (
            .in0(N__2968),
            .in1(N__2914),
            .in2(N__2944),
            .in3(N__4308),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_15_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_15_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_15_0  (
            .in0(N__2893),
            .in1(N__2964),
            .in2(N__2943),
            .in3(N__2803),
            .lcout(N_76),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_3_LC_1_15_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_3_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_3_LC_1_15_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_3_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__2887),
            .in2(_gnd_net_),
            .in3(N__2913),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_10_LC_1_16_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_10_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_10_LC_1_16_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_10_LC_1_16_0  (
            .in0(N__2883),
            .in1(N__2839),
            .in2(N__2863),
            .in3(N__2820),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_16_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_16_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_16_2  (
            .in0(N__2859),
            .in1(N__2838),
            .in2(N__2821),
            .in3(N__3093),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_0_LC_3_13_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_0_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_0_LC_3_13_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_0_LC_3_13_1  (
            .in0(N__3424),
            .in1(N__3791),
            .in2(N__3502),
            .in3(N__4336),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.N_41_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_3_13_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_3_13_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_3_13_2  (
            .in0(N__2797),
            .in1(N__2770),
            .in2(N__2773),
            .in3(N__3493),
            .lcout(\U409_TRANSFER_ACK.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_2_LC_3_13_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_2_LC_3_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_2_LC_3_13_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_2_LC_3_13_4  (
            .in0(N__4337),
            .in1(_gnd_net_),
            .in2(N__3796),
            .in3(N__3202),
            .lcout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.PORTSIZE_i_a2_0_LC_5_12_0 .C_ON=1'b0;
    defparam \U409_CIA.PORTSIZE_i_a2_0_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.PORTSIZE_i_a2_0_LC_5_12_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_CIA.PORTSIZE_i_a2_0_LC_5_12_0  (
            .in0(N__3234),
            .in1(N__3212),
            .in2(_gnd_net_),
            .in3(N__3161),
            .lcout(\U409_CIA.N_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_0_LC_5_13_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_0_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_0_LC_5_13_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_0_LC_5_13_1  (
            .in0(N__3241),
            .in1(N__3475),
            .in2(N__3130),
            .in3(N__3036),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_0_0_a2_LC_5_13_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_0_0_a2_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_0_0_a2_LC_5_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_0_0_a2_LC_5_13_6  (
            .in0(N__3474),
            .in1(N__3213),
            .in2(N__3166),
            .in3(N__3240),
            .lcout(N_80),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_2_LC_5_14_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_2_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_2_LC_5_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_2_LC_5_14_4  (
            .in0(N__3069),
            .in1(N__3099),
            .in2(N__3217),
            .in3(N__3165),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_1_LC_5_14_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_1_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_1_LC_5_14_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_1_LC_5_14_6  (
            .in0(N__4265),
            .in1(N__3123),
            .in2(N__3025),
            .in3(N__3037),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_5_14_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_5_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_5_14_7  (
            .in0(N__3100),
            .in1(N__3070),
            .in2(N__3049),
            .in3(N__2997),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_3_LC_6_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_3_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_3_LC_6_13_5 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_3_LC_6_13_5  (
            .in0(N__3315),
            .in1(N__3046),
            .in2(_gnd_net_),
            .in3(N__3344),
            .lcout(\U409_TRANSFER_ACK.N_28_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_4_LC_6_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_4_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_4_LC_6_13_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_4_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(N__5371),
            .in2(_gnd_net_),
            .in3(N__4634),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_1_LC_6_14_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_1_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_1_LC_6_14_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_1_LC_6_14_5  (
            .in0(N__3024),
            .in1(N__3007),
            .in2(_gnd_net_),
            .in3(N__3001),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_7_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_7_11_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_7_11_0  (
            .in0(N__2974),
            .in1(N__3901),
            .in2(_gnd_net_),
            .in3(N__3605),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_7_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_7_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_7_12_3  (
            .in0(N__4078),
            .in1(N__4036),
            .in2(N__3856),
            .in3(N__3577),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_7_12_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_7_12_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_7_12_6  (
            .in0(N__3367),
            .in1(N__3358),
            .in2(N__4805),
            .in3(N__3252),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un2_ROMEN_0_i_0_x3_LC_7_13_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un2_ROMEN_0_i_0_x3_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un2_ROMEN_0_i_0_x3_LC_7_13_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U409_ADDRESS_DECODE.un2_ROMEN_0_i_0_x3_LC_7_13_5  (
            .in0(N__3346),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3322),
            .lcout(\U409_ADDRESS_DECODE.N_16_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a3_0_a2_0_LC_7_13_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a3_0_a2_0_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a3_0_a2_0_LC_7_13_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a3_0_a2_0_LC_7_13_7  (
            .in0(N__3345),
            .in1(N__3321),
            .in2(N__4605),
            .in3(N__5367),
            .lcout(N_90),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.PORTSIZE_i_a2_LC_7_14_4 .C_ON=1'b0;
    defparam \U409_CIA.PORTSIZE_i_a2_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.PORTSIZE_i_a2_LC_7_14_4 .LUT_INIT=16'b0010000010000000;
    LogicCell40 \U409_CIA.PORTSIZE_i_a2_LC_7_14_4  (
            .in0(N__4372),
            .in1(N__3503),
            .in2(N__3526),
            .in3(N__4328),
            .lcout(PORTSIZE_i_a2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_8_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_8_9_3 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_8_9_3  (
            .in0(N__3274),
            .in1(N__3259),
            .in2(N__4806),
            .in3(N__3691),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net ),
            .ce(),
            .sr(N__5243));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_8_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_8_10_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_8_10_2  (
            .in0(N__3900),
            .in1(N__3576),
            .in2(_gnd_net_),
            .in3(N__3607),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__4443));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_8_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_8_10_3 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_8_10_3 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_8_10_3  (
            .in0(N__3627),
            .in1(N__3679),
            .in2(_gnd_net_),
            .in3(N__4003),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__4443));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_8_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_8_10_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_8_10_6 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_8_10_6  (
            .in0(N__4077),
            .in1(N__3978),
            .in2(N__4042),
            .in3(N__3959),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__4443));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_8_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_8_11_2 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__3927),
            .in2(N__3961),
            .in3(N__3537),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__4444));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_8_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_8_11_4 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_8_11_4  (
            .in0(N__4774),
            .in1(N__3823),
            .in2(N__3628),
            .in3(N__3814),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_8_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_8_11_5 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__3899),
            .in2(N__3541),
            .in3(N__3606),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__4444));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_8_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_8_11_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_8_11_7  (
            .in0(N__3977),
            .in1(N__4038),
            .in2(_gnd_net_),
            .in3(N__3954),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__4444));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_8_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_8_12_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_8_12_0 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_8_12_0  (
            .in0(N__3538),
            .in1(N__4096),
            .in2(N__3931),
            .in3(N__3960),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net ),
            .ce(),
            .sr(N__4439));
    defparam \U409_CIA.VMA_RNO_0_LC_8_13_3 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_8_13_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_8_13_3  (
            .in0(N__3525),
            .in1(N__3505),
            .in2(N__4392),
            .in3(N__4351),
            .lcout(\U409_CIA.VMA_3_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3_4_LC_8_13_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3_4_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3_4_LC_8_13_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3_4_LC_8_13_6  (
            .in0(N__3504),
            .in1(N__5366),
            .in2(N__4354),
            .in3(N__3417),
            .lcout(\U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3Z0Z_4 ),
            .ltout(\U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.N_53_i_LC_8_13_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.N_53_i_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.N_53_i_LC_8_13_7 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \U409_ADDRESS_DECODE.N_53_i_LC_8_13_7  (
            .in0(N__3786),
            .in1(N__3726),
            .in2(N__3391),
            .in3(N__4600),
            .lcout(N_53_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_9_0 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_9_0  (
            .in0(N__4211),
            .in1(N__5349),
            .in2(_gnd_net_),
            .in3(N__4190),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_9_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_9_9_2 .LUT_INIT=16'b1000111110011111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_9_9_2  (
            .in0(N__4210),
            .in1(N__4189),
            .in2(N__5364),
            .in3(N__4169),
            .lcout(\U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_9_4 .LUT_INIT=16'b0010000000110000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_9_4  (
            .in0(N__4212),
            .in1(N__4191),
            .in2(N__5363),
            .in3(N__4170),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_9_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_9_9_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_9_9_5  (
            .in0(N__3690),
            .in1(N__4224),
            .in2(N__4117),
            .in3(N__3678),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER6 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_9_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_9_9_6 .LUT_INIT=16'b0000000111011101;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_9_9_6  (
            .in0(N__4209),
            .in1(N__4188),
            .in2(N__3667),
            .in3(N__3641),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_9_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_9_9_7 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_9_9_7  (
            .in0(N__3642),
            .in1(_gnd_net_),
            .in2(N__3664),
            .in3(N__5348),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_9_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_9_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__4076),
            .in2(_gnd_net_),
            .in3(N__4037),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_9_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_9_10_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_9_10_5  (
            .in0(N__3895),
            .in1(N__3575),
            .in2(_gnd_net_),
            .in3(N__3604),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_9_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_9_11_0 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_9_11_0  (
            .in0(N__3924),
            .in1(N__3891),
            .in2(N__3550),
            .in3(N__3613),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_9_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_9_11_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_9_11_1  (
            .in0(N__4071),
            .in1(N__4034),
            .in2(N__3852),
            .in3(N__4094),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_9_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_9_11_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__3603),
            .in2(_gnd_net_),
            .in3(N__3571),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIG5942_7_LC_9_11_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIG5942_7_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIG5942_7_LC_9_11_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIG5942_7_LC_9_11_3  (
            .in0(N__4095),
            .in1(N__4075),
            .in2(N__4045),
            .in3(N__4035),
            .lcout(\U409_TRANSFER_ACK.N_54_4 ),
            .ltout(\U409_TRANSFER_ACK.N_54_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_9_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_9_11_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_9_11_4  (
            .in0(N__3925),
            .in1(N__3892),
            .in2(N__4006),
            .in3(N__3846),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_5 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_11_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_11_5 .LUT_INIT=16'b1111111100000101;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_11_5  (
            .in0(N__3893),
            .in1(_gnd_net_),
            .in2(N__3997),
            .in3(N__3802),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__4438));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_12_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_12_0 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_12_0  (
            .in0(N__3994),
            .in1(N__3851),
            .in2(N__3985),
            .in3(N__3958),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__4425));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIUGMJ1_5_LC_9_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIUGMJ1_5_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIUGMJ1_5_LC_9_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIUGMJ1_5_LC_9_12_2  (
            .in0(N__3926),
            .in1(N__3894),
            .in2(N__4651),
            .in3(N__3850),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a3_0_1_0 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a3_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_0_LC_9_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_0_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_0_LC_9_12_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_0_LC_9_12_3  (
            .in0(N__4778),
            .in1(_gnd_net_),
            .in2(N__3817),
            .in3(N__3813),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3_LC_9_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3_LC_9_13_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3_LC_9_13_3  (
            .in0(N__3795),
            .in1(N__3736),
            .in2(N__4604),
            .in3(N__3730),
            .lcout(un1_RAMSPACEn_i_i_a3),
            .ltout(un1_RAMSPACEn_i_i_a3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.N_11_i_LC_9_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.N_11_i_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.N_11_i_LC_9_13_4 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \U409_ADDRESS_DECODE.N_11_i_LC_9_13_4  (
            .in0(N__4387),
            .in1(N__4352),
            .in2(N__3715),
            .in3(N__4280),
            .lcout(N_11_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a3_0_a2_LC_9_13_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a3_0_a2_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a3_0_a2_LC_9_13_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a3_0_a2_LC_9_13_6  (
            .in0(N__4388),
            .in1(N__4353),
            .in2(_gnd_net_),
            .in3(N__4281),
            .lcout(),
            .ltout(un1_REGSPACEn_i_i_a3_0_a2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_7 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_7  (
            .in0(N__4471),
            .in1(N__4465),
            .in2(N__4447),
            .in3(N__5365),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.N_52_i_LC_9_14_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.N_52_i_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.N_52_i_LC_9_14_0 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U409_ADDRESS_DECODE.N_52_i_LC_9_14_0  (
            .in0(N__4393),
            .in1(N__4329),
            .in2(_gnd_net_),
            .in3(N__4282),
            .lcout(N_52_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_8_0 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_8_0  (
            .in0(N__4657),
            .in1(N__4225),
            .in2(_gnd_net_),
            .in3(N__4858),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__5237));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_10_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_10_9_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_LC_10_9_1  (
            .in0(N__4213),
            .in1(N__4192),
            .in2(N__5362),
            .in3(N__4171),
            .lcout(TACK_EN_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .ce(N__4156),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_LC_10_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_10_10_0 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_10_10_0 .LUT_INIT=16'b1111111101110000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_LC_10_10_0  (
            .in0(N__4102),
            .in1(N__4542),
            .in2(N__4134),
            .in3(N__4558),
            .lcout(ROMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .ce(),
            .sr(N__5244));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_10_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_10_5 .LUT_INIT=16'b1011111100100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_10_5  (
            .in0(N__4510),
            .in1(N__5068),
            .in2(N__4552),
            .in3(N__4116),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .ce(),
            .sr(N__5244));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_10_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_10_11_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_10_11_1  (
            .in0(N__5061),
            .in1(N__4530),
            .in2(N__5105),
            .in3(N__5131),
            .lcout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI6OQO2_0_LC_10_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI6OQO2_0_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI6OQO2_0_LC_10_11_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI6OQO2_0_LC_10_11_2  (
            .in0(N__4498),
            .in1(N__4650),
            .in2(N__4609),
            .in3(N__4773),
            .lcout(\U409_TRANSFER_ACK.N_28_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_10_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_10_11_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_10_11_4  (
            .in0(N__5130),
            .in1(N__5093),
            .in2(N__4508),
            .in3(N__5060),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_11_6 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_11_6  (
            .in0(N__5132),
            .in1(N__5094),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_EN_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_10_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_10_12_0 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_10_12_0  (
            .in0(N__4504),
            .in1(N__4543),
            .in2(N__4531),
            .in3(N__5032),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5238));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_10_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_10_12_1 .LUT_INIT=16'b0111100001111000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_10_12_1  (
            .in0(N__5063),
            .in1(N__4502),
            .in2(N__5106),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5238));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_10_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_10_12_3 .LUT_INIT=16'b0111101110000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_10_12_3  (
            .in0(N__5064),
            .in1(N__4503),
            .in2(N__5107),
            .in3(N__5134),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5238));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_10_12_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_10_12_4 .LUT_INIT=16'b0000111111010000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_10_12_4  (
            .in0(N__5133),
            .in1(N__5098),
            .in2(N__4509),
            .in3(N__5062),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5238));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_1_LC_11_6_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_1_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_1_LC_11_6_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_1_LC_11_6_2  (
            .in0(N__4926),
            .in1(N__4685),
            .in2(N__4912),
            .in3(N__4837),
            .lcout(\U409_TRANSFER_ACK.N_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_o2_0_LC_11_6_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_o2_0_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_o2_0_LC_11_6_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_o2_0_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__4908),
            .in2(_gnd_net_),
            .in3(N__4925),
            .lcout(\U409_TRANSFER_ACK.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_0_LC_11_7_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_0_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_0_LC_11_7_0 .LUT_INIT=16'b0001001100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_0_LC_11_7_0  (
            .in0(N__5391),
            .in1(N__4680),
            .in2(N__4900),
            .in3(N__4835),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.N_63_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_1_LC_11_7_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_1_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_1_LC_11_7_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_1_LC_11_7_1  (
            .in0(N__4856),
            .in1(N__4879),
            .in2(N__4873),
            .in3(N__4866),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.m9_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_7_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_7_2 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__5297),
            .in2(N__4870),
            .in3(N__4813),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_7_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_7_3 .LUT_INIT=16'b0011000000010000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_7_3  (
            .in0(N__4857),
            .in1(N__4843),
            .in2(N__5315),
            .in3(N__4867),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_LC_11_7_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_LC_11_7_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__4681),
            .in2(_gnd_net_),
            .in3(N__4834),
            .lcout(\U409_TRANSFER_ACK.N_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m12_0_a3_LC_11_7_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m12_0_a3_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m12_0_a3_LC_11_7_5 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m12_0_a3_LC_11_7_5  (
            .in0(N__4836),
            .in1(N__4898),
            .in2(N__4687),
            .in3(N__5393),
            .lcout(\U409_TRANSFER_ACK.N_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_0_LC_11_7_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_0_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_0_LC_11_7_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_0_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__4679),
            .in2(_gnd_net_),
            .in3(N__4833),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_2_LC_11_7_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_2_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_2_LC_11_7_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_2_LC_11_7_7  (
            .in0(N__4803),
            .in1(N__4897),
            .in2(N__4816),
            .in3(N__5392),
            .lcout(\U409_TRANSFER_ACK.N_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_8_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_8_3  (
            .in0(N__4899),
            .in1(N__5394),
            .in2(N__4807),
            .in3(N__4686),
            .lcout(\U409_TRANSFER_ACK.N_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_11_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_11_12_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_11_12_2  (
            .in0(N__5129),
            .in1(N__5092),
            .in2(_gnd_net_),
            .in3(N__5059),
            .lcout(\U409_TRANSFER_ACK.N_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_12_4_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_12_4_5 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_12_4_5  (
            .in0(N__5011),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4972),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS1n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNI692L_0_LC_12_4_6 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNI692L_0_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNI692L_0_LC_12_4_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_CIA.VMA_RNI692L_0_LC_12_4_6  (
            .in0(N__5280),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5158),
            .lcout(CIA_ENABLE),
            .ltout(CIA_ENABLE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_4_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_4_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_4_7 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4966),
            .in3(N__4963),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS0n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_6_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_6_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_6_1  (
            .in0(N__5157),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5281),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__5245));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_6_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4927),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__5245));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_12_7_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_12_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_12_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5395),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(N__5230));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_12_8_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_12_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5427),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__5239));
    defparam RESETn_ibuf_RNIM9SF_LC_12_10_3.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_10_3.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_10_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5301),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_12_11_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_12_11_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_12_11_0  (
            .in0(N__5565),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5634),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5603),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_2_LC_12_11_1 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_2_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_2_LC_12_11_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.VMA_RNO_2_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__5563),
            .in2(_gnd_net_),
            .in3(N__5733),
            .lcout(),
            .ltout(\U409_CIA.N_93_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_1_LC_12_11_2 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_1_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_1_LC_12_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.VMA_RNO_1_LC_12_11_2  (
            .in0(N__5451),
            .in1(N__5473),
            .in2(N__5176),
            .in3(N__5633),
            .lcout(),
            .ltout(\U409_CIA.VMA_RNOZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_12_11_3 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_12_11_3 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \U409_CIA.VMA_LC_12_11_3  (
            .in0(N__5150),
            .in1(N__5564),
            .in2(N__5173),
            .in3(N__5170),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5603),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_12_12_0 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_12_12_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_1_LC_12_12_0  (
            .in0(N__5751),
            .in1(N__5732),
            .in2(N__5656),
            .in3(N__5679),
            .lcout(\U409_CIA.un1_CIA_CLK_COUNT_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_12_12_1 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_12_12_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_12_12_1  (
            .in0(N__5651),
            .in1(N__5678),
            .in2(_gnd_net_),
            .in3(N__5750),
            .lcout(\U409_CIA.N_91 ),
            .ltout(\U409_CIA.N_91_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_12_12_2 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_12_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_12_12_2  (
            .in0(N__5566),
            .in1(N__5632),
            .in2(N__5137),
            .in3(N__5479),
            .lcout(\U409_CIA.CIA_CLK_COUNT11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIBFRM_2_LC_12_12_3 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIBFRM_2_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIBFRM_2_LC_12_12_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIBFRM_2_LC_12_12_3  (
            .in0(N__5769),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5697),
            .lcout(\U409_CIA.CLK_CIA6_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_12_12_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_12_12_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_12_12_4  (
            .in0(N__5696),
            .in1(N__5730),
            .in2(_gnd_net_),
            .in3(N__5768),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_12_12_6 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_12_12_6 .LUT_INIT=16'b0000010110001101;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_0_LC_12_12_6  (
            .in0(N__5542),
            .in1(N__5472),
            .in2(N__5426),
            .in3(N__5731),
            .lcout(),
            .ltout(\U409_CIA.CLK_CIA_r_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_LC_12_12_7 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLK_CIA_LC_12_12_7 .LUT_INIT=16'b0000111011001100;
    LogicCell40 \U409_CIA.CLK_CIA_LC_12_12_7  (
            .in0(N__5461),
            .in1(N__5419),
            .in2(N__5455),
            .in3(N__5452),
            .lcout(CLK_CIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5605),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_13_1_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_13_1_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_13_1_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_13_1_0  (
            .in0(_gnd_net_),
            .in1(N__6316),
            .in2(_gnd_net_),
            .in3(N__5814),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6678),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_13_1_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_13_1_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_13_1_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_13_1_2  (
            .in0(N__6229),
            .in1(N__6390),
            .in2(N__5491),
            .in3(N__6351),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6678),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_13_1_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_13_1_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_13_1_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_13_1_3  (
            .in0(N__6475),
            .in1(N__6517),
            .in2(N__6622),
            .in3(N__6562),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_13_1_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_13_1_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_13_1_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_13_1_4  (
            .in0(N__6009),
            .in1(N__5972),
            .in2(N__5401),
            .in3(N__6604),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6678),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_13_1_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_13_1_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_13_1_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_13_1_5  (
            .in0(N__6097),
            .in1(N__6133),
            .in2(_gnd_net_),
            .in3(N__6169),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_13_1_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_13_1_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_13_1_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_13_1_6  (
            .in0(N__5848),
            .in1(N__6496),
            .in2(N__5398),
            .in3(N__6538),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_13_1_7 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_13_1_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_13_1_7 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \U409_TICK.TICK50_LC_13_1_7  (
            .in0(N__5520),
            .in1(N__6010),
            .in2(N__5536),
            .in3(N__5925),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6678),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_2_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_2_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_2_0  (
            .in0(_gnd_net_),
            .in1(N__5810),
            .in2(N__6312),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_2_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_13_2_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_13_2_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_13_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_13_2_1  (
            .in0(_gnd_net_),
            .in1(N__5826),
            .in2(_gnd_net_),
            .in3(N__5509),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__6679),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_13_2_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_13_2_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_13_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_13_2_2  (
            .in0(_gnd_net_),
            .in1(N__6042),
            .in2(_gnd_net_),
            .in3(N__5506),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__6679),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_13_2_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_13_2_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_13_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_13_2_3  (
            .in0(_gnd_net_),
            .in1(N__6021),
            .in2(_gnd_net_),
            .in3(N__5503),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_13_2_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_13_2_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_13_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_13_2_4  (
            .in0(_gnd_net_),
            .in1(N__6075),
            .in2(_gnd_net_),
            .in3(N__5500),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__6679),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_13_2_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_13_2_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_13_2_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_13_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6420),
            .in3(N__5497),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_13_2_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_13_2_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_13_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_13_2_6  (
            .in0(_gnd_net_),
            .in1(N__6252),
            .in2(_gnd_net_),
            .in3(N__5494),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__6679),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_13_2_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_13_2_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_13_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_13_2_7  (
            .in0(_gnd_net_),
            .in1(N__6435),
            .in2(_gnd_net_),
            .in3(N__5482),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_13_3_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_13_3_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_13_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_13_3_0  (
            .in0(_gnd_net_),
            .in1(N__6450),
            .in2(_gnd_net_),
            .in3(N__5590),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_13_3_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_13_3_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_13_3_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_13_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_13_3_1  (
            .in0(_gnd_net_),
            .in1(N__6270),
            .in2(_gnd_net_),
            .in3(N__5587),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__6681),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_13_3_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_13_3_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_13_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_13_3_2  (
            .in0(_gnd_net_),
            .in1(N__6063),
            .in2(_gnd_net_),
            .in3(N__5584),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__6681),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_13_3_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_13_3_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_13_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_13_3_3  (
            .in0(_gnd_net_),
            .in1(N__5838),
            .in2(_gnd_net_),
            .in3(N__5581),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__6681),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_13_3_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_13_3_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_13_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_13_3_4  (
            .in0(_gnd_net_),
            .in1(N__6282),
            .in2(_gnd_net_),
            .in3(N__5578),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__6681),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_13_3_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_13_3_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_13_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_13_3_5  (
            .in0(_gnd_net_),
            .in1(N__6402),
            .in2(_gnd_net_),
            .in3(N__5575),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_13_3_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_13_3_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_13_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_13_3_6  (
            .in0(_gnd_net_),
            .in1(N__6240),
            .in2(_gnd_net_),
            .in3(N__5572),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_13_3_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_13_3_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_13_3_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_13_3_7  (
            .in0(_gnd_net_),
            .in1(N__5794),
            .in2(_gnd_net_),
            .in3(N__5569),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6681),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_13_12_0 .C_ON=1'b1;
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_13_12_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_2_LC_13_12_0  (
            .in0(N__5627),
            .in1(N__5562),
            .in2(N__5635),
            .in3(_gnd_net_),
            .lcout(\U409_CIA.CLK_CIA6_1 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_13_12_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_13_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__5770),
            .in2(_gnd_net_),
            .in3(N__5755),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__5604),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_13_12_2 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_13_12_2 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_13_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_13_12_2  (
            .in0(N__5706),
            .in1(N__5752),
            .in2(_gnd_net_),
            .in3(N__5737),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(N__5604),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_13_12_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_13_12_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_13_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__5734),
            .in2(_gnd_net_),
            .in3(N__5710),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__5604),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_13_12_4 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_13_12_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_13_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_13_12_4  (
            .in0(N__5707),
            .in1(N__5698),
            .in2(_gnd_net_),
            .in3(N__5683),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .clk(N__5604),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_13_12_5 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_13_12_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_13_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_6_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__5680),
            .in2(_gnd_net_),
            .in3(N__5662),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ),
            .clk(N__5604),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_13_12_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_13_12_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_13_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_7_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__5655),
            .in2(_gnd_net_),
            .in3(N__5659),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5604),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_13_12_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_13_12_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_13_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5631),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5604),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_14_1_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_14_1_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_14_1_0 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_14_1_0  (
            .in0(N__6003),
            .in1(N__5969),
            .in2(N__6175),
            .in3(N__5926),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6680),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_14_1_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_14_1_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_14_1_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_14_1_1  (
            .in0(N__5968),
            .in1(N__6006),
            .in2(N__5938),
            .in3(N__6085),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6680),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_14_1_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_14_1_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_14_1_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_14_1_2  (
            .in0(N__6004),
            .in1(N__5970),
            .in2(N__6733),
            .in3(N__5927),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6680),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_14_1_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_14_1_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_14_1_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_14_1_3  (
            .in0(N__5967),
            .in1(N__6005),
            .in2(N__5937),
            .in3(N__6709),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6680),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_1_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_1_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_1_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_1_4  (
            .in0(N__6577),
            .in1(N__6148),
            .in2(N__6193),
            .in3(N__6696),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_14_1_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_14_1_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_14_1_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_14_1_5  (
            .in0(N__6592),
            .in1(N__6745),
            .in2(N__6115),
            .in3(N__6721),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_14_1_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_14_1_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_14_1_6 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_14_1_6  (
            .in0(N__6547),
            .in1(N__5971),
            .in2(N__5842),
            .in3(N__5934),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6680),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_14_1_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_14_1_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_14_1_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_14_1_7  (
            .in0(_gnd_net_),
            .in1(N__6170),
            .in2(_gnd_net_),
            .in3(N__6192),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6680),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_14_2_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_14_2_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_14_2_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_14_2_0  (
            .in0(N__5839),
            .in1(N__5827),
            .in2(N__5815),
            .in3(N__5793),
            .lcout(\U409_TICK.TICK603_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_14_2_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_14_2_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_14_2_1 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_14_2_1  (
            .in0(N__6388),
            .in1(N__6350),
            .in2(N__5782),
            .in3(N__6228),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6682),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_14_2_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_14_2_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_14_2_2 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_14_2_2  (
            .in0(N__6007),
            .in1(N__6505),
            .in2(N__5977),
            .in3(N__5935),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6682),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_2_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_2_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_2_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_2_3  (
            .in0(N__6076),
            .in1(N__6022),
            .in2(_gnd_net_),
            .in3(N__6307),
            .lcout(),
            .ltout(\U409_TICK.TICK603_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_14_2_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_14_2_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_14_2_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_14_2_4  (
            .in0(N__6064),
            .in1(N__6052),
            .in2(N__6046),
            .in3(N__6043),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_14_2_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_14_2_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_14_2_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_14_2_5  (
            .in0(N__6387),
            .in1(N__6226),
            .in2(N__6031),
            .in3(N__6028),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6682),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_14_2_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_14_2_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_14_2_6 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_14_2_6  (
            .in0(N__6008),
            .in1(N__5976),
            .in2(N__6463),
            .in3(N__5936),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6682),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_14_2_7 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_14_2_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_14_2_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK60_LC_14_2_7  (
            .in0(N__6389),
            .in1(N__5886),
            .in2(N__6355),
            .in3(N__6227),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6682),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_14_3_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_14_3_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_14_3_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_14_3_0  (
            .in0(N__6347),
            .in1(N__6224),
            .in2(N__5875),
            .in3(N__6385),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6684),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_14_3_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_14_3_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_14_3_1 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_14_3_1  (
            .in0(N__6222),
            .in1(N__5863),
            .in2(N__6391),
            .in3(N__6349),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6684),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_14_3_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_14_3_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_14_3_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_14_3_2  (
            .in0(N__6348),
            .in1(N__6225),
            .in2(N__5857),
            .in3(N__6386),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6684),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_3_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_3_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_14_3_5  (
            .in0(N__6451),
            .in1(N__6439),
            .in2(N__6424),
            .in3(N__6403),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_14_3_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_14_3_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_14_3_6 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_14_3_6  (
            .in0(N__6346),
            .in1(N__6223),
            .in2(N__6319),
            .in3(N__6311),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6684),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_14_3_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_14_3_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_14_3_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_14_3_7  (
            .in0(N__6283),
            .in1(N__6271),
            .in2(N__6259),
            .in3(N__6241),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_1_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_1_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_1_0  (
            .in0(_gnd_net_),
            .in1(N__6188),
            .in2(N__6174),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_1_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_15_1_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_15_1_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_15_1_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_15_1_1  (
            .in0(_gnd_net_),
            .in1(N__6147),
            .in2(_gnd_net_),
            .in3(N__6136),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__6683),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_15_1_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_15_1_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_15_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_15_1_2  (
            .in0(_gnd_net_),
            .in1(N__6129),
            .in2(_gnd_net_),
            .in3(N__6118),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__6683),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_15_1_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_15_1_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_15_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_15_1_3  (
            .in0(_gnd_net_),
            .in1(N__6111),
            .in2(_gnd_net_),
            .in3(N__6100),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__6683),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_15_1_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_15_1_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_15_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_15_1_4  (
            .in0(_gnd_net_),
            .in1(N__6096),
            .in2(_gnd_net_),
            .in3(N__6079),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_15_1_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_15_1_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_15_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_15_1_5  (
            .in0(_gnd_net_),
            .in1(N__6621),
            .in2(_gnd_net_),
            .in3(N__6595),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_15_1_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_15_1_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_15_1_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_15_1_6  (
            .in0(_gnd_net_),
            .in1(N__6591),
            .in2(_gnd_net_),
            .in3(N__6580),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__6683),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_15_1_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_15_1_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_15_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_15_1_7  (
            .in0(_gnd_net_),
            .in1(N__6576),
            .in2(_gnd_net_),
            .in3(N__6565),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__6683),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_15_2_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_15_2_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_15_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_15_2_0  (
            .in0(_gnd_net_),
            .in1(N__6558),
            .in2(_gnd_net_),
            .in3(N__6541),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_15_2_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_15_2_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_15_2_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_15_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_15_2_1  (
            .in0(_gnd_net_),
            .in1(N__6531),
            .in2(_gnd_net_),
            .in3(N__6520),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__6685),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_15_2_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_15_2_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_15_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_15_2_2  (
            .in0(_gnd_net_),
            .in1(N__6516),
            .in2(_gnd_net_),
            .in3(N__6499),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_15_2_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_15_2_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_15_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_15_2_3  (
            .in0(_gnd_net_),
            .in1(N__6489),
            .in2(_gnd_net_),
            .in3(N__6478),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__6685),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_15_2_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_15_2_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_15_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_15_2_4  (
            .in0(_gnd_net_),
            .in1(N__6474),
            .in2(_gnd_net_),
            .in3(N__6454),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_15_2_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_15_2_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_15_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_15_2_5  (
            .in0(_gnd_net_),
            .in1(N__6744),
            .in2(_gnd_net_),
            .in3(N__6724),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_15_2_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_15_2_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_15_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_15_2_6  (
            .in0(_gnd_net_),
            .in1(N__6720),
            .in2(_gnd_net_),
            .in3(N__6703),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_15_2_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_15_2_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_15_2_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_15_2_7  (
            .in0(_gnd_net_),
            .in1(N__6697),
            .in2(_gnd_net_),
            .in3(N__6700),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6685),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_iobuf_RNO_LC_17_15_4.C_ON=1'b0;
    defparam TACKn_iobuf_RNO_LC_17_15_4.SEQ_MODE=4'b0000;
    defparam TACKn_iobuf_RNO_LC_17_15_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_iobuf_RNO_LC_17_15_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6655),
            .lcout(N_525_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 25 2024 14:30:47

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RAMENn : out std_logic;
    RASn : out std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__10026\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_OUT_i_i\ : std_logic;
signal \N_839_i\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4_cascade_\ : std_logic;
signal \A_c_6\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.N_319\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.N_318\ : std_logic;
signal \CLK40_OUT_i_i\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_0_a2_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_181\ : std_logic;
signal \CLK40_OUT_i\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_307_i_0_en_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \U712_CYCLE_TERM.N_307_i_0_en_0\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_CHIP_RAM.N_287_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_1_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \TSn_c\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_GOZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \U712_REG_SM.LDS_OUT_2_0_a2Z0Z_0\ : std_logic;
signal \U712_REG_SM.N_342\ : std_logic;
signal \U712_REG_SM.LDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_LDSn_i\ : std_logic;
signal \U712_REG_SM.UDS_OUTZ0\ : std_logic;
signal \U712_REG_SM.DS_ENZ0\ : std_logic;
signal \U712_REG_SM_un1_UDSn_i\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_287\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_273_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_0\ : std_logic;
signal \U712_CHIP_RAM.N_347_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_378_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_tz\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_0_a2_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER50_cascade_\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_296_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_e_1_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_0_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \N_188\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_1\ : std_logic;
signal \U712_REG_SM.N_288_cascade_\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_5\ : std_logic;
signal \U712_REG_SM.N_301_cascade_\ : std_logic;
signal \U712_REG_SM.N_288\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.N_301\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_341\ : std_logic;
signal \U712_REG_SM.N_294_cascade_\ : std_logic;
signal \U712_REG_SM.N_373\ : std_logic;
signal \U712_REG_SM.N_292_cascade_\ : std_logic;
signal \U712_REG_SM.N_507\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U712_REG_SM.N_104\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_372\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_186_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_0_a2_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_393\ : std_logic;
signal \U712_CHIP_RAM.N_310\ : std_logic;
signal \U712_CHIP_RAM.N_310_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_46\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_3_0_a2_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_179_cascade_\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_438_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_289\ : std_logic;
signal \U712_CHIP_RAM.N_425_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_424\ : std_logic;
signal \U712_CHIP_RAM.N_302\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_START_2_0_a2_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_438\ : std_logic;
signal \U712_CHIP_RAM.N_284\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_272\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.DBENn_7_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_347\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_3_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_2_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER50\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_273\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_305\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST_cascade_\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0_cascade_\ : std_logic;
signal \N_192_i\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0\ : std_logic;
signal \N_194_i\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_cascade_\ : std_logic;
signal \N_196_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_404\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_411_cascade_\ : std_logic;
signal \N_198_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_405\ : std_logic;
signal \U712_REG_SM.N_292\ : std_logic;
signal \U712_REG_SM.N_298\ : std_logic;
signal \U712_REG_SM.N_294\ : std_logic;
signal \U712_REG_SM.N_309\ : std_logic;
signal \U712_REG_SM.N_282\ : std_logic;
signal \U712_REG_SM.N_282_cascade_\ : std_logic;
signal \U712_REG_SM.N_306\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \U712_BYTE_ENABLE.N_407\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_409\ : std_logic;
signal \C1_c\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.N_317\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5_cascade_\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6_cascade_\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_315_cascade_\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_316\ : std_logic;
signal \U712_CHIP_RAM.N_425\ : std_logic;
signal \U712_CHIP_RAM.N_276\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_314\ : std_logic;
signal \U712_CHIP_RAM.N_293\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH9lt7_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH9lto7_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_321\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.N_320\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH9lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.N_322_cascade_\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_8_cascade_\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    CLK_EN <= \CLK_EN_wire\;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    LDSn <= \LDSn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_OUT_i\,
            REFERENCECLK => \N__3617\,
            RESETB => \N__7409\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_OUT\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10026\,
            DIN => \N__10025\,
            DOUT => \N__10024\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10026\,
            PADOUT => \N__10025\,
            PADIN => \N__10024\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6038\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10017\,
            DIN => \N__10016\,
            DOUT => \N__10015\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10017\,
            PADOUT => \N__10016\,
            PADIN => \N__10015\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10008\,
            DIN => \N__10007\,
            DOUT => \N__10006\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10008\,
            PADOUT => \N__10007\,
            PADIN => \N__10006\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8396\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9999\,
            DIN => \N__9998\,
            DOUT => \N__9997\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9999\,
            PADOUT => \N__9998\,
            PADIN => \N__9997\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4589\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9990\,
            DIN => \N__9989\,
            DOUT => \N__9988\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9990\,
            PADOUT => \N__9989\,
            PADIN => \N__9988\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9981\,
            DIN => \N__9980\,
            DOUT => \N__9979\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9981\,
            PADOUT => \N__9980\,
            PADIN => \N__9979\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9972\,
            DIN => \N__9971\,
            DOUT => \N__9970\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9972\,
            PADOUT => \N__9971\,
            PADIN => \N__9970\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9963\,
            DIN => \N__9962\,
            DOUT => \N__9961\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9963\,
            PADOUT => \N__9962\,
            PADIN => \N__9961\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9954\,
            DIN => \N__9953\,
            DOUT => \N__9952\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9954\,
            PADOUT => \N__9953\,
            PADIN => \N__9952\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9945\,
            DIN => \N__9944\,
            DOUT => \N__9943\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9945\,
            PADOUT => \N__9944\,
            PADIN => \N__9943\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9936\,
            DIN => \N__9935\,
            DOUT => \N__9934\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9936\,
            PADOUT => \N__9935\,
            PADIN => \N__9934\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8225\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9927\,
            DIN => \N__9926\,
            DOUT => \N__9925\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9927\,
            PADOUT => \N__9926\,
            PADIN => \N__9925\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5996\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9918\,
            DIN => \N__9917\,
            DOUT => \N__9916\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9918\,
            PADOUT => \N__9917\,
            PADIN => \N__9916\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9909\,
            DIN => \N__9908\,
            DOUT => \N__9907\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9909\,
            PADOUT => \N__9908\,
            PADIN => \N__9907\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9900\,
            DIN => \N__9899\,
            DOUT => \N__9898\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9900\,
            PADOUT => \N__9899\,
            PADIN => \N__9898\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3917\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9891\,
            DIN => \N__9890\,
            DOUT => \N__9889\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9891\,
            PADOUT => \N__9890\,
            PADIN => \N__9889\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9882\,
            DIN => \N__9881\,
            DOUT => \N__9880\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9882\,
            PADOUT => \N__9881\,
            PADIN => \N__9880\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9873\,
            DIN => \N__9872\,
            DOUT => \N__9871\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9873\,
            PADOUT => \N__9872\,
            PADIN => \N__9871\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6719\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9864\,
            DIN => \N__9863\,
            DOUT => \N__9862\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9864\,
            PADOUT => \N__9863\,
            PADIN => \N__9862\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9855\,
            DIN => \N__9854\,
            DOUT => \N__9853\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9855\,
            PADOUT => \N__9854\,
            PADIN => \N__9853\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7025\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9846\,
            DIN => \N__9845\,
            DOUT => \N__9844\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9846\,
            PADOUT => \N__9845\,
            PADIN => \N__9844\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9837\,
            DIN => \N__9836\,
            DOUT => \N__9835\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9837\,
            PADOUT => \N__9836\,
            PADIN => \N__9835\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9828\,
            DIN => \N__9827\,
            DOUT => \N__9826\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9828\,
            PADOUT => \N__9827\,
            PADIN => \N__9826\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9819\,
            DIN => \N__9818\,
            DOUT => \N__9817\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9819\,
            PADOUT => \N__9818\,
            PADIN => \N__9817\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9810\,
            DIN => \N__9809\,
            DOUT => \N__9808\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9810\,
            PADOUT => \N__9809\,
            PADIN => \N__9808\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9801\,
            DIN => \N__9800\,
            DOUT => \N__9799\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9801\,
            PADOUT => \N__9800\,
            PADIN => \N__9799\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5141\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9792\,
            DIN => \N__9791\,
            DOUT => \N__9790\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9792\,
            PADOUT => \N__9791\,
            PADIN => \N__9790\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9783\,
            DIN => \N__9782\,
            DOUT => \N__9781\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9783\,
            PADOUT => \N__9782\,
            PADIN => \N__9781\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9774\,
            DIN => \N__9773\,
            DOUT => \N__9772\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9774\,
            PADOUT => \N__9773\,
            PADIN => \N__9772\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9765\,
            DIN => \N__9764\,
            DOUT => \N__9763\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9765\,
            PADOUT => \N__9764\,
            PADIN => \N__9763\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9756\,
            DIN => \N__9755\,
            DOUT => \N__9754\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9756\,
            PADOUT => \N__9755\,
            PADIN => \N__9754\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9747\,
            DIN => \N__9746\,
            DOUT => \N__9745\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9747\,
            PADOUT => \N__9746\,
            PADIN => \N__9745\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7313\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9738\,
            DIN => \N__9737\,
            DOUT => \N__9736\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9738\,
            PADOUT => \N__9737\,
            PADIN => \N__9736\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9729\,
            DIN => \N__9728\,
            DOUT => \N__9727\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9729\,
            PADOUT => \N__9728\,
            PADIN => \N__9727\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9720\,
            DIN => \N__9719\,
            DOUT => \N__9718\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9720\,
            PADOUT => \N__9719\,
            PADIN => \N__9718\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9711\,
            DIN => \N__9710\,
            DOUT => \N__9709\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9711\,
            PADOUT => \N__9710\,
            PADIN => \N__9709\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9702\,
            DIN => \N__9701\,
            DOUT => \N__9700\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9702\,
            PADOUT => \N__9701\,
            PADIN => \N__9700\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3674\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9693\,
            DIN => \N__9692\,
            DOUT => \N__9691\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9693\,
            PADOUT => \N__9692\,
            PADIN => \N__9691\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4331\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9684\,
            DIN => \N__9683\,
            DOUT => \N__9682\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9684\,
            PADOUT => \N__9683\,
            PADIN => \N__9682\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9675\,
            DIN => \N__9674\,
            DOUT => \N__9673\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9675\,
            PADOUT => \N__9674\,
            PADIN => \N__9673\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8660\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9666\,
            DIN => \N__9665\,
            DOUT => \N__9664\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9666\,
            PADOUT => \N__9665\,
            PADIN => \N__9664\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9657\,
            DIN => \N__9656\,
            DOUT => \N__9655\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9657\,
            PADOUT => \N__9656\,
            PADIN => \N__9655\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9648\,
            DIN => \N__9647\,
            DOUT => \N__9646\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9648\,
            PADOUT => \N__9647\,
            PADIN => \N__9646\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3653\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9639\,
            DIN => \N__9638\,
            DOUT => \N__9637\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9639\,
            PADOUT => \N__9638\,
            PADIN => \N__9637\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9630\,
            DIN => \N__9629\,
            DOUT => \N__9628\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9630\,
            PADOUT => \N__9629\,
            PADIN => \N__9628\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4898\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9621\,
            DIN => \N__9620\,
            DOUT => \N__9619\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9621\,
            PADOUT => \N__9620\,
            PADIN => \N__9619\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3758\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9612\,
            DIN => \N__9611\,
            DOUT => \N__9610\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9612\,
            PADOUT => \N__9611\,
            PADIN => \N__9610\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9603\,
            DIN => \N__9602\,
            DOUT => \N__9601\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9603\,
            PADOUT => \N__9602\,
            PADIN => \N__9601\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9594\,
            DIN => \N__9593\,
            DOUT => \N__9592\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9594\,
            PADOUT => \N__9593\,
            PADIN => \N__9592\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9585\,
            DIN => \N__9584\,
            DOUT => \N__9583\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9585\,
            PADOUT => \N__9584\,
            PADIN => \N__9583\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6476\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9576\,
            DIN => \N__9575\,
            DOUT => \N__9574\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9576\,
            PADOUT => \N__9575\,
            PADIN => \N__9574\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9567\,
            DIN => \N__9566\,
            DOUT => \N__9565\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9567\,
            PADOUT => \N__9566\,
            PADIN => \N__9565\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3737\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9558\,
            DIN => \N__9557\,
            DOUT => \N__9556\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9558\,
            PADOUT => \N__9557\,
            PADIN => \N__9556\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4721\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9549\,
            DIN => \N__9548\,
            DOUT => \N__9547\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9549\,
            PADOUT => \N__9548\,
            PADIN => \N__9547\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5888\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9540\,
            DIN => \N__9539\,
            DOUT => \N__9538\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9540\,
            PADOUT => \N__9539\,
            PADIN => \N__9538\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7988\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9531\,
            DIN => \N__9530\,
            DOUT => \N__9529\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9531\,
            PADOUT => \N__9530\,
            PADIN => \N__9529\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4894\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9522\,
            DIN => \N__9521\,
            DOUT => \N__9520\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9522\,
            PADOUT => \N__9521\,
            PADIN => \N__9520\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9513\,
            DIN => \N__9512\,
            DOUT => \N__9511\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9513\,
            PADOUT => \N__9512\,
            PADIN => \N__9511\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9504\,
            DIN => \N__9503\,
            DOUT => \N__9502\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9504\,
            PADOUT => \N__9503\,
            PADIN => \N__9502\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5933\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9495\,
            DIN => \N__9494\,
            DOUT => \N__9493\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9495\,
            PADOUT => \N__9494\,
            PADIN => \N__9493\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8543\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9486\,
            DIN => \N__9485\,
            DOUT => \N__9484\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9486\,
            PADOUT => \N__9485\,
            PADIN => \N__9484\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4628\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9477\,
            DIN => \N__9476\,
            DOUT => \N__9475\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9477\,
            PADOUT => \N__9476\,
            PADIN => \N__9475\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6083\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9468\,
            DIN => \N__9467\,
            DOUT => \N__9466\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9468\,
            PADOUT => \N__9467\,
            PADIN => \N__9466\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9459\,
            DIN => \N__9458\,
            DOUT => \N__9457\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9459\,
            PADOUT => \N__9458\,
            PADIN => \N__9457\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9450\,
            DIN => \N__9449\,
            DOUT => \N__9448\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9450\,
            PADOUT => \N__9449\,
            PADIN => \N__9448\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9441\,
            DIN => \N__9440\,
            DOUT => \N__9439\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9441\,
            PADOUT => \N__9440\,
            PADIN => \N__9439\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9432\,
            DIN => \N__9431\,
            DOUT => \N__9430\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9432\,
            PADOUT => \N__9431\,
            PADIN => \N__9430\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6488\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9423\,
            DIN => \N__9422\,
            DOUT => \N__9421\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9423\,
            PADOUT => \N__9422\,
            PADIN => \N__9421\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9414\,
            DIN => \N__9413\,
            DOUT => \N__9412\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9414\,
            PADOUT => \N__9413\,
            PADIN => \N__9412\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6110\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9405\,
            DIN => \N__9404\,
            DOUT => \N__9403\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9405\,
            PADOUT => \N__9404\,
            PADIN => \N__9403\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3635\,
            DIN0 => OPEN,
            DOUT0 => \N__3860\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9396\,
            DIN => \N__9395\,
            DOUT => \N__9394\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9396\,
            PADOUT => \N__9395\,
            PADIN => \N__9394\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6497\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9387\,
            DIN => \N__9386\,
            DOUT => \N__9385\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9387\,
            PADOUT => \N__9386\,
            PADIN => \N__9385\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9378\,
            DIN => \N__9377\,
            DOUT => \N__9376\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9378\,
            PADOUT => \N__9377\,
            PADIN => \N__9376\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9369\,
            DIN => \N__9368\,
            DOUT => \N__9367\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9369\,
            PADOUT => \N__9368\,
            PADIN => \N__9367\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7256\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9360\,
            DIN => \N__9359\,
            DOUT => \N__9358\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9360\,
            PADOUT => \N__9359\,
            PADIN => \N__9358\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9351\,
            DIN => \N__9350\,
            DOUT => \N__9349\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9351\,
            PADOUT => \N__9350\,
            PADIN => \N__9349\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9342\,
            DIN => \N__9341\,
            DOUT => \N__9340\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9342\,
            PADOUT => \N__9341\,
            PADIN => \N__9340\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9333\,
            DIN => \N__9332\,
            DOUT => \N__9331\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9333\,
            PADOUT => \N__9332\,
            PADIN => \N__9331\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9324\,
            DIN => \N__9323\,
            DOUT => \N__9322\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9324\,
            PADOUT => \N__9323\,
            PADIN => \N__9322\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7286\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9315\,
            DIN => \N__9314\,
            DOUT => \N__9313\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9315\,
            PADOUT => \N__9314\,
            PADIN => \N__9313\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4268\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2203\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9292\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9289\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__9292\,
            I => \N__9286\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__9289\,
            I => \N__9283\
        );

    \I__2199\ : Span4Mux_v
    port map (
            O => \N__9286\,
            I => \N__9280\
        );

    \I__2198\ : Span4Mux_h
    port map (
            O => \N__9283\,
            I => \N__9277\
        );

    \I__2197\ : Span4Mux_v
    port map (
            O => \N__9280\,
            I => \N__9274\
        );

    \I__2196\ : Span4Mux_v
    port map (
            O => \N__9277\,
            I => \N__9271\
        );

    \I__2195\ : Sp12to4
    port map (
            O => \N__9274\,
            I => \N__9266\
        );

    \I__2194\ : Sp12to4
    port map (
            O => \N__9271\,
            I => \N__9266\
        );

    \I__2193\ : Span12Mux_h
    port map (
            O => \N__9266\,
            I => \N__9263\
        );

    \I__2192\ : Span12Mux_v
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__2191\ : Odrv12
    port map (
            O => \N__9260\,
            I => \DRA_c_0\
        );

    \I__2190\ : InMux
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__9254\,
            I => \N__9251\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__9251\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9245\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9245\,
            I => \N__9219\
        );

    \I__2185\ : ClkMux
    port map (
            O => \N__9244\,
            I => \N__9119\
        );

    \I__2184\ : ClkMux
    port map (
            O => \N__9243\,
            I => \N__9119\
        );

    \I__2183\ : ClkMux
    port map (
            O => \N__9242\,
            I => \N__9119\
        );

    \I__2182\ : ClkMux
    port map (
            O => \N__9241\,
            I => \N__9119\
        );

    \I__2181\ : ClkMux
    port map (
            O => \N__9240\,
            I => \N__9119\
        );

    \I__2180\ : ClkMux
    port map (
            O => \N__9239\,
            I => \N__9119\
        );

    \I__2179\ : ClkMux
    port map (
            O => \N__9238\,
            I => \N__9119\
        );

    \I__2178\ : ClkMux
    port map (
            O => \N__9237\,
            I => \N__9119\
        );

    \I__2177\ : ClkMux
    port map (
            O => \N__9236\,
            I => \N__9119\
        );

    \I__2176\ : ClkMux
    port map (
            O => \N__9235\,
            I => \N__9119\
        );

    \I__2175\ : ClkMux
    port map (
            O => \N__9234\,
            I => \N__9119\
        );

    \I__2174\ : ClkMux
    port map (
            O => \N__9233\,
            I => \N__9119\
        );

    \I__2173\ : ClkMux
    port map (
            O => \N__9232\,
            I => \N__9119\
        );

    \I__2172\ : ClkMux
    port map (
            O => \N__9231\,
            I => \N__9119\
        );

    \I__2171\ : ClkMux
    port map (
            O => \N__9230\,
            I => \N__9119\
        );

    \I__2170\ : ClkMux
    port map (
            O => \N__9229\,
            I => \N__9119\
        );

    \I__2169\ : ClkMux
    port map (
            O => \N__9228\,
            I => \N__9119\
        );

    \I__2168\ : ClkMux
    port map (
            O => \N__9227\,
            I => \N__9119\
        );

    \I__2167\ : ClkMux
    port map (
            O => \N__9226\,
            I => \N__9119\
        );

    \I__2166\ : ClkMux
    port map (
            O => \N__9225\,
            I => \N__9119\
        );

    \I__2165\ : ClkMux
    port map (
            O => \N__9224\,
            I => \N__9119\
        );

    \I__2164\ : ClkMux
    port map (
            O => \N__9223\,
            I => \N__9119\
        );

    \I__2163\ : ClkMux
    port map (
            O => \N__9222\,
            I => \N__9119\
        );

    \I__2162\ : Glb2LocalMux
    port map (
            O => \N__9219\,
            I => \N__9119\
        );

    \I__2161\ : ClkMux
    port map (
            O => \N__9218\,
            I => \N__9119\
        );

    \I__2160\ : ClkMux
    port map (
            O => \N__9217\,
            I => \N__9119\
        );

    \I__2159\ : ClkMux
    port map (
            O => \N__9216\,
            I => \N__9119\
        );

    \I__2158\ : ClkMux
    port map (
            O => \N__9215\,
            I => \N__9119\
        );

    \I__2157\ : ClkMux
    port map (
            O => \N__9214\,
            I => \N__9119\
        );

    \I__2156\ : ClkMux
    port map (
            O => \N__9213\,
            I => \N__9119\
        );

    \I__2155\ : ClkMux
    port map (
            O => \N__9212\,
            I => \N__9119\
        );

    \I__2154\ : ClkMux
    port map (
            O => \N__9211\,
            I => \N__9119\
        );

    \I__2153\ : ClkMux
    port map (
            O => \N__9210\,
            I => \N__9119\
        );

    \I__2152\ : ClkMux
    port map (
            O => \N__9209\,
            I => \N__9119\
        );

    \I__2151\ : ClkMux
    port map (
            O => \N__9208\,
            I => \N__9119\
        );

    \I__2150\ : ClkMux
    port map (
            O => \N__9207\,
            I => \N__9119\
        );

    \I__2149\ : ClkMux
    port map (
            O => \N__9206\,
            I => \N__9119\
        );

    \I__2148\ : ClkMux
    port map (
            O => \N__9205\,
            I => \N__9119\
        );

    \I__2147\ : ClkMux
    port map (
            O => \N__9204\,
            I => \N__9119\
        );

    \I__2146\ : ClkMux
    port map (
            O => \N__9203\,
            I => \N__9119\
        );

    \I__2145\ : ClkMux
    port map (
            O => \N__9202\,
            I => \N__9119\
        );

    \I__2144\ : GlobalMux
    port map (
            O => \N__9119\,
            I => \CLK80_OUT\
        );

    \I__2143\ : CEMux
    port map (
            O => \N__9116\,
            I => \N__9113\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9113\,
            I => \N__9109\
        );

    \I__2141\ : CEMux
    port map (
            O => \N__9112\,
            I => \N__9105\
        );

    \I__2140\ : Span4Mux_h
    port map (
            O => \N__9109\,
            I => \N__9102\
        );

    \I__2139\ : CEMux
    port map (
            O => \N__9108\,
            I => \N__9099\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9105\,
            I => \N__9096\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__9102\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9099\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__2135\ : Odrv12
    port map (
            O => \N__9096\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__2134\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9077\
        );

    \I__2133\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9072\
        );

    \I__2132\ : InMux
    port map (
            O => \N__9087\,
            I => \N__9072\
        );

    \I__2131\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9069\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9085\,
            I => \N__9066\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9063\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9083\,
            I => \N__9060\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9082\,
            I => \N__9057\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9081\,
            I => \N__9054\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9051\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9077\,
            I => \N__9047\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__9072\,
            I => \N__9043\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9069\,
            I => \N__9040\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__9066\,
            I => \N__9037\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9063\,
            I => \N__9033\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__9060\,
            I => \N__9015\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9057\,
            I => \N__9009\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9054\,
            I => \N__9000\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__9051\,
            I => \N__8995\
        );

    \I__2115\ : SRMux
    port map (
            O => \N__9050\,
            I => \N__8906\
        );

    \I__2114\ : Glb2LocalMux
    port map (
            O => \N__9047\,
            I => \N__8906\
        );

    \I__2113\ : SRMux
    port map (
            O => \N__9046\,
            I => \N__8906\
        );

    \I__2112\ : Glb2LocalMux
    port map (
            O => \N__9043\,
            I => \N__8906\
        );

    \I__2111\ : Glb2LocalMux
    port map (
            O => \N__9040\,
            I => \N__8906\
        );

    \I__2110\ : Glb2LocalMux
    port map (
            O => \N__9037\,
            I => \N__8906\
        );

    \I__2109\ : SRMux
    port map (
            O => \N__9036\,
            I => \N__8906\
        );

    \I__2108\ : Glb2LocalMux
    port map (
            O => \N__9033\,
            I => \N__8906\
        );

    \I__2107\ : SRMux
    port map (
            O => \N__9032\,
            I => \N__8906\
        );

    \I__2106\ : SRMux
    port map (
            O => \N__9031\,
            I => \N__8906\
        );

    \I__2105\ : SRMux
    port map (
            O => \N__9030\,
            I => \N__8906\
        );

    \I__2104\ : SRMux
    port map (
            O => \N__9029\,
            I => \N__8906\
        );

    \I__2103\ : SRMux
    port map (
            O => \N__9028\,
            I => \N__8906\
        );

    \I__2102\ : SRMux
    port map (
            O => \N__9027\,
            I => \N__8906\
        );

    \I__2101\ : SRMux
    port map (
            O => \N__9026\,
            I => \N__8906\
        );

    \I__2100\ : SRMux
    port map (
            O => \N__9025\,
            I => \N__8906\
        );

    \I__2099\ : SRMux
    port map (
            O => \N__9024\,
            I => \N__8906\
        );

    \I__2098\ : SRMux
    port map (
            O => \N__9023\,
            I => \N__8906\
        );

    \I__2097\ : SRMux
    port map (
            O => \N__9022\,
            I => \N__8906\
        );

    \I__2096\ : SRMux
    port map (
            O => \N__9021\,
            I => \N__8906\
        );

    \I__2095\ : SRMux
    port map (
            O => \N__9020\,
            I => \N__8906\
        );

    \I__2094\ : SRMux
    port map (
            O => \N__9019\,
            I => \N__8906\
        );

    \I__2093\ : SRMux
    port map (
            O => \N__9018\,
            I => \N__8906\
        );

    \I__2092\ : Glb2LocalMux
    port map (
            O => \N__9015\,
            I => \N__8906\
        );

    \I__2091\ : SRMux
    port map (
            O => \N__9014\,
            I => \N__8906\
        );

    \I__2090\ : SRMux
    port map (
            O => \N__9013\,
            I => \N__8906\
        );

    \I__2089\ : SRMux
    port map (
            O => \N__9012\,
            I => \N__8906\
        );

    \I__2088\ : Glb2LocalMux
    port map (
            O => \N__9009\,
            I => \N__8906\
        );

    \I__2087\ : SRMux
    port map (
            O => \N__9008\,
            I => \N__8906\
        );

    \I__2086\ : SRMux
    port map (
            O => \N__9007\,
            I => \N__8906\
        );

    \I__2085\ : SRMux
    port map (
            O => \N__9006\,
            I => \N__8906\
        );

    \I__2084\ : SRMux
    port map (
            O => \N__9005\,
            I => \N__8906\
        );

    \I__2083\ : SRMux
    port map (
            O => \N__9004\,
            I => \N__8906\
        );

    \I__2082\ : SRMux
    port map (
            O => \N__9003\,
            I => \N__8906\
        );

    \I__2081\ : Glb2LocalMux
    port map (
            O => \N__9000\,
            I => \N__8906\
        );

    \I__2080\ : SRMux
    port map (
            O => \N__8999\,
            I => \N__8906\
        );

    \I__2079\ : SRMux
    port map (
            O => \N__8998\,
            I => \N__8906\
        );

    \I__2078\ : Glb2LocalMux
    port map (
            O => \N__8995\,
            I => \N__8906\
        );

    \I__2077\ : SRMux
    port map (
            O => \N__8994\,
            I => \N__8906\
        );

    \I__2076\ : SRMux
    port map (
            O => \N__8993\,
            I => \N__8906\
        );

    \I__2075\ : SRMux
    port map (
            O => \N__8992\,
            I => \N__8906\
        );

    \I__2074\ : SRMux
    port map (
            O => \N__8991\,
            I => \N__8906\
        );

    \I__2073\ : GlobalMux
    port map (
            O => \N__8906\,
            I => \N__8903\
        );

    \I__2072\ : gio2CtrlBuf
    port map (
            O => \N__8903\,
            I => \RESETn_c_i_g\
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__8900\,
            I => \N__8897\
        );

    \I__2070\ : InMux
    port map (
            O => \N__8897\,
            I => \N__8894\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__8894\,
            I => \N__8889\
        );

    \I__2068\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8886\
        );

    \I__2067\ : InMux
    port map (
            O => \N__8892\,
            I => \N__8883\
        );

    \I__2066\ : Span4Mux_v
    port map (
            O => \N__8889\,
            I => \N__8878\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__8886\,
            I => \N__8878\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__8883\,
            I => \N__8875\
        );

    \I__2063\ : Span4Mux_h
    port map (
            O => \N__8878\,
            I => \N__8870\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__8875\,
            I => \N__8870\
        );

    \I__2061\ : Sp12to4
    port map (
            O => \N__8870\,
            I => \N__8867\
        );

    \I__2060\ : Span12Mux_v
    port map (
            O => \N__8867\,
            I => \N__8864\
        );

    \I__2059\ : Span12Mux_h
    port map (
            O => \N__8864\,
            I => \N__8861\
        );

    \I__2058\ : Odrv12
    port map (
            O => \N__8861\,
            I => \CASLn_c\
        );

    \I__2057\ : InMux
    port map (
            O => \N__8858\,
            I => \N__8854\
        );

    \I__2056\ : InMux
    port map (
            O => \N__8857\,
            I => \N__8850\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__8854\,
            I => \N__8847\
        );

    \I__2054\ : InMux
    port map (
            O => \N__8853\,
            I => \N__8844\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__8850\,
            I => \N__8841\
        );

    \I__2052\ : Span4Mux_h
    port map (
            O => \N__8847\,
            I => \N__8836\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__8844\,
            I => \N__8836\
        );

    \I__2050\ : Span4Mux_v
    port map (
            O => \N__8841\,
            I => \N__8833\
        );

    \I__2049\ : Span4Mux_v
    port map (
            O => \N__8836\,
            I => \N__8830\
        );

    \I__2048\ : Span4Mux_v
    port map (
            O => \N__8833\,
            I => \N__8827\
        );

    \I__2047\ : Sp12to4
    port map (
            O => \N__8830\,
            I => \N__8822\
        );

    \I__2046\ : Sp12to4
    port map (
            O => \N__8827\,
            I => \N__8822\
        );

    \I__2045\ : Span12Mux_h
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__2044\ : Span12Mux_v
    port map (
            O => \N__8819\,
            I => \N__8816\
        );

    \I__2043\ : Odrv12
    port map (
            O => \N__8816\,
            I => \CASUn_c\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__8813\,
            I => \N__8810\
        );

    \I__2041\ : InMux
    port map (
            O => \N__8810\,
            I => \N__8807\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__8807\,
            I => \N__8803\
        );

    \I__2039\ : InMux
    port map (
            O => \N__8806\,
            I => \N__8799\
        );

    \I__2038\ : Span4Mux_v
    port map (
            O => \N__8803\,
            I => \N__8796\
        );

    \I__2037\ : InMux
    port map (
            O => \N__8802\,
            I => \N__8793\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__8799\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__8796\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__8793\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__2033\ : InMux
    port map (
            O => \N__8786\,
            I => \N__8783\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__8783\,
            I => \N__8780\
        );

    \I__2031\ : Span4Mux_h
    port map (
            O => \N__8780\,
            I => \N__8776\
        );

    \I__2030\ : InMux
    port map (
            O => \N__8779\,
            I => \N__8773\
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__8776\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__8773\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__2027\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8764\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__8767\,
            I => \N__8761\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__8764\,
            I => \N__8750\
        );

    \I__2024\ : InMux
    port map (
            O => \N__8761\,
            I => \N__8744\
        );

    \I__2023\ : InMux
    port map (
            O => \N__8760\,
            I => \N__8744\
        );

    \I__2022\ : InMux
    port map (
            O => \N__8759\,
            I => \N__8741\
        );

    \I__2021\ : InMux
    port map (
            O => \N__8758\,
            I => \N__8736\
        );

    \I__2020\ : InMux
    port map (
            O => \N__8757\,
            I => \N__8736\
        );

    \I__2019\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8731\
        );

    \I__2018\ : InMux
    port map (
            O => \N__8755\,
            I => \N__8731\
        );

    \I__2017\ : InMux
    port map (
            O => \N__8754\,
            I => \N__8728\
        );

    \I__2016\ : InMux
    port map (
            O => \N__8753\,
            I => \N__8725\
        );

    \I__2015\ : Span4Mux_h
    port map (
            O => \N__8750\,
            I => \N__8722\
        );

    \I__2014\ : InMux
    port map (
            O => \N__8749\,
            I => \N__8719\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__8744\,
            I => \N__8714\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__8741\,
            I => \N__8709\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__8736\,
            I => \N__8709\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__8731\,
            I => \N__8706\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__8728\,
            I => \N__8697\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__8725\,
            I => \N__8697\
        );

    \I__2007\ : Span4Mux_v
    port map (
            O => \N__8722\,
            I => \N__8697\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__8719\,
            I => \N__8697\
        );

    \I__2005\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8693\
        );

    \I__2004\ : InMux
    port map (
            O => \N__8717\,
            I => \N__8690\
        );

    \I__2003\ : Span4Mux_v
    port map (
            O => \N__8714\,
            I => \N__8687\
        );

    \I__2002\ : Span12Mux_h
    port map (
            O => \N__8709\,
            I => \N__8684\
        );

    \I__2001\ : Span4Mux_h
    port map (
            O => \N__8706\,
            I => \N__8679\
        );

    \I__2000\ : Span4Mux_h
    port map (
            O => \N__8697\,
            I => \N__8679\
        );

    \I__1999\ : InMux
    port map (
            O => \N__8696\,
            I => \N__8676\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__8693\,
            I => \N__8673\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__8690\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1996\ : Odrv4
    port map (
            O => \N__8687\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1995\ : Odrv12
    port map (
            O => \N__8684\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__8679\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__8676\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__8673\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1991\ : IoInMux
    port map (
            O => \N__8660\,
            I => \N__8657\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__8657\,
            I => \N__8654\
        );

    \I__1989\ : Span4Mux_s2_v
    port map (
            O => \N__8654\,
            I => \N__8651\
        );

    \I__1988\ : Span4Mux_v
    port map (
            O => \N__8651\,
            I => \N__8648\
        );

    \I__1987\ : Span4Mux_h
    port map (
            O => \N__8648\,
            I => \N__8645\
        );

    \I__1986\ : Odrv4
    port map (
            O => \N__8645\,
            I => \RASn_c\
        );

    \I__1985\ : InMux
    port map (
            O => \N__8642\,
            I => \N__8635\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__8641\,
            I => \N__8632\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__8640\,
            I => \N__8628\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__8639\,
            I => \N__8624\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__8638\,
            I => \N__8621\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__8635\,
            I => \N__8616\
        );

    \I__1979\ : InMux
    port map (
            O => \N__8632\,
            I => \N__8609\
        );

    \I__1978\ : InMux
    port map (
            O => \N__8631\,
            I => \N__8609\
        );

    \I__1977\ : InMux
    port map (
            O => \N__8628\,
            I => \N__8604\
        );

    \I__1976\ : InMux
    port map (
            O => \N__8627\,
            I => \N__8604\
        );

    \I__1975\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8597\
        );

    \I__1974\ : InMux
    port map (
            O => \N__8621\,
            I => \N__8597\
        );

    \I__1973\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8597\
        );

    \I__1972\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8594\
        );

    \I__1971\ : Span4Mux_h
    port map (
            O => \N__8616\,
            I => \N__8591\
        );

    \I__1970\ : InMux
    port map (
            O => \N__8615\,
            I => \N__8586\
        );

    \I__1969\ : InMux
    port map (
            O => \N__8614\,
            I => \N__8586\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__8609\,
            I => \N__8583\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__8604\,
            I => \N__8580\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__8597\,
            I => \N__8577\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__8594\,
            I => \N__8570\
        );

    \I__1964\ : Span4Mux_v
    port map (
            O => \N__8591\,
            I => \N__8570\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__8586\,
            I => \N__8570\
        );

    \I__1962\ : Span4Mux_v
    port map (
            O => \N__8583\,
            I => \N__8563\
        );

    \I__1961\ : Span4Mux_v
    port map (
            O => \N__8580\,
            I => \N__8563\
        );

    \I__1960\ : Span4Mux_v
    port map (
            O => \N__8577\,
            I => \N__8560\
        );

    \I__1959\ : Span4Mux_h
    port map (
            O => \N__8570\,
            I => \N__8557\
        );

    \I__1958\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8552\
        );

    \I__1957\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8552\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__8563\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1955\ : Odrv4
    port map (
            O => \N__8560\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__8557\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__8552\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1952\ : IoInMux
    port map (
            O => \N__8543\,
            I => \N__8540\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__8540\,
            I => \N__8537\
        );

    \I__1950\ : IoSpan4Mux
    port map (
            O => \N__8537\,
            I => \N__8534\
        );

    \I__1949\ : IoSpan4Mux
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__1948\ : Span4Mux_s1_h
    port map (
            O => \N__8531\,
            I => \N__8528\
        );

    \I__1947\ : Sp12to4
    port map (
            O => \N__8528\,
            I => \N__8525\
        );

    \I__1946\ : Odrv12
    port map (
            O => \N__8525\,
            I => \WEn_c\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8515\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__8521\,
            I => \N__8511\
        );

    \I__1943\ : InMux
    port map (
            O => \N__8520\,
            I => \N__8508\
        );

    \I__1942\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8497\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8518\,
            I => \N__8497\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__8515\,
            I => \N__8493\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__8514\,
            I => \N__8490\
        );

    \I__1938\ : InMux
    port map (
            O => \N__8511\,
            I => \N__8487\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__8508\,
            I => \N__8484\
        );

    \I__1936\ : InMux
    port map (
            O => \N__8507\,
            I => \N__8481\
        );

    \I__1935\ : InMux
    port map (
            O => \N__8506\,
            I => \N__8477\
        );

    \I__1934\ : InMux
    port map (
            O => \N__8505\,
            I => \N__8472\
        );

    \I__1933\ : InMux
    port map (
            O => \N__8504\,
            I => \N__8472\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8503\,
            I => \N__8465\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8502\,
            I => \N__8465\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__8497\,
            I => \N__8462\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8459\
        );

    \I__1928\ : Span4Mux_v
    port map (
            O => \N__8493\,
            I => \N__8456\
        );

    \I__1927\ : InMux
    port map (
            O => \N__8490\,
            I => \N__8453\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__8487\,
            I => \N__8446\
        );

    \I__1925\ : Span4Mux_h
    port map (
            O => \N__8484\,
            I => \N__8446\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8481\,
            I => \N__8446\
        );

    \I__1923\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8443\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__8477\,
            I => \N__8438\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__8472\,
            I => \N__8438\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8471\,
            I => \N__8435\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__8470\,
            I => \N__8432\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__8465\,
            I => \N__8429\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__8462\,
            I => \N__8420\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__8459\,
            I => \N__8420\
        );

    \I__1915\ : Span4Mux_h
    port map (
            O => \N__8456\,
            I => \N__8420\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__8453\,
            I => \N__8420\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__8446\,
            I => \N__8417\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__8443\,
            I => \N__8410\
        );

    \I__1911\ : Span4Mux_v
    port map (
            O => \N__8438\,
            I => \N__8410\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__8435\,
            I => \N__8410\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8432\,
            I => \N__8407\
        );

    \I__1908\ : Odrv4
    port map (
            O => \N__8429\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__8420\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__8417\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1905\ : Odrv4
    port map (
            O => \N__8410\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8407\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1903\ : IoInMux
    port map (
            O => \N__8396\,
            I => \N__8393\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__8393\,
            I => \N__8390\
        );

    \I__1901\ : Span4Mux_s1_v
    port map (
            O => \N__8390\,
            I => \N__8387\
        );

    \I__1900\ : Sp12to4
    port map (
            O => \N__8387\,
            I => \N__8384\
        );

    \I__1899\ : Span12Mux_h
    port map (
            O => \N__8384\,
            I => \N__8381\
        );

    \I__1898\ : Odrv12
    port map (
            O => \N__8381\,
            I => \CASn_c\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8378\,
            I => \N__8374\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8371\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__8374\,
            I => \N__8368\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__8371\,
            I => \N__8365\
        );

    \I__1893\ : Span4Mux_v
    port map (
            O => \N__8368\,
            I => \N__8362\
        );

    \I__1892\ : Span4Mux_h
    port map (
            O => \N__8365\,
            I => \N__8359\
        );

    \I__1891\ : Span4Mux_v
    port map (
            O => \N__8362\,
            I => \N__8356\
        );

    \I__1890\ : Span4Mux_v
    port map (
            O => \N__8359\,
            I => \N__8353\
        );

    \I__1889\ : Sp12to4
    port map (
            O => \N__8356\,
            I => \N__8348\
        );

    \I__1888\ : Sp12to4
    port map (
            O => \N__8353\,
            I => \N__8348\
        );

    \I__1887\ : Span12Mux_h
    port map (
            O => \N__8348\,
            I => \N__8345\
        );

    \I__1886\ : Odrv12
    port map (
            O => \N__8345\,
            I => \RAS0n_c\
        );

    \I__1885\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8339\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__8339\,
            I => \N__8336\
        );

    \I__1883\ : Span12Mux_v
    port map (
            O => \N__8336\,
            I => \N__8333\
        );

    \I__1882\ : Span12Mux_h
    port map (
            O => \N__8333\,
            I => \N__8330\
        );

    \I__1881\ : Odrv12
    port map (
            O => \N__8330\,
            I => \RAS1n_c\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8327\,
            I => \N__8323\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8326\,
            I => \N__8320\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8323\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8320\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__1876\ : InMux
    port map (
            O => \N__8315\,
            I => \N__8312\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8312\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8309\,
            I => \N__8305\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8308\,
            I => \N__8302\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8305\,
            I => \N__8299\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8302\,
            I => \N__8296\
        );

    \I__1870\ : Span4Mux_v
    port map (
            O => \N__8299\,
            I => \N__8293\
        );

    \I__1869\ : Span4Mux_v
    port map (
            O => \N__8296\,
            I => \N__8290\
        );

    \I__1868\ : Span4Mux_v
    port map (
            O => \N__8293\,
            I => \N__8287\
        );

    \I__1867\ : Span4Mux_v
    port map (
            O => \N__8290\,
            I => \N__8284\
        );

    \I__1866\ : Sp12to4
    port map (
            O => \N__8287\,
            I => \N__8279\
        );

    \I__1865\ : Sp12to4
    port map (
            O => \N__8284\,
            I => \N__8279\
        );

    \I__1864\ : Span12Mux_h
    port map (
            O => \N__8279\,
            I => \N__8276\
        );

    \I__1863\ : Odrv12
    port map (
            O => \N__8276\,
            I => \DRA_c_7\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8273\,
            I => \N__8270\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8270\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8267\,
            I => \N__8264\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__8264\,
            I => \N__8261\
        );

    \I__1858\ : Sp12to4
    port map (
            O => \N__8261\,
            I => \N__8258\
        );

    \I__1857\ : Span12Mux_v
    port map (
            O => \N__8258\,
            I => \N__8255\
        );

    \I__1856\ : Span12Mux_h
    port map (
            O => \N__8255\,
            I => \N__8252\
        );

    \I__1855\ : Odrv12
    port map (
            O => \N__8252\,
            I => \A_c_18\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__8249\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8246\,
            I => \N__8243\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__8243\,
            I => \N__8240\
        );

    \I__1851\ : Sp12to4
    port map (
            O => \N__8240\,
            I => \N__8237\
        );

    \I__1850\ : Span12Mux_v
    port map (
            O => \N__8237\,
            I => \N__8234\
        );

    \I__1849\ : Span12Mux_h
    port map (
            O => \N__8234\,
            I => \N__8231\
        );

    \I__1848\ : Odrv12
    port map (
            O => \N__8231\,
            I => \A_c_16\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__8228\,
            I => \U712_CHIP_RAM.N_322_cascade_\
        );

    \I__1846\ : IoInMux
    port map (
            O => \N__8225\,
            I => \N__8222\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8222\,
            I => \N__8219\
        );

    \I__1844\ : Span4Mux_s2_h
    port map (
            O => \N__8219\,
            I => \N__8216\
        );

    \I__1843\ : Span4Mux_v
    port map (
            O => \N__8216\,
            I => \N__8213\
        );

    \I__1842\ : Sp12to4
    port map (
            O => \N__8213\,
            I => \N__8210\
        );

    \I__1841\ : Span12Mux_h
    port map (
            O => \N__8210\,
            I => \N__8207\
        );

    \I__1840\ : Odrv12
    port map (
            O => \N__8207\,
            I => \CMA_c_7\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8204\,
            I => \N__8201\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8201\,
            I => \U712_CHIP_RAM.CMA_5_i_0_8\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8198\,
            I => \N__8195\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__8195\,
            I => \N__8192\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__8192\,
            I => \N__8189\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__8189\,
            I => \N__8186\
        );

    \I__1833\ : Sp12to4
    port map (
            O => \N__8186\,
            I => \N__8183\
        );

    \I__1832\ : Span12Mux_h
    port map (
            O => \N__8183\,
            I => \N__8180\
        );

    \I__1831\ : Odrv12
    port map (
            O => \N__8180\,
            I => \A_c_19\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__8177\,
            I => \U712_CHIP_RAM.CMA_5_i_0_8_cascade_\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__8174\,
            I => \N__8170\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__8173\,
            I => \N__8163\
        );

    \I__1827\ : InMux
    port map (
            O => \N__8170\,
            I => \N__8159\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__8169\,
            I => \N__8155\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__8168\,
            I => \N__8152\
        );

    \I__1824\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8141\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8166\,
            I => \N__8141\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8138\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8162\,
            I => \N__8129\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8159\,
            I => \N__8126\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8158\,
            I => \N__8123\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8120\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8115\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8151\,
            I => \N__8115\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8150\,
            I => \N__8108\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8149\,
            I => \N__8108\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8148\,
            I => \N__8108\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__8147\,
            I => \N__8103\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__8146\,
            I => \N__8100\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8141\,
            I => \N__8094\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__8138\,
            I => \N__8094\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8137\,
            I => \N__8089\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8136\,
            I => \N__8086\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8135\,
            I => \N__8081\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8134\,
            I => \N__8081\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__8133\,
            I => \N__8077\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8132\,
            I => \N__8073\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8129\,
            I => \N__8064\
        );

    \I__1801\ : Span4Mux_v
    port map (
            O => \N__8126\,
            I => \N__8064\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__8123\,
            I => \N__8064\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8120\,
            I => \N__8064\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8115\,
            I => \N__8056\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8108\,
            I => \N__8056\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8107\,
            I => \N__8051\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8106\,
            I => \N__8051\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8046\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8100\,
            I => \N__8046\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8043\
        );

    \I__1791\ : Span4Mux_h
    port map (
            O => \N__8094\,
            I => \N__8040\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8093\,
            I => \N__8035\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8092\,
            I => \N__8035\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8089\,
            I => \N__8028\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__8086\,
            I => \N__8028\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8081\,
            I => \N__8028\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8080\,
            I => \N__8021\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8077\,
            I => \N__8021\
        );

    \I__1783\ : InMux
    port map (
            O => \N__8076\,
            I => \N__8021\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8073\,
            I => \N__8016\
        );

    \I__1781\ : Span4Mux_h
    port map (
            O => \N__8064\,
            I => \N__8016\
        );

    \I__1780\ : InMux
    port map (
            O => \N__8063\,
            I => \N__8009\
        );

    \I__1779\ : InMux
    port map (
            O => \N__8062\,
            I => \N__8009\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8061\,
            I => \N__8009\
        );

    \I__1777\ : Odrv12
    port map (
            O => \N__8056\,
            I => \CPU_CYCLEm\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__8051\,
            I => \CPU_CYCLEm\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__8046\,
            I => \CPU_CYCLEm\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__8043\,
            I => \CPU_CYCLEm\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__8040\,
            I => \CPU_CYCLEm\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8035\,
            I => \CPU_CYCLEm\
        );

    \I__1771\ : Odrv12
    port map (
            O => \N__8028\,
            I => \CPU_CYCLEm\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8021\,
            I => \CPU_CYCLEm\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__8016\,
            I => \CPU_CYCLEm\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8009\,
            I => \CPU_CYCLEm\
        );

    \I__1767\ : IoInMux
    port map (
            O => \N__7988\,
            I => \N__7985\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__7985\,
            I => \N__7982\
        );

    \I__1765\ : IoSpan4Mux
    port map (
            O => \N__7982\,
            I => \N__7979\
        );

    \I__1764\ : Span4Mux_s2_h
    port map (
            O => \N__7979\,
            I => \N__7976\
        );

    \I__1763\ : Sp12to4
    port map (
            O => \N__7976\,
            I => \N__7973\
        );

    \I__1762\ : Span12Mux_h
    port map (
            O => \N__7973\,
            I => \N__7970\
        );

    \I__1761\ : Odrv12
    port map (
            O => \N__7970\,
            I => \CMA_c_9\
        );

    \I__1760\ : CEMux
    port map (
            O => \N__7967\,
            I => \N__7961\
        );

    \I__1759\ : CEMux
    port map (
            O => \N__7966\,
            I => \N__7958\
        );

    \I__1758\ : CEMux
    port map (
            O => \N__7965\,
            I => \N__7955\
        );

    \I__1757\ : CEMux
    port map (
            O => \N__7964\,
            I => \N__7952\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__7961\,
            I => \N__7948\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__7958\,
            I => \N__7945\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__7955\,
            I => \N__7942\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__7952\,
            I => \N__7939\
        );

    \I__1752\ : CEMux
    port map (
            O => \N__7951\,
            I => \N__7936\
        );

    \I__1751\ : Span4Mux_h
    port map (
            O => \N__7948\,
            I => \N__7931\
        );

    \I__1750\ : Span4Mux_h
    port map (
            O => \N__7945\,
            I => \N__7931\
        );

    \I__1749\ : Span4Mux_v
    port map (
            O => \N__7942\,
            I => \N__7928\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__7939\,
            I => \N__7923\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__7936\,
            I => \N__7923\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__7931\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__7928\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__7923\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1743\ : InMux
    port map (
            O => \N__7916\,
            I => \N__7913\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__7913\,
            I => \N__7910\
        );

    \I__1741\ : Odrv12
    port map (
            O => \N__7910\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1740\ : InMux
    port map (
            O => \N__7907\,
            I => \N__7903\
        );

    \I__1739\ : InMux
    port map (
            O => \N__7906\,
            I => \N__7900\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__7903\,
            I => \N__7895\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__7900\,
            I => \N__7895\
        );

    \I__1736\ : Span4Mux_v
    port map (
            O => \N__7895\,
            I => \N__7892\
        );

    \I__1735\ : Sp12to4
    port map (
            O => \N__7892\,
            I => \N__7889\
        );

    \I__1734\ : Span12Mux_h
    port map (
            O => \N__7889\,
            I => \N__7886\
        );

    \I__1733\ : Span12Mux_v
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__1732\ : Odrv12
    port map (
            O => \N__7883\,
            I => \DRA_c_4\
        );

    \I__1731\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7877\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__7877\,
            I => \N__7874\
        );

    \I__1729\ : Odrv12
    port map (
            O => \N__7874\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1728\ : InMux
    port map (
            O => \N__7871\,
            I => \N__7868\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__7868\,
            I => \N__7864\
        );

    \I__1726\ : InMux
    port map (
            O => \N__7867\,
            I => \N__7861\
        );

    \I__1725\ : Span4Mux_v
    port map (
            O => \N__7864\,
            I => \N__7856\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__7861\,
            I => \N__7856\
        );

    \I__1723\ : Span4Mux_v
    port map (
            O => \N__7856\,
            I => \N__7853\
        );

    \I__1722\ : Sp12to4
    port map (
            O => \N__7853\,
            I => \N__7850\
        );

    \I__1721\ : Span12Mux_h
    port map (
            O => \N__7850\,
            I => \N__7847\
        );

    \I__1720\ : Odrv12
    port map (
            O => \N__7847\,
            I => \DRA_c_8\
        );

    \I__1719\ : InMux
    port map (
            O => \N__7844\,
            I => \N__7841\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__7841\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1717\ : CEMux
    port map (
            O => \N__7838\,
            I => \N__7834\
        );

    \I__1716\ : CEMux
    port map (
            O => \N__7837\,
            I => \N__7829\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__7834\,
            I => \N__7826\
        );

    \I__1714\ : CEMux
    port map (
            O => \N__7833\,
            I => \N__7823\
        );

    \I__1713\ : CEMux
    port map (
            O => \N__7832\,
            I => \N__7820\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__7829\,
            I => \N__7817\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__7826\,
            I => \N__7814\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__7823\,
            I => \N__7809\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__7820\,
            I => \N__7809\
        );

    \I__1708\ : Span4Mux_h
    port map (
            O => \N__7817\,
            I => \N__7804\
        );

    \I__1707\ : Span4Mux_h
    port map (
            O => \N__7814\,
            I => \N__7804\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__7809\,
            I => \N__7801\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__7804\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__7801\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1703\ : InMux
    port map (
            O => \N__7796\,
            I => \N__7791\
        );

    \I__1702\ : InMux
    port map (
            O => \N__7795\,
            I => \N__7786\
        );

    \I__1701\ : InMux
    port map (
            O => \N__7794\,
            I => \N__7786\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__7791\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__7786\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1698\ : InMux
    port map (
            O => \N__7781\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__1697\ : InMux
    port map (
            O => \N__7778\,
            I => \N__7774\
        );

    \I__1696\ : InMux
    port map (
            O => \N__7777\,
            I => \N__7771\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__7774\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__7771\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1693\ : InMux
    port map (
            O => \N__7766\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__1692\ : InMux
    port map (
            O => \N__7763\,
            I => \N__7759\
        );

    \I__1691\ : InMux
    port map (
            O => \N__7762\,
            I => \N__7756\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__7759\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__7756\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1688\ : InMux
    port map (
            O => \N__7751\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__1687\ : InMux
    port map (
            O => \N__7748\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__1686\ : InMux
    port map (
            O => \N__7745\,
            I => \N__7740\
        );

    \I__1685\ : InMux
    port map (
            O => \N__7744\,
            I => \N__7735\
        );

    \I__1684\ : InMux
    port map (
            O => \N__7743\,
            I => \N__7735\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__7740\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__7735\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1681\ : ClkMux
    port map (
            O => \N__7730\,
            I => \N__7727\
        );

    \I__1680\ : GlobalMux
    port map (
            O => \N__7727\,
            I => \N__7724\
        );

    \I__1679\ : gio2CtrlBuf
    port map (
            O => \N__7724\,
            I => \C1_c_g\
        );

    \I__1678\ : SRMux
    port map (
            O => \N__7721\,
            I => \N__7718\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__7718\,
            I => \N__7715\
        );

    \I__1676\ : Span4Mux_h
    port map (
            O => \N__7715\,
            I => \N__7712\
        );

    \I__1675\ : Odrv4
    port map (
            O => \N__7712\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1674\ : InMux
    port map (
            O => \N__7709\,
            I => \N__7703\
        );

    \I__1673\ : InMux
    port map (
            O => \N__7708\,
            I => \N__7703\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__7703\,
            I => \N__7698\
        );

    \I__1671\ : InMux
    port map (
            O => \N__7702\,
            I => \N__7695\
        );

    \I__1670\ : InMux
    port map (
            O => \N__7701\,
            I => \N__7692\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__7698\,
            I => \N__7686\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__7695\,
            I => \N__7686\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__7692\,
            I => \N__7682\
        );

    \I__1666\ : InMux
    port map (
            O => \N__7691\,
            I => \N__7679\
        );

    \I__1665\ : Span4Mux_h
    port map (
            O => \N__7686\,
            I => \N__7676\
        );

    \I__1664\ : InMux
    port map (
            O => \N__7685\,
            I => \N__7673\
        );

    \I__1663\ : Span4Mux_v
    port map (
            O => \N__7682\,
            I => \N__7670\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7679\,
            I => \N__7667\
        );

    \I__1661\ : Span4Mux_v
    port map (
            O => \N__7676\,
            I => \N__7664\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7673\,
            I => \N__7661\
        );

    \I__1659\ : Sp12to4
    port map (
            O => \N__7670\,
            I => \N__7658\
        );

    \I__1658\ : Span12Mux_h
    port map (
            O => \N__7667\,
            I => \N__7655\
        );

    \I__1657\ : Sp12to4
    port map (
            O => \N__7664\,
            I => \N__7650\
        );

    \I__1656\ : Span12Mux_v
    port map (
            O => \N__7661\,
            I => \N__7650\
        );

    \I__1655\ : Span12Mux_h
    port map (
            O => \N__7658\,
            I => \N__7647\
        );

    \I__1654\ : Span12Mux_h
    port map (
            O => \N__7655\,
            I => \N__7644\
        );

    \I__1653\ : Span12Mux_h
    port map (
            O => \N__7650\,
            I => \N__7641\
        );

    \I__1652\ : Odrv12
    port map (
            O => \N__7647\,
            I => \RESETn_c\
        );

    \I__1651\ : Odrv12
    port map (
            O => \N__7644\,
            I => \RESETn_c\
        );

    \I__1650\ : Odrv12
    port map (
            O => \N__7641\,
            I => \RESETn_c\
        );

    \I__1649\ : IoInMux
    port map (
            O => \N__7634\,
            I => \N__7631\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__7631\,
            I => \N__7628\
        );

    \I__1647\ : Span12Mux_s7_v
    port map (
            O => \N__7628\,
            I => \N__7625\
        );

    \I__1646\ : Odrv12
    port map (
            O => \N__7625\,
            I => \RESETn_c_i\
        );

    \I__1645\ : InMux
    port map (
            O => \N__7622\,
            I => \N__7619\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7619\,
            I => \N__7615\
        );

    \I__1643\ : InMux
    port map (
            O => \N__7618\,
            I => \N__7612\
        );

    \I__1642\ : Span4Mux_h
    port map (
            O => \N__7615\,
            I => \N__7609\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7612\,
            I => \N__7606\
        );

    \I__1640\ : Sp12to4
    port map (
            O => \N__7609\,
            I => \N__7601\
        );

    \I__1639\ : Sp12to4
    port map (
            O => \N__7606\,
            I => \N__7601\
        );

    \I__1638\ : Span12Mux_v
    port map (
            O => \N__7601\,
            I => \N__7598\
        );

    \I__1637\ : Span12Mux_h
    port map (
            O => \N__7598\,
            I => \N__7595\
        );

    \I__1636\ : Odrv12
    port map (
            O => \N__7595\,
            I => \DRA_c_5\
        );

    \I__1635\ : InMux
    port map (
            O => \N__7592\,
            I => \N__7589\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__7589\,
            I => \N__7586\
        );

    \I__1633\ : Odrv4
    port map (
            O => \N__7586\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1632\ : InMux
    port map (
            O => \N__7583\,
            I => \N__7580\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__7580\,
            I => \N__7577\
        );

    \I__1630\ : Odrv12
    port map (
            O => \N__7577\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__1629\ : CascadeMux
    port map (
            O => \N__7574\,
            I => \N__7571\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7568\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__7568\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1626\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7561\
        );

    \I__1625\ : InMux
    port map (
            O => \N__7564\,
            I => \N__7558\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7561\,
            I => \N__7553\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7558\,
            I => \N__7553\
        );

    \I__1622\ : Span4Mux_v
    port map (
            O => \N__7553\,
            I => \N__7550\
        );

    \I__1621\ : Sp12to4
    port map (
            O => \N__7550\,
            I => \N__7547\
        );

    \I__1620\ : Span12Mux_h
    port map (
            O => \N__7547\,
            I => \N__7544\
        );

    \I__1619\ : Span12Mux_v
    port map (
            O => \N__7544\,
            I => \N__7541\
        );

    \I__1618\ : Odrv12
    port map (
            O => \N__7541\,
            I => \DRA_c_6\
        );

    \I__1617\ : InMux
    port map (
            O => \N__7538\,
            I => \N__7535\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__7535\,
            I => \N__7532\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__7532\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__1614\ : InMux
    port map (
            O => \N__7529\,
            I => \N__7526\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__7526\,
            I => \N__7522\
        );

    \I__1612\ : InMux
    port map (
            O => \N__7525\,
            I => \N__7519\
        );

    \I__1611\ : Span4Mux_h
    port map (
            O => \N__7522\,
            I => \N__7514\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__7519\,
            I => \N__7514\
        );

    \I__1609\ : Span4Mux_v
    port map (
            O => \N__7514\,
            I => \N__7511\
        );

    \I__1608\ : Sp12to4
    port map (
            O => \N__7511\,
            I => \N__7508\
        );

    \I__1607\ : Span12Mux_h
    port map (
            O => \N__7508\,
            I => \N__7505\
        );

    \I__1606\ : Span12Mux_v
    port map (
            O => \N__7505\,
            I => \N__7502\
        );

    \I__1605\ : Odrv12
    port map (
            O => \N__7502\,
            I => \DRA_c_1\
        );

    \I__1604\ : InMux
    port map (
            O => \N__7499\,
            I => \N__7496\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__7496\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1602\ : InMux
    port map (
            O => \N__7493\,
            I => \N__7490\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__7490\,
            I => \N__7486\
        );

    \I__1600\ : InMux
    port map (
            O => \N__7489\,
            I => \N__7483\
        );

    \I__1599\ : Span4Mux_v
    port map (
            O => \N__7486\,
            I => \N__7480\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__7483\,
            I => \N__7475\
        );

    \I__1597\ : Sp12to4
    port map (
            O => \N__7480\,
            I => \N__7475\
        );

    \I__1596\ : Span12Mux_h
    port map (
            O => \N__7475\,
            I => \N__7472\
        );

    \I__1595\ : Span12Mux_v
    port map (
            O => \N__7472\,
            I => \N__7469\
        );

    \I__1594\ : Odrv12
    port map (
            O => \N__7469\,
            I => \DRA_c_3\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7466\,
            I => \N__7463\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__7463\,
            I => \N__7460\
        );

    \I__1591\ : Odrv12
    port map (
            O => \N__7460\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7457\,
            I => \N__7454\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7454\,
            I => \N__7450\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7453\,
            I => \N__7447\
        );

    \I__1587\ : Span4Mux_v
    port map (
            O => \N__7450\,
            I => \N__7444\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__7447\,
            I => \N__7441\
        );

    \I__1585\ : Sp12to4
    port map (
            O => \N__7444\,
            I => \N__7438\
        );

    \I__1584\ : Span12Mux_h
    port map (
            O => \N__7441\,
            I => \N__7435\
        );

    \I__1583\ : Span12Mux_h
    port map (
            O => \N__7438\,
            I => \N__7432\
        );

    \I__1582\ : Span12Mux_v
    port map (
            O => \N__7435\,
            I => \N__7429\
        );

    \I__1581\ : Span12Mux_v
    port map (
            O => \N__7432\,
            I => \N__7426\
        );

    \I__1580\ : Odrv12
    port map (
            O => \N__7429\,
            I => \DRA_c_2\
        );

    \I__1579\ : Odrv12
    port map (
            O => \N__7426\,
            I => \DRA_c_2\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__7421\,
            I => \N__7418\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7418\,
            I => \N__7415\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__7415\,
            I => \N__7412\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__7412\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1574\ : IoInMux
    port map (
            O => \N__7409\,
            I => \N__7406\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7406\,
            I => \N__7403\
        );

    \I__1572\ : Span4Mux_s3_v
    port map (
            O => \N__7403\,
            I => \N__7400\
        );

    \I__1571\ : Span4Mux_v
    port map (
            O => \N__7400\,
            I => \N__7397\
        );

    \I__1570\ : Span4Mux_v
    port map (
            O => \N__7397\,
            I => \N__7394\
        );

    \I__1569\ : Span4Mux_h
    port map (
            O => \N__7394\,
            I => \N__7390\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7393\,
            I => \N__7387\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__7390\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7387\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7382\,
            I => \N__7379\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__7379\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7376\,
            I => \bfn_12_8_0_\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7373\,
            I => \N__7370\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7370\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7367\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__1559\ : InMux
    port map (
            O => \N__7364\,
            I => \N__7359\
        );

    \I__1558\ : InMux
    port map (
            O => \N__7363\,
            I => \N__7354\
        );

    \I__1557\ : InMux
    port map (
            O => \N__7362\,
            I => \N__7354\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7359\,
            I => \U712_CHIP_RAM.REFRESH9lto2\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7354\,
            I => \U712_CHIP_RAM.REFRESH9lto2\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7349\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__1553\ : CascadeMux
    port map (
            O => \N__7346\,
            I => \N__7342\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7345\,
            I => \N__7338\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7342\,
            I => \N__7333\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7341\,
            I => \N__7333\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7338\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7333\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7328\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7322\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7322\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7316\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__7316\,
            I => \U712_CHIP_RAM.N_321\
        );

    \I__1542\ : IoInMux
    port map (
            O => \N__7313\,
            I => \N__7310\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__7310\,
            I => \N__7307\
        );

    \I__1540\ : Span4Mux_s0_h
    port map (
            O => \N__7307\,
            I => \N__7304\
        );

    \I__1539\ : Sp12to4
    port map (
            O => \N__7304\,
            I => \N__7301\
        );

    \I__1538\ : Span12Mux_s9_v
    port map (
            O => \N__7301\,
            I => \N__7298\
        );

    \I__1537\ : Span12Mux_h
    port map (
            O => \N__7298\,
            I => \N__7295\
        );

    \I__1536\ : Odrv12
    port map (
            O => \N__7295\,
            I => \CMA_c_6\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7292\,
            I => \N__7289\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7289\,
            I => \U712_CHIP_RAM.N_320\
        );

    \I__1533\ : IoInMux
    port map (
            O => \N__7286\,
            I => \N__7283\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__7283\,
            I => \N__7280\
        );

    \I__1531\ : Span12Mux_s4_h
    port map (
            O => \N__7280\,
            I => \N__7277\
        );

    \I__1530\ : Span12Mux_h
    port map (
            O => \N__7277\,
            I => \N__7274\
        );

    \I__1529\ : Odrv12
    port map (
            O => \N__7274\,
            I => \CMA_c_5\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7268\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7268\,
            I => \N__7265\
        );

    \I__1526\ : Span12Mux_v
    port map (
            O => \N__7265\,
            I => \N__7262\
        );

    \I__1525\ : Span12Mux_h
    port map (
            O => \N__7262\,
            I => \N__7259\
        );

    \I__1524\ : Odrv12
    port map (
            O => \N__7259\,
            I => \A_c_17\
        );

    \I__1523\ : IoInMux
    port map (
            O => \N__7256\,
            I => \N__7253\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7253\,
            I => \N__7250\
        );

    \I__1521\ : Span12Mux_s4_h
    port map (
            O => \N__7250\,
            I => \N__7247\
        );

    \I__1520\ : Span12Mux_h
    port map (
            O => \N__7247\,
            I => \N__7244\
        );

    \I__1519\ : Odrv12
    port map (
            O => \N__7244\,
            I => \CMA_c_8\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7241\,
            I => \N__7238\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__7238\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7235\,
            I => \N__7232\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__7232\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7229\,
            I => \N__7226\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7226\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7223\,
            I => \N__7220\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7220\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7217\,
            I => \N__7213\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7216\,
            I => \N__7210\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7213\,
            I => \U712_CHIP_RAM.N_425\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7210\,
            I => \U712_CHIP_RAM.N_425\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7205\,
            I => \N__7200\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7204\,
            I => \N__7197\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7203\,
            I => \N__7194\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7200\,
            I => \N__7190\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7197\,
            I => \N__7185\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7194\,
            I => \N__7182\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7174\
        );

    \I__1499\ : Span4Mux_v
    port map (
            O => \N__7190\,
            I => \N__7171\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7168\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7188\,
            I => \N__7165\
        );

    \I__1496\ : Span4Mux_v
    port map (
            O => \N__7185\,
            I => \N__7160\
        );

    \I__1495\ : Span4Mux_v
    port map (
            O => \N__7182\,
            I => \N__7160\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7181\,
            I => \N__7155\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7180\,
            I => \N__7155\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7179\,
            I => \N__7150\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7178\,
            I => \N__7150\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7177\,
            I => \N__7147\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7174\,
            I => \U712_CHIP_RAM.N_276\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__7171\,
            I => \U712_CHIP_RAM.N_276\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7168\,
            I => \U712_CHIP_RAM.N_276\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7165\,
            I => \U712_CHIP_RAM.N_276\
        );

    \I__1485\ : Odrv4
    port map (
            O => \N__7160\,
            I => \U712_CHIP_RAM.N_276\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7155\,
            I => \U712_CHIP_RAM.N_276\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7150\,
            I => \U712_CHIP_RAM.N_276\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7147\,
            I => \U712_CHIP_RAM.N_276\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7118\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7129\,
            I => \N__7118\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7128\,
            I => \N__7118\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7127\,
            I => \N__7115\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__7126\,
            I => \N__7109\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7125\,
            I => \N__7105\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__7118\,
            I => \N__7102\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7115\,
            I => \N__7099\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7114\,
            I => \N__7092\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7113\,
            I => \N__7092\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7112\,
            I => \N__7085\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7109\,
            I => \N__7085\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7108\,
            I => \N__7085\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7105\,
            I => \N__7078\
        );

    \I__1467\ : Span4Mux_v
    port map (
            O => \N__7102\,
            I => \N__7078\
        );

    \I__1466\ : Span4Mux_v
    port map (
            O => \N__7099\,
            I => \N__7078\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7098\,
            I => \N__7073\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7097\,
            I => \N__7073\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7092\,
            I => \N__7070\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7085\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1461\ : Odrv4
    port map (
            O => \N__7078\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__7073\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1459\ : Odrv12
    port map (
            O => \N__7070\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7061\,
            I => \N__7057\
        );

    \I__1457\ : InMux
    port map (
            O => \N__7060\,
            I => \N__7054\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7057\,
            I => \N__7051\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7054\,
            I => \N__7048\
        );

    \I__1454\ : Span4Mux_h
    port map (
            O => \N__7051\,
            I => \N__7045\
        );

    \I__1453\ : Span4Mux_h
    port map (
            O => \N__7048\,
            I => \N__7038\
        );

    \I__1452\ : Span4Mux_v
    port map (
            O => \N__7045\,
            I => \N__7038\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7044\,
            I => \N__7035\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7043\,
            I => \N__7032\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__7038\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7035\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7032\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1446\ : IoInMux
    port map (
            O => \N__7025\,
            I => \N__7022\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7022\,
            I => \N__7019\
        );

    \I__1444\ : Span4Mux_s3_v
    port map (
            O => \N__7019\,
            I => \N__7016\
        );

    \I__1443\ : Span4Mux_v
    port map (
            O => \N__7016\,
            I => \N__7013\
        );

    \I__1442\ : Span4Mux_v
    port map (
            O => \N__7013\,
            I => \N__7010\
        );

    \I__1441\ : Sp12to4
    port map (
            O => \N__7010\,
            I => \N__7007\
        );

    \I__1440\ : Odrv12
    port map (
            O => \N__7007\,
            I => \CRCSn_c\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7004\,
            I => \N__7001\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__7001\,
            I => \N__6997\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6994\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__6997\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_a2_0\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__6994\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_a2_0\
        );

    \I__1434\ : CascadeMux
    port map (
            O => \N__6989\,
            I => \N__6986\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6986\,
            I => \N__6983\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__6983\,
            I => \N__6980\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__6980\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__1430\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6972\
        );

    \I__1429\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6969\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6975\,
            I => \N__6966\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__6972\,
            I => \N__6959\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__6969\,
            I => \N__6956\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__6966\,
            I => \N__6951\
        );

    \I__1424\ : InMux
    port map (
            O => \N__6965\,
            I => \N__6946\
        );

    \I__1423\ : InMux
    port map (
            O => \N__6964\,
            I => \N__6946\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6963\,
            I => \N__6943\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6962\,
            I => \N__6940\
        );

    \I__1420\ : Span4Mux_v
    port map (
            O => \N__6959\,
            I => \N__6935\
        );

    \I__1419\ : Span4Mux_v
    port map (
            O => \N__6956\,
            I => \N__6935\
        );

    \I__1418\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6930\
        );

    \I__1417\ : InMux
    port map (
            O => \N__6954\,
            I => \N__6930\
        );

    \I__1416\ : Span4Mux_h
    port map (
            O => \N__6951\,
            I => \N__6925\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__6946\,
            I => \N__6925\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__6943\,
            I => \U712_CHIP_RAM.N_293\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__6940\,
            I => \U712_CHIP_RAM.N_293\
        );

    \I__1412\ : Odrv4
    port map (
            O => \N__6935\,
            I => \U712_CHIP_RAM.N_293\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6930\,
            I => \U712_CHIP_RAM.N_293\
        );

    \I__1410\ : Odrv4
    port map (
            O => \N__6925\,
            I => \U712_CHIP_RAM.N_293\
        );

    \I__1409\ : InMux
    port map (
            O => \N__6914\,
            I => \N__6909\
        );

    \I__1408\ : InMux
    port map (
            O => \N__6913\,
            I => \N__6906\
        );

    \I__1407\ : InMux
    port map (
            O => \N__6912\,
            I => \N__6903\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__6909\,
            I => \N__6898\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__6906\,
            I => \N__6898\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__6903\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__6898\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6890\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__6890\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__6887\,
            I => \U712_CHIP_RAM.REFRESH_RNO_0Z0Z_0_cascade_\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6884\,
            I => \N__6881\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6881\,
            I => \U712_CHIP_RAM.REFRESHZ0Z_0\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__6878\,
            I => \U712_CHIP_RAM.REFRESH9lt7_cascade_\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6875\,
            I => \N__6872\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__6872\,
            I => \N__6869\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__6869\,
            I => \U712_CHIP_RAM.REFRESHZ0Z_1\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6866\,
            I => \N__6860\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6865\,
            I => \N__6860\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6860\,
            I => \U712_CHIP_RAM.REFRESH9lto7_0\
        );

    \I__1390\ : InMux
    port map (
            O => \N__6857\,
            I => \N__6854\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__6854\,
            I => \N__6851\
        );

    \I__1388\ : Span4Mux_v
    port map (
            O => \N__6851\,
            I => \N__6848\
        );

    \I__1387\ : Sp12to4
    port map (
            O => \N__6848\,
            I => \N__6845\
        );

    \I__1386\ : Span12Mux_h
    port map (
            O => \N__6845\,
            I => \N__6842\
        );

    \I__1385\ : Odrv12
    port map (
            O => \N__6842\,
            I => \A_c_14\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__6839\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5_cascade_\
        );

    \I__1383\ : InMux
    port map (
            O => \N__6836\,
            I => \N__6833\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__6833\,
            I => \N__6830\
        );

    \I__1381\ : Sp12to4
    port map (
            O => \N__6830\,
            I => \N__6827\
        );

    \I__1380\ : Span12Mux_v
    port map (
            O => \N__6827\,
            I => \N__6824\
        );

    \I__1379\ : Span12Mux_h
    port map (
            O => \N__6824\,
            I => \N__6821\
        );

    \I__1378\ : Odrv12
    port map (
            O => \N__6821\,
            I => \A_c_7\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6818\,
            I => \N__6815\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__6815\,
            I => \N__6812\
        );

    \I__1375\ : Odrv12
    port map (
            O => \N__6812\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1374\ : InMux
    port map (
            O => \N__6809\,
            I => \N__6806\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__6806\,
            I => \N__6803\
        );

    \I__1372\ : Span4Mux_v
    port map (
            O => \N__6803\,
            I => \N__6800\
        );

    \I__1371\ : Span4Mux_h
    port map (
            O => \N__6800\,
            I => \N__6797\
        );

    \I__1370\ : Sp12to4
    port map (
            O => \N__6797\,
            I => \N__6794\
        );

    \I__1369\ : Odrv12
    port map (
            O => \N__6794\,
            I => \A_c_15\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__6791\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6_cascade_\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6785\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__6785\,
            I => \N__6782\
        );

    \I__1365\ : Span4Mux_v
    port map (
            O => \N__6782\,
            I => \N__6779\
        );

    \I__1364\ : Span4Mux_v
    port map (
            O => \N__6779\,
            I => \N__6776\
        );

    \I__1363\ : Sp12to4
    port map (
            O => \N__6776\,
            I => \N__6773\
        );

    \I__1362\ : Span12Mux_h
    port map (
            O => \N__6773\,
            I => \N__6770\
        );

    \I__1361\ : Odrv12
    port map (
            O => \N__6770\,
            I => \A_c_8\
        );

    \I__1360\ : InMux
    port map (
            O => \N__6767\,
            I => \N__6764\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__6764\,
            I => \N__6761\
        );

    \I__1358\ : Span4Mux_v
    port map (
            O => \N__6761\,
            I => \N__6758\
        );

    \I__1357\ : Span4Mux_v
    port map (
            O => \N__6758\,
            I => \N__6755\
        );

    \I__1356\ : Sp12to4
    port map (
            O => \N__6755\,
            I => \N__6752\
        );

    \I__1355\ : Span12Mux_h
    port map (
            O => \N__6752\,
            I => \N__6749\
        );

    \I__1354\ : Odrv12
    port map (
            O => \N__6749\,
            I => \A_c_9\
        );

    \I__1353\ : InMux
    port map (
            O => \N__6746\,
            I => \N__6743\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__6743\,
            I => \N__6740\
        );

    \I__1351\ : Span4Mux_v
    port map (
            O => \N__6740\,
            I => \N__6737\
        );

    \I__1350\ : Sp12to4
    port map (
            O => \N__6737\,
            I => \N__6734\
        );

    \I__1349\ : Span12Mux_v
    port map (
            O => \N__6734\,
            I => \N__6731\
        );

    \I__1348\ : Span12Mux_h
    port map (
            O => \N__6731\,
            I => \N__6728\
        );

    \I__1347\ : Odrv12
    port map (
            O => \N__6728\,
            I => \A_c_2\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__6725\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0_cascade_\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__6722\,
            I => \U712_CHIP_RAM.N_315_cascade_\
        );

    \I__1344\ : IoInMux
    port map (
            O => \N__6719\,
            I => \N__6716\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__6716\,
            I => \N__6713\
        );

    \I__1342\ : Span4Mux_s0_v
    port map (
            O => \N__6713\,
            I => \N__6710\
        );

    \I__1341\ : Sp12to4
    port map (
            O => \N__6710\,
            I => \N__6707\
        );

    \I__1340\ : Span12Mux_h
    port map (
            O => \N__6707\,
            I => \N__6704\
        );

    \I__1339\ : Odrv12
    port map (
            O => \N__6704\,
            I => \CMA_c_0\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6701\,
            I => \N__6698\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6698\,
            I => \N__6695\
        );

    \I__1336\ : Span4Mux_v
    port map (
            O => \N__6695\,
            I => \N__6692\
        );

    \I__1335\ : Sp12to4
    port map (
            O => \N__6692\,
            I => \N__6689\
        );

    \I__1334\ : Span12Mux_h
    port map (
            O => \N__6689\,
            I => \N__6686\
        );

    \I__1333\ : Span12Mux_v
    port map (
            O => \N__6686\,
            I => \N__6683\
        );

    \I__1332\ : Odrv12
    port map (
            O => \N__6683\,
            I => \A_c_3\
        );

    \I__1331\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6677\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__6677\,
            I => \N__6674\
        );

    \I__1329\ : Span4Mux_v
    port map (
            O => \N__6674\,
            I => \N__6671\
        );

    \I__1328\ : Span4Mux_h
    port map (
            O => \N__6671\,
            I => \N__6668\
        );

    \I__1327\ : Sp12to4
    port map (
            O => \N__6668\,
            I => \N__6665\
        );

    \I__1326\ : Odrv12
    port map (
            O => \N__6665\,
            I => \A_c_10\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__6662\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__6659\,
            I => \N__6656\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6656\,
            I => \N__6653\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6653\,
            I => \N__6650\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__6650\,
            I => \U712_CHIP_RAM.N_316\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__6647\,
            I => \N__6641\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6646\,
            I => \N__6635\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6645\,
            I => \N__6632\
        );

    \I__1317\ : InMux
    port map (
            O => \N__6644\,
            I => \N__6629\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6641\,
            I => \N__6626\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6619\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6639\,
            I => \N__6619\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6638\,
            I => \N__6619\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6635\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__6632\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__6629\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6626\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__6619\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1307\ : InMux
    port map (
            O => \N__6608\,
            I => \N__6600\
        );

    \I__1306\ : InMux
    port map (
            O => \N__6607\,
            I => \N__6597\
        );

    \I__1305\ : InMux
    port map (
            O => \N__6606\,
            I => \N__6590\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6605\,
            I => \N__6590\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6604\,
            I => \N__6590\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6603\,
            I => \N__6587\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__6600\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6597\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6590\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6587\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6578\,
            I => \N__6571\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6568\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6561\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6575\,
            I => \N__6561\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6574\,
            I => \N__6561\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__6571\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__6568\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__6561\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6548\
        );

    \I__1288\ : InMux
    port map (
            O => \N__6553\,
            I => \N__6543\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6552\,
            I => \N__6543\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6551\,
            I => \N__6540\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__6548\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__6543\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6540\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6533\,
            I => \N__6527\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6532\,
            I => \N__6524\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__6531\,
            I => \N__6520\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6530\,
            I => \N__6516\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__6527\,
            I => \N__6511\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6524\,
            I => \N__6511\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6523\,
            I => \N__6504\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6520\,
            I => \N__6504\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6504\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__6516\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__6511\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__6504\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1270\ : IoInMux
    port map (
            O => \N__6497\,
            I => \N__6494\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__6494\,
            I => \N__6491\
        );

    \I__1268\ : Odrv12
    port map (
            O => \N__6491\,
            I => \CMA_c_2\
        );

    \I__1267\ : IoInMux
    port map (
            O => \N__6488\,
            I => \N__6485\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__6485\,
            I => \N__6482\
        );

    \I__1265\ : Span4Mux_s3_v
    port map (
            O => \N__6482\,
            I => \N__6479\
        );

    \I__1264\ : Odrv4
    port map (
            O => \N__6479\,
            I => \CMA_c_1\
        );

    \I__1263\ : IoInMux
    port map (
            O => \N__6476\,
            I => \N__6473\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__6473\,
            I => \N__6470\
        );

    \I__1261\ : Span4Mux_s3_v
    port map (
            O => \N__6470\,
            I => \N__6467\
        );

    \I__1260\ : Span4Mux_h
    port map (
            O => \N__6467\,
            I => \N__6464\
        );

    \I__1259\ : Span4Mux_h
    port map (
            O => \N__6464\,
            I => \N__6461\
        );

    \I__1258\ : Odrv4
    port map (
            O => \N__6461\,
            I => \CMA_c_10\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6458\,
            I => \N__6455\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__6455\,
            I => \N__6452\
        );

    \I__1255\ : Span4Mux_v
    port map (
            O => \N__6452\,
            I => \N__6449\
        );

    \I__1254\ : Span4Mux_h
    port map (
            O => \N__6449\,
            I => \N__6446\
        );

    \I__1253\ : Sp12to4
    port map (
            O => \N__6446\,
            I => \N__6443\
        );

    \I__1252\ : Odrv12
    port map (
            O => \N__6443\,
            I => \A_c_11\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__6440\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6437\,
            I => \N__6434\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__6434\,
            I => \N__6431\
        );

    \I__1248\ : Span4Mux_v
    port map (
            O => \N__6431\,
            I => \N__6428\
        );

    \I__1247\ : Sp12to4
    port map (
            O => \N__6428\,
            I => \N__6425\
        );

    \I__1246\ : Span12Mux_h
    port map (
            O => \N__6425\,
            I => \N__6422\
        );

    \I__1245\ : Span12Mux_v
    port map (
            O => \N__6422\,
            I => \N__6419\
        );

    \I__1244\ : Odrv12
    port map (
            O => \N__6419\,
            I => \A_c_4\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6416\,
            I => \N__6413\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__6413\,
            I => \U712_CHIP_RAM.N_317\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__6410\,
            I => \N__6407\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6407\,
            I => \N__6402\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6406\,
            I => \N__6399\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6405\,
            I => \N__6396\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6402\,
            I => \U712_REG_SM.N_292\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6399\,
            I => \U712_REG_SM.N_292\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6396\,
            I => \U712_REG_SM.N_292\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6389\,
            I => \N__6384\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6379\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6387\,
            I => \N__6379\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__6384\,
            I => \U712_REG_SM.N_298\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__6379\,
            I => \U712_REG_SM.N_298\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__6374\,
            I => \N__6368\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6373\,
            I => \N__6365\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6362\
        );

    \I__1226\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6357\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6357\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6365\,
            I => \U712_REG_SM.N_294\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6362\,
            I => \U712_REG_SM.N_294\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__6357\,
            I => \U712_REG_SM.N_294\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6350\,
            I => \N__6344\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6344\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6344\,
            I => \U712_REG_SM.N_309\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__6341\,
            I => \N__6338\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6338\,
            I => \N__6334\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6331\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__6334\,
            I => \U712_REG_SM.N_282\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6331\,
            I => \U712_REG_SM.N_282\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__6326\,
            I => \U712_REG_SM.N_282_cascade_\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__6323\,
            I => \N__6319\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6322\,
            I => \N__6316\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6319\,
            I => \N__6313\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6316\,
            I => \N__6310\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__6313\,
            I => \U712_REG_SM.N_306\
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__6310\,
            I => \U712_REG_SM.N_306\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__6305\,
            I => \N__6301\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6304\,
            I => \N__6295\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6295\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6300\,
            I => \N__6292\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__6295\,
            I => \N__6287\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6292\,
            I => \N__6287\
        );

    \I__1200\ : Span12Mux_v
    port map (
            O => \N__6287\,
            I => \N__6284\
        );

    \I__1199\ : Span12Mux_h
    port map (
            O => \N__6284\,
            I => \N__6281\
        );

    \I__1198\ : Span12Mux_v
    port map (
            O => \N__6281\,
            I => \N__6278\
        );

    \I__1197\ : Odrv12
    port map (
            O => \N__6278\,
            I => \SIZ_c_1\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6275\,
            I => \N__6272\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__6272\,
            I => \N__6269\
        );

    \I__1194\ : Odrv4
    port map (
            O => \N__6269\,
            I => \U712_BYTE_ENABLE.N_407\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6266\,
            I => \N__6258\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6265\,
            I => \N__6258\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6264\,
            I => \N__6253\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6263\,
            I => \N__6253\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__6258\,
            I => \N__6248\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6253\,
            I => \N__6248\
        );

    \I__1187\ : Span4Mux_v
    port map (
            O => \N__6248\,
            I => \N__6245\
        );

    \I__1186\ : Sp12to4
    port map (
            O => \N__6245\,
            I => \N__6242\
        );

    \I__1185\ : Span12Mux_h
    port map (
            O => \N__6242\,
            I => \N__6239\
        );

    \I__1184\ : Span12Mux_v
    port map (
            O => \N__6239\,
            I => \N__6236\
        );

    \I__1183\ : Odrv12
    port map (
            O => \N__6236\,
            I => \A_c_1\
        );

    \I__1182\ : InMux
    port map (
            O => \N__6233\,
            I => \N__6225\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6232\,
            I => \N__6225\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6231\,
            I => \N__6222\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6230\,
            I => \N__6219\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6225\,
            I => \N__6214\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6222\,
            I => \N__6214\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__6219\,
            I => \N__6211\
        );

    \I__1175\ : Span4Mux_v
    port map (
            O => \N__6214\,
            I => \N__6208\
        );

    \I__1174\ : Span4Mux_v
    port map (
            O => \N__6211\,
            I => \N__6205\
        );

    \I__1173\ : Span4Mux_v
    port map (
            O => \N__6208\,
            I => \N__6198\
        );

    \I__1172\ : Span4Mux_v
    port map (
            O => \N__6205\,
            I => \N__6198\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6193\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6193\
        );

    \I__1169\ : Span4Mux_h
    port map (
            O => \N__6198\,
            I => \N__6190\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6193\,
            I => \N__6187\
        );

    \I__1167\ : Sp12to4
    port map (
            O => \N__6190\,
            I => \N__6182\
        );

    \I__1166\ : Span12Mux_v
    port map (
            O => \N__6187\,
            I => \N__6182\
        );

    \I__1165\ : Odrv12
    port map (
            O => \N__6182\,
            I => \A_c_0\
        );

    \I__1164\ : InMux
    port map (
            O => \N__6179\,
            I => \N__6176\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6176\,
            I => \U712_BYTE_ENABLE.N_409\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6173\,
            I => \N__6170\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__6170\,
            I => \N__6166\
        );

    \I__1160\ : IoInMux
    port map (
            O => \N__6169\,
            I => \N__6163\
        );

    \I__1159\ : Span4Mux_v
    port map (
            O => \N__6166\,
            I => \N__6160\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6163\,
            I => \N__6157\
        );

    \I__1157\ : Sp12to4
    port map (
            O => \N__6160\,
            I => \N__6154\
        );

    \I__1156\ : Span4Mux_s3_h
    port map (
            O => \N__6157\,
            I => \N__6151\
        );

    \I__1155\ : Span12Mux_h
    port map (
            O => \N__6154\,
            I => \N__6146\
        );

    \I__1154\ : Sp12to4
    port map (
            O => \N__6151\,
            I => \N__6146\
        );

    \I__1153\ : Span12Mux_v
    port map (
            O => \N__6146\,
            I => \N__6143\
        );

    \I__1152\ : Odrv12
    port map (
            O => \N__6143\,
            I => \C1_c\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6137\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6137\,
            I => \N__6134\
        );

    \I__1149\ : Span12Mux_h
    port map (
            O => \N__6134\,
            I => \N__6131\
        );

    \I__1148\ : Span12Mux_v
    port map (
            O => \N__6131\,
            I => \N__6128\
        );

    \I__1147\ : Odrv12
    port map (
            O => \N__6128\,
            I => \C3_c\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6125\,
            I => \N__6121\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6124\,
            I => \N__6118\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6121\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6118\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__6113\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0_cascade_\
        );

    \I__1141\ : IoInMux
    port map (
            O => \N__6110\,
            I => \N__6107\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__6107\,
            I => \N__6104\
        );

    \I__1139\ : Span4Mux_s3_h
    port map (
            O => \N__6104\,
            I => \N__6101\
        );

    \I__1138\ : Span4Mux_v
    port map (
            O => \N__6101\,
            I => \N__6098\
        );

    \I__1137\ : Sp12to4
    port map (
            O => \N__6098\,
            I => \N__6095\
        );

    \I__1136\ : Span12Mux_h
    port map (
            O => \N__6095\,
            I => \N__6092\
        );

    \I__1135\ : Odrv12
    port map (
            O => \N__6092\,
            I => \N_192_i\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6089\,
            I => \N__6086\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6086\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0\
        );

    \I__1132\ : IoInMux
    port map (
            O => \N__6083\,
            I => \N__6080\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6080\,
            I => \N__6077\
        );

    \I__1130\ : Span12Mux_s6_h
    port map (
            O => \N__6077\,
            I => \N__6074\
        );

    \I__1129\ : Span12Mux_h
    port map (
            O => \N__6074\,
            I => \N__6071\
        );

    \I__1128\ : Span12Mux_v
    port map (
            O => \N__6071\,
            I => \N__6068\
        );

    \I__1127\ : Odrv12
    port map (
            O => \N__6068\,
            I => \N_194_i\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6065\,
            I => \N__6062\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6062\,
            I => \N__6059\
        );

    \I__1124\ : Span4Mux_v
    port map (
            O => \N__6059\,
            I => \N__6055\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6058\,
            I => \N__6052\
        );

    \I__1122\ : Sp12to4
    port map (
            O => \N__6055\,
            I => \N__6047\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6052\,
            I => \N__6047\
        );

    \I__1120\ : Span12Mux_h
    port map (
            O => \N__6047\,
            I => \N__6044\
        );

    \I__1119\ : Span12Mux_v
    port map (
            O => \N__6044\,
            I => \N__6041\
        );

    \I__1118\ : Odrv12
    port map (
            O => \N__6041\,
            I => \SIZ_c_0\
        );

    \I__1117\ : IoInMux
    port map (
            O => \N__6038\,
            I => \N__6035\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6035\,
            I => \N__6032\
        );

    \I__1115\ : Span4Mux_s3_v
    port map (
            O => \N__6032\,
            I => \N__6029\
        );

    \I__1114\ : Span4Mux_v
    port map (
            O => \N__6029\,
            I => \N__6026\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__6026\,
            I => \N__6021\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6025\,
            I => \N__6018\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6024\,
            I => \N__6015\
        );

    \I__1110\ : Span4Mux_h
    port map (
            O => \N__6021\,
            I => \N__6011\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6018\,
            I => \N__6006\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6015\,
            I => \N__6006\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6014\,
            I => \N__6003\
        );

    \I__1106\ : Odrv4
    port map (
            O => \N__6011\,
            I => \DBENn_c\
        );

    \I__1105\ : Odrv4
    port map (
            O => \N__6006\,
            I => \DBENn_c\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6003\,
            I => \DBENn_c\
        );

    \I__1103\ : IoInMux
    port map (
            O => \N__5996\,
            I => \N__5993\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5993\,
            I => \N__5990\
        );

    \I__1101\ : Span4Mux_s2_v
    port map (
            O => \N__5990\,
            I => \N__5987\
        );

    \I__1100\ : Span4Mux_h
    port map (
            O => \N__5987\,
            I => \N__5984\
        );

    \I__1099\ : Span4Mux_h
    port map (
            O => \N__5984\,
            I => \N__5979\
        );

    \I__1098\ : InMux
    port map (
            O => \N__5983\,
            I => \N__5974\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5982\,
            I => \N__5974\
        );

    \I__1096\ : Sp12to4
    port map (
            O => \N__5979\,
            I => \N__5969\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5974\,
            I => \N__5966\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5973\,
            I => \N__5963\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5960\
        );

    \I__1092\ : Span12Mux_s9_v
    port map (
            O => \N__5969\,
            I => \N__5948\
        );

    \I__1091\ : Sp12to4
    port map (
            O => \N__5966\,
            I => \N__5948\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__5963\,
            I => \N__5948\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5960\,
            I => \N__5948\
        );

    \I__1088\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5941\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5941\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5957\,
            I => \N__5941\
        );

    \I__1085\ : Odrv12
    port map (
            O => \N__5948\,
            I => \RAMENn_c\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__5941\,
            I => \RAMENn_c\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__5936\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_cascade_\
        );

    \I__1082\ : IoInMux
    port map (
            O => \N__5933\,
            I => \N__5930\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__5930\,
            I => \N__5927\
        );

    \I__1080\ : Span12Mux_s6_h
    port map (
            O => \N__5927\,
            I => \N__5924\
        );

    \I__1079\ : Span12Mux_h
    port map (
            O => \N__5924\,
            I => \N__5921\
        );

    \I__1078\ : Span12Mux_v
    port map (
            O => \N__5921\,
            I => \N__5918\
        );

    \I__1077\ : Odrv12
    port map (
            O => \N__5918\,
            I => \N_196_i\
        );

    \I__1076\ : InMux
    port map (
            O => \N__5915\,
            I => \N__5907\
        );

    \I__1075\ : InMux
    port map (
            O => \N__5914\,
            I => \N__5907\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5913\,
            I => \N__5902\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5912\,
            I => \N__5902\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5907\,
            I => \U712_BYTE_ENABLE.N_404\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__5902\,
            I => \U712_BYTE_ENABLE.N_404\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5897\,
            I => \N__5894\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5894\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__5891\,
            I => \U712_BYTE_ENABLE.N_411_cascade_\
        );

    \I__1067\ : IoInMux
    port map (
            O => \N__5888\,
            I => \N__5885\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5885\,
            I => \N__5882\
        );

    \I__1065\ : IoSpan4Mux
    port map (
            O => \N__5882\,
            I => \N__5879\
        );

    \I__1064\ : Sp12to4
    port map (
            O => \N__5879\,
            I => \N__5876\
        );

    \I__1063\ : Span12Mux_s7_v
    port map (
            O => \N__5876\,
            I => \N__5873\
        );

    \I__1062\ : Odrv12
    port map (
            O => \N__5873\,
            I => \N_198_i\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5867\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__5867\,
            I => \U712_BYTE_ENABLE.N_405\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__5864\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_cascade_\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5858\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__5858\,
            I => \U712_CHIP_RAM.DBENn_7_0_a2_0\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__5855\,
            I => \N__5852\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5847\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5851\,
            I => \N__5844\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5850\,
            I => \N__5841\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5847\,
            I => \N__5838\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__5844\,
            I => \N__5835\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__5841\,
            I => \U712_CHIP_RAM.N_347\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__5838\,
            I => \U712_CHIP_RAM.N_347\
        );

    \I__1048\ : Odrv4
    port map (
            O => \N__5835\,
            I => \U712_CHIP_RAM.N_347\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5828\,
            I => \N__5825\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__5825\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_3_1\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__5822\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_2_1_cascade_\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5819\,
            I => \N__5814\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5811\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5808\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5814\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER50\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5811\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER50\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__5808\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER50\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5795\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5784\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__5799\,
            I => \N__5778\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5775\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5795\,
            I => \N__5772\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5794\,
            I => \N__5765\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5765\
        );

    \I__1031\ : InMux
    port map (
            O => \N__5792\,
            I => \N__5765\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5791\,
            I => \N__5758\
        );

    \I__1029\ : InMux
    port map (
            O => \N__5790\,
            I => \N__5758\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5789\,
            I => \N__5758\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5788\,
            I => \N__5753\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5787\,
            I => \N__5753\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5784\,
            I => \N__5750\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__5783\,
            I => \N__5747\
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__5782\,
            I => \N__5743\
        );

    \I__1022\ : CascadeMux
    port map (
            O => \N__5781\,
            I => \N__5738\
        );

    \I__1021\ : InMux
    port map (
            O => \N__5778\,
            I => \N__5728\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5775\,
            I => \N__5723\
        );

    \I__1019\ : Span4Mux_v
    port map (
            O => \N__5772\,
            I => \N__5723\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5765\,
            I => \N__5720\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5758\,
            I => \N__5713\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5753\,
            I => \N__5713\
        );

    \I__1015\ : Span4Mux_h
    port map (
            O => \N__5750\,
            I => \N__5713\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5747\,
            I => \N__5706\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5746\,
            I => \N__5706\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5743\,
            I => \N__5706\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5742\,
            I => \N__5701\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5741\,
            I => \N__5701\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5738\,
            I => \N__5696\
        );

    \I__1008\ : InMux
    port map (
            O => \N__5737\,
            I => \N__5696\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5736\,
            I => \N__5693\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5735\,
            I => \N__5686\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5686\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5686\
        );

    \I__1003\ : InMux
    port map (
            O => \N__5732\,
            I => \N__5681\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5681\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__5728\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1000\ : Odrv4
    port map (
            O => \N__5723\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__999\ : Odrv12
    port map (
            O => \N__5720\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__998\ : Odrv4
    port map (
            O => \N__5713\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5706\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5701\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5696\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5693\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5686\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5681\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__991\ : InMux
    port map (
            O => \N__5660\,
            I => \N__5653\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__5659\,
            I => \N__5650\
        );

    \I__989\ : CascadeMux
    port map (
            O => \N__5658\,
            I => \N__5647\
        );

    \I__988\ : CascadeMux
    port map (
            O => \N__5657\,
            I => \N__5643\
        );

    \I__987\ : InMux
    port map (
            O => \N__5656\,
            I => \N__5639\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5653\,
            I => \N__5634\
        );

    \I__985\ : InMux
    port map (
            O => \N__5650\,
            I => \N__5629\
        );

    \I__984\ : InMux
    port map (
            O => \N__5647\,
            I => \N__5629\
        );

    \I__983\ : InMux
    port map (
            O => \N__5646\,
            I => \N__5626\
        );

    \I__982\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5623\
        );

    \I__981\ : InMux
    port map (
            O => \N__5642\,
            I => \N__5620\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__5639\,
            I => \N__5617\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__5638\,
            I => \N__5608\
        );

    \I__978\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5602\
        );

    \I__977\ : Span4Mux_v
    port map (
            O => \N__5634\,
            I => \N__5597\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5629\,
            I => \N__5597\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__5626\,
            I => \N__5592\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__5623\,
            I => \N__5592\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__5620\,
            I => \N__5587\
        );

    \I__972\ : Span4Mux_v
    port map (
            O => \N__5617\,
            I => \N__5587\
        );

    \I__971\ : InMux
    port map (
            O => \N__5616\,
            I => \N__5582\
        );

    \I__970\ : InMux
    port map (
            O => \N__5615\,
            I => \N__5582\
        );

    \I__969\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5579\
        );

    \I__968\ : InMux
    port map (
            O => \N__5613\,
            I => \N__5572\
        );

    \I__967\ : InMux
    port map (
            O => \N__5612\,
            I => \N__5572\
        );

    \I__966\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5572\
        );

    \I__965\ : InMux
    port map (
            O => \N__5608\,
            I => \N__5567\
        );

    \I__964\ : InMux
    port map (
            O => \N__5607\,
            I => \N__5567\
        );

    \I__963\ : InMux
    port map (
            O => \N__5606\,
            I => \N__5562\
        );

    \I__962\ : InMux
    port map (
            O => \N__5605\,
            I => \N__5562\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__5602\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__960\ : Odrv4
    port map (
            O => \N__5597\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__959\ : Odrv4
    port map (
            O => \N__5592\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__958\ : Odrv4
    port map (
            O => \N__5587\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__5582\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__5579\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5572\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5567\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5562\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__952\ : InMux
    port map (
            O => \N__5543\,
            I => \N__5536\
        );

    \I__951\ : InMux
    port map (
            O => \N__5542\,
            I => \N__5536\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__5541\,
            I => \N__5532\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5536\,
            I => \N__5528\
        );

    \I__948\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5525\
        );

    \I__947\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5520\
        );

    \I__946\ : InMux
    port map (
            O => \N__5531\,
            I => \N__5520\
        );

    \I__945\ : Odrv4
    port map (
            O => \N__5528\,
            I => \U712_CHIP_RAM.N_273\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5525\,
            I => \U712_CHIP_RAM.N_273\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__5520\,
            I => \U712_CHIP_RAM.N_273\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__5513\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_1_0_cascade_\
        );

    \I__941\ : InMux
    port map (
            O => \N__5510\,
            I => \N__5506\
        );

    \I__940\ : InMux
    port map (
            O => \N__5509\,
            I => \N__5503\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5506\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5503\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__5498\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_0_cascade_\
        );

    \I__936\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5487\
        );

    \I__935\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5487\
        );

    \I__934\ : InMux
    port map (
            O => \N__5493\,
            I => \N__5482\
        );

    \I__933\ : InMux
    port map (
            O => \N__5492\,
            I => \N__5482\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__5487\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5482\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__5477\,
            I => \U712_CHIP_RAM.REFRESH_RST_cascade_\
        );

    \I__929\ : InMux
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5471\,
            I => \U712_CHIP_RAM.N_289\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__5468\,
            I => \U712_CHIP_RAM.N_425_cascade_\
        );

    \I__926\ : InMux
    port map (
            O => \N__5465\,
            I => \N__5461\
        );

    \I__925\ : InMux
    port map (
            O => \N__5464\,
            I => \N__5458\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5461\,
            I => \U712_CHIP_RAM.N_424\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5458\,
            I => \U712_CHIP_RAM.N_424\
        );

    \I__922\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5450\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__5450\,
            I => \U712_CHIP_RAM.N_302\
        );

    \I__920\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5443\
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__5446\,
            I => \N__5439\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5443\,
            I => \N__5435\
        );

    \I__917\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5428\
        );

    \I__916\ : InMux
    port map (
            O => \N__5439\,
            I => \N__5428\
        );

    \I__915\ : InMux
    port map (
            O => \N__5438\,
            I => \N__5428\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__5435\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5428\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__5423\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_START_2_0_a2_1_cascade_\
        );

    \I__911\ : InMux
    port map (
            O => \N__5420\,
            I => \N__5416\
        );

    \I__910\ : InMux
    port map (
            O => \N__5419\,
            I => \N__5413\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5416\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__5413\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__907\ : InMux
    port map (
            O => \N__5408\,
            I => \N__5403\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__5407\,
            I => \N__5398\
        );

    \I__905\ : InMux
    port map (
            O => \N__5406\,
            I => \N__5392\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5403\,
            I => \N__5388\
        );

    \I__903\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5385\
        );

    \I__902\ : InMux
    port map (
            O => \N__5401\,
            I => \N__5376\
        );

    \I__901\ : InMux
    port map (
            O => \N__5398\,
            I => \N__5376\
        );

    \I__900\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5376\
        );

    \I__899\ : InMux
    port map (
            O => \N__5396\,
            I => \N__5376\
        );

    \I__898\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5373\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5392\,
            I => \N__5370\
        );

    \I__896\ : InMux
    port map (
            O => \N__5391\,
            I => \N__5367\
        );

    \I__895\ : Odrv4
    port map (
            O => \N__5388\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__5385\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5376\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5373\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__891\ : Odrv12
    port map (
            O => \N__5370\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5367\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__5354\,
            I => \N__5350\
        );

    \I__888\ : CascadeMux
    port map (
            O => \N__5353\,
            I => \N__5346\
        );

    \I__887\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5343\
        );

    \I__886\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5340\
        );

    \I__885\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5335\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5343\,
            I => \N__5331\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__5340\,
            I => \N__5328\
        );

    \I__882\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5320\
        );

    \I__881\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5317\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5335\,
            I => \N__5314\
        );

    \I__879\ : InMux
    port map (
            O => \N__5334\,
            I => \N__5311\
        );

    \I__878\ : Span4Mux_v
    port map (
            O => \N__5331\,
            I => \N__5306\
        );

    \I__877\ : Span4Mux_v
    port map (
            O => \N__5328\,
            I => \N__5306\
        );

    \I__876\ : InMux
    port map (
            O => \N__5327\,
            I => \N__5303\
        );

    \I__875\ : InMux
    port map (
            O => \N__5326\,
            I => \N__5300\
        );

    \I__874\ : InMux
    port map (
            O => \N__5325\,
            I => \N__5297\
        );

    \I__873\ : InMux
    port map (
            O => \N__5324\,
            I => \N__5292\
        );

    \I__872\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5292\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5320\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5317\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__869\ : Odrv12
    port map (
            O => \N__5314\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5311\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__867\ : Odrv4
    port map (
            O => \N__5306\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5303\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5300\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5297\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5292\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__862\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5270\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5270\,
            I => \U712_CHIP_RAM.N_438\
        );

    \I__860\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5264\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5264\,
            I => \N__5254\
        );

    \I__858\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5251\
        );

    \I__857\ : InMux
    port map (
            O => \N__5262\,
            I => \N__5248\
        );

    \I__856\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5243\
        );

    \I__855\ : InMux
    port map (
            O => \N__5260\,
            I => \N__5240\
        );

    \I__854\ : InMux
    port map (
            O => \N__5259\,
            I => \N__5233\
        );

    \I__853\ : InMux
    port map (
            O => \N__5258\,
            I => \N__5233\
        );

    \I__852\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5233\
        );

    \I__851\ : Span4Mux_h
    port map (
            O => \N__5254\,
            I => \N__5228\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5251\,
            I => \N__5228\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5248\,
            I => \N__5225\
        );

    \I__848\ : InMux
    port map (
            O => \N__5247\,
            I => \N__5220\
        );

    \I__847\ : InMux
    port map (
            O => \N__5246\,
            I => \N__5220\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5243\,
            I => \U712_CHIP_RAM.N_284\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5240\,
            I => \U712_CHIP_RAM.N_284\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5233\,
            I => \U712_CHIP_RAM.N_284\
        );

    \I__843\ : Odrv4
    port map (
            O => \N__5228\,
            I => \U712_CHIP_RAM.N_284\
        );

    \I__842\ : Odrv4
    port map (
            O => \N__5225\,
            I => \U712_CHIP_RAM.N_284\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5220\,
            I => \U712_CHIP_RAM.N_284\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__5207\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_1_cascade_\
        );

    \I__839\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5197\
        );

    \I__838\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5197\
        );

    \I__837\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5193\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__5197\,
            I => \N__5190\
        );

    \I__835\ : InMux
    port map (
            O => \N__5196\,
            I => \N__5187\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5193\,
            I => \N__5182\
        );

    \I__833\ : Span4Mux_v
    port map (
            O => \N__5190\,
            I => \N__5182\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5187\,
            I => \U712_CHIP_RAM.N_272\
        );

    \I__831\ : Odrv4
    port map (
            O => \N__5182\,
            I => \U712_CHIP_RAM.N_272\
        );

    \I__830\ : InMux
    port map (
            O => \N__5177\,
            I => \N__5174\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__5174\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0\
        );

    \I__828\ : InMux
    port map (
            O => \N__5171\,
            I => \N__5168\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5168\,
            I => \U712_CHIP_RAM.N_310\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__5165\,
            I => \U712_CHIP_RAM.N_310_cascade_\
        );

    \I__825\ : InMux
    port map (
            O => \N__5162\,
            I => \N__5155\
        );

    \I__824\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5155\
        );

    \I__823\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5152\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5155\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5152\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__5147\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_3_0_a2_i_0_cascade_\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__5144\,
            I => \U712_CHIP_RAM.N_179_cascade_\
        );

    \I__818\ : IoInMux
    port map (
            O => \N__5141\,
            I => \N__5138\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5138\,
            I => \N__5135\
        );

    \I__816\ : IoSpan4Mux
    port map (
            O => \N__5135\,
            I => \N__5132\
        );

    \I__815\ : Span4Mux_s3_h
    port map (
            O => \N__5132\,
            I => \N__5129\
        );

    \I__814\ : Span4Mux_h
    port map (
            O => \N__5129\,
            I => \N__5126\
        );

    \I__813\ : Sp12to4
    port map (
            O => \N__5126\,
            I => \N__5123\
        );

    \I__812\ : Span12Mux_h
    port map (
            O => \N__5123\,
            I => \N__5119\
        );

    \I__811\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5116\
        );

    \I__810\ : Odrv12
    port map (
            O => \N__5119\,
            I => \CLK_EN_c\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__5116\,
            I => \CLK_EN_c\
        );

    \I__808\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5106\
        );

    \I__807\ : InMux
    port map (
            O => \N__5110\,
            I => \N__5101\
        );

    \I__806\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5101\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5106\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5101\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__803\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5092\
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__5095\,
            I => \N__5086\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5092\,
            I => \N__5082\
        );

    \I__800\ : CascadeMux
    port map (
            O => \N__5091\,
            I => \N__5078\
        );

    \I__799\ : InMux
    port map (
            O => \N__5090\,
            I => \N__5071\
        );

    \I__798\ : InMux
    port map (
            O => \N__5089\,
            I => \N__5068\
        );

    \I__797\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5065\
        );

    \I__796\ : InMux
    port map (
            O => \N__5085\,
            I => \N__5062\
        );

    \I__795\ : Span4Mux_h
    port map (
            O => \N__5082\,
            I => \N__5059\
        );

    \I__794\ : InMux
    port map (
            O => \N__5081\,
            I => \N__5056\
        );

    \I__793\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5053\
        );

    \I__792\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5048\
        );

    \I__791\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5048\
        );

    \I__790\ : InMux
    port map (
            O => \N__5075\,
            I => \N__5043\
        );

    \I__789\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5043\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5071\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5068\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5065\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5062\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__5059\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5056\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5053\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5048\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5043\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__5024\,
            I => \U712_CHIP_RAM.N_438_cascade_\
        );

    \I__778\ : CascadeMux
    port map (
            O => \N__5021\,
            I => \U712_REG_SM.N_292_cascade_\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__5018\,
            I => \N__5015\
        );

    \I__776\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5011\
        );

    \I__775\ : InMux
    port map (
            O => \N__5014\,
            I => \N__5008\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5011\,
            I => \U712_REG_SM.N_507\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__5008\,
            I => \U712_REG_SM.N_507\
        );

    \I__772\ : InMux
    port map (
            O => \N__5003\,
            I => \N__5000\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5000\,
            I => \N__4994\
        );

    \I__770\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4991\
        );

    \I__769\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4988\
        );

    \I__768\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4985\
        );

    \I__767\ : Span4Mux_v
    port map (
            O => \N__4994\,
            I => \N__4978\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4991\,
            I => \N__4978\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4988\,
            I => \N__4978\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4985\,
            I => \N__4975\
        );

    \I__763\ : Span4Mux_v
    port map (
            O => \N__4978\,
            I => \N__4972\
        );

    \I__762\ : Span4Mux_v
    port map (
            O => \N__4975\,
            I => \N__4969\
        );

    \I__761\ : Sp12to4
    port map (
            O => \N__4972\,
            I => \N__4964\
        );

    \I__760\ : Sp12to4
    port map (
            O => \N__4969\,
            I => \N__4964\
        );

    \I__759\ : Span12Mux_h
    port map (
            O => \N__4964\,
            I => \N__4961\
        );

    \I__758\ : Span12Mux_v
    port map (
            O => \N__4961\,
            I => \N__4958\
        );

    \I__757\ : Odrv12
    port map (
            O => \N__4958\,
            I => \RnW_c\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__755\ : InMux
    port map (
            O => \N__4952\,
            I => \N__4949\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__4949\,
            I => \U712_REG_SM.N_104\
        );

    \I__753\ : InMux
    port map (
            O => \N__4946\,
            I => \N__4941\
        );

    \I__752\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4938\
        );

    \I__751\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4935\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__4941\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4938\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4935\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__747\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4925\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4925\,
            I => \U712_REG_SM.N_372\
        );

    \I__745\ : CascadeMux
    port map (
            O => \N__4922\,
            I => \N__4917\
        );

    \I__744\ : InMux
    port map (
            O => \N__4921\,
            I => \N__4914\
        );

    \I__743\ : InMux
    port map (
            O => \N__4920\,
            I => \N__4911\
        );

    \I__742\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4908\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4914\,
            I => \N__4903\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4911\,
            I => \N__4903\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4908\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__738\ : Odrv4
    port map (
            O => \N__4903\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__737\ : IoInMux
    port map (
            O => \N__4898\,
            I => \N__4895\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__4895\,
            I => \N__4891\
        );

    \I__735\ : IoInMux
    port map (
            O => \N__4894\,
            I => \N__4888\
        );

    \I__734\ : IoSpan4Mux
    port map (
            O => \N__4891\,
            I => \N__4885\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4888\,
            I => \N__4882\
        );

    \I__732\ : Span4Mux_s2_v
    port map (
            O => \N__4885\,
            I => \N__4879\
        );

    \I__731\ : IoSpan4Mux
    port map (
            O => \N__4882\,
            I => \N__4876\
        );

    \I__730\ : Sp12to4
    port map (
            O => \N__4879\,
            I => \N__4873\
        );

    \I__729\ : Span4Mux_s2_v
    port map (
            O => \N__4876\,
            I => \N__4870\
        );

    \I__728\ : Span12Mux_v
    port map (
            O => \N__4873\,
            I => \N__4867\
        );

    \I__727\ : Sp12to4
    port map (
            O => \N__4870\,
            I => \N__4864\
        );

    \I__726\ : Span12Mux_h
    port map (
            O => \N__4867\,
            I => \N__4859\
        );

    \I__725\ : Span12Mux_v
    port map (
            O => \N__4864\,
            I => \N__4859\
        );

    \I__724\ : Odrv12
    port map (
            O => \N__4859\,
            I => \ASn_c\
        );

    \I__723\ : CEMux
    port map (
            O => \N__4856\,
            I => \N__4853\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4853\,
            I => \U712_REG_SM.N_186_0\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__4850\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_cascade_\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__4847\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_0_a2_2_cascade_\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__4844\,
            I => \N__4841\
        );

    \I__718\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4838\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4838\,
            I => \U712_CHIP_RAM.N_393\
        );

    \I__716\ : InMux
    port map (
            O => \N__4835\,
            I => \N__4829\
        );

    \I__715\ : InMux
    port map (
            O => \N__4834\,
            I => \N__4824\
        );

    \I__714\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4824\
        );

    \I__713\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4821\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4829\,
            I => \N__4818\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__4824\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4821\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__709\ : Odrv4
    port map (
            O => \N__4818\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__708\ : CascadeMux
    port map (
            O => \N__4811\,
            I => \U712_REG_SM.N_301_cascade_\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__4808\,
            I => \N__4804\
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__4807\,
            I => \N__4801\
        );

    \I__705\ : InMux
    port map (
            O => \N__4804\,
            I => \N__4797\
        );

    \I__704\ : InMux
    port map (
            O => \N__4801\,
            I => \N__4794\
        );

    \I__703\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4791\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__4797\,
            I => \U712_REG_SM.N_288\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__4794\,
            I => \U712_REG_SM.N_288\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4791\,
            I => \U712_REG_SM.N_288\
        );

    \I__699\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4779\
        );

    \I__698\ : InMux
    port map (
            O => \N__4783\,
            I => \N__4776\
        );

    \I__697\ : InMux
    port map (
            O => \N__4782\,
            I => \N__4773\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__4779\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4776\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4773\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__693\ : InMux
    port map (
            O => \N__4766\,
            I => \N__4760\
        );

    \I__692\ : InMux
    port map (
            O => \N__4765\,
            I => \N__4760\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__4760\,
            I => \U712_REG_SM.N_301\
        );

    \I__690\ : InMux
    port map (
            O => \N__4757\,
            I => \N__4748\
        );

    \I__689\ : InMux
    port map (
            O => \N__4756\,
            I => \N__4748\
        );

    \I__688\ : InMux
    port map (
            O => \N__4755\,
            I => \N__4748\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__4748\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__686\ : InMux
    port map (
            O => \N__4745\,
            I => \N__4742\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4742\,
            I => \N__4739\
        );

    \I__684\ : Span4Mux_v
    port map (
            O => \N__4739\,
            I => \N__4733\
        );

    \I__683\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4726\
        );

    \I__682\ : InMux
    port map (
            O => \N__4737\,
            I => \N__4726\
        );

    \I__681\ : InMux
    port map (
            O => \N__4736\,
            I => \N__4726\
        );

    \I__680\ : Odrv4
    port map (
            O => \N__4733\,
            I => \REG_CYCLEm\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__4726\,
            I => \REG_CYCLEm\
        );

    \I__678\ : IoInMux
    port map (
            O => \N__4721\,
            I => \N__4718\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4718\,
            I => \N__4715\
        );

    \I__676\ : IoSpan4Mux
    port map (
            O => \N__4715\,
            I => \N__4712\
        );

    \I__675\ : IoSpan4Mux
    port map (
            O => \N__4712\,
            I => \N__4709\
        );

    \I__674\ : IoSpan4Mux
    port map (
            O => \N__4709\,
            I => \N__4706\
        );

    \I__673\ : Span4Mux_s3_v
    port map (
            O => \N__4706\,
            I => \N__4703\
        );

    \I__672\ : Sp12to4
    port map (
            O => \N__4703\,
            I => \N__4700\
        );

    \I__671\ : Span12Mux_v
    port map (
            O => \N__4700\,
            I => \N__4697\
        );

    \I__670\ : Odrv12
    port map (
            O => \N__4697\,
            I => \DRDENn_c\
        );

    \I__669\ : CascadeMux
    port map (
            O => \N__4694\,
            I => \N__4691\
        );

    \I__668\ : InMux
    port map (
            O => \N__4691\,
            I => \N__4687\
        );

    \I__667\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4684\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__4687\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4684\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__664\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4673\
        );

    \I__663\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4673\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__4673\,
            I => \U712_REG_SM.N_341\
        );

    \I__661\ : CascadeMux
    port map (
            O => \N__4670\,
            I => \U712_REG_SM.N_294_cascade_\
        );

    \I__660\ : InMux
    port map (
            O => \N__4667\,
            I => \N__4664\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__4664\,
            I => \N__4661\
        );

    \I__658\ : Odrv4
    port map (
            O => \N__4661\,
            I => \U712_REG_SM.N_373\
        );

    \I__657\ : InMux
    port map (
            O => \N__4658\,
            I => \N__4652\
        );

    \I__656\ : InMux
    port map (
            O => \N__4657\,
            I => \N__4652\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__4649\,
            I => \U712_CHIP_RAM.N_296_i\
        );

    \I__653\ : CascadeMux
    port map (
            O => \N__4646\,
            I => \U712_CHIP_RAM.SDRAM_CMD_e_1_2_cascade_\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__4643\,
            I => \N__4640\
        );

    \I__651\ : InMux
    port map (
            O => \N__4640\,
            I => \N__4637\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4637\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_0_3\
        );

    \I__649\ : CEMux
    port map (
            O => \N__4634\,
            I => \N__4631\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4631\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0\
        );

    \I__647\ : IoInMux
    port map (
            O => \N__4628\,
            I => \N__4625\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__645\ : Span4Mux_s2_v
    port map (
            O => \N__4622\,
            I => \N__4618\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__4621\,
            I => \N__4615\
        );

    \I__643\ : Sp12to4
    port map (
            O => \N__4618\,
            I => \N__4611\
        );

    \I__642\ : InMux
    port map (
            O => \N__4615\,
            I => \N__4608\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__4614\,
            I => \N__4605\
        );

    \I__640\ : Span12Mux_h
    port map (
            O => \N__4611\,
            I => \N__4602\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4608\,
            I => \N__4599\
        );

    \I__638\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4596\
        );

    \I__637\ : Odrv12
    port map (
            O => \N__4602\,
            I => \DBDIR_c\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__4599\,
            I => \DBDIR_c\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4596\,
            I => \DBDIR_c\
        );

    \I__634\ : IoInMux
    port map (
            O => \N__4589\,
            I => \N__4586\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4586\,
            I => \N__4583\
        );

    \I__632\ : IoSpan4Mux
    port map (
            O => \N__4583\,
            I => \N__4580\
        );

    \I__631\ : Span4Mux_s2_h
    port map (
            O => \N__4580\,
            I => \N__4577\
        );

    \I__630\ : Sp12to4
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__629\ : Span12Mux_s11_h
    port map (
            O => \N__4574\,
            I => \N__4571\
        );

    \I__628\ : Span12Mux_v
    port map (
            O => \N__4571\,
            I => \N__4568\
        );

    \I__627\ : Odrv12
    port map (
            O => \N__4568\,
            I => \N_188\
        );

    \I__626\ : InMux
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4562\,
            I => \N__4559\
        );

    \I__624\ : Span4Mux_v
    port map (
            O => \N__4559\,
            I => \N__4554\
        );

    \I__623\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4549\
        );

    \I__622\ : InMux
    port map (
            O => \N__4557\,
            I => \N__4549\
        );

    \I__621\ : Odrv4
    port map (
            O => \N__4554\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__4549\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__4544\,
            I => \U712_REG_SM.N_288_cascade_\
        );

    \I__618\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4538\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__4538\,
            I => \N__4534\
        );

    \I__616\ : InMux
    port map (
            O => \N__4537\,
            I => \N__4529\
        );

    \I__615\ : Span4Mux_v
    port map (
            O => \N__4534\,
            I => \N__4526\
        );

    \I__614\ : InMux
    port map (
            O => \N__4533\,
            I => \N__4521\
        );

    \I__613\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4521\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4529\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__611\ : Odrv4
    port map (
            O => \N__4526\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4521\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__4514\,
            I => \U712_CHIP_RAM.N_347_cascade_\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__4511\,
            I => \U712_CHIP_RAM.N_378_cascade_\
        );

    \I__607\ : InMux
    port map (
            O => \N__4508\,
            I => \N__4505\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__4505\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_tz\
        );

    \I__605\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4499\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_0_a2_0_a2_0\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__4496\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_0_cascade_\
        );

    \I__602\ : CascadeMux
    port map (
            O => \N__4493\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER50_cascade_\
        );

    \I__601\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4486\
        );

    \I__600\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4483\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4486\,
            I => \N__4478\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__4483\,
            I => \N__4478\
        );

    \I__597\ : Span12Mux_h
    port map (
            O => \N__4478\,
            I => \N__4475\
        );

    \I__596\ : Span12Mux_v
    port map (
            O => \N__4475\,
            I => \N__4472\
        );

    \I__595\ : Odrv12
    port map (
            O => \N__4472\,
            I => \AWEn_c\
        );

    \I__594\ : InMux
    port map (
            O => \N__4469\,
            I => \N__4466\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4466\,
            I => \U712_CHIP_RAM.N_287\
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__4463\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_1_0_cascade_\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__4460\,
            I => \U712_CHIP_RAM.N_273_cascade_\
        );

    \I__590\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4452\
        );

    \I__589\ : InMux
    port map (
            O => \N__4456\,
            I => \N__4449\
        );

    \I__588\ : InMux
    port map (
            O => \N__4455\,
            I => \N__4446\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4452\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4449\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__4446\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3\
        );

    \I__584\ : InMux
    port map (
            O => \N__4439\,
            I => \N__4436\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__4436\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_0\
        );

    \I__582\ : InMux
    port map (
            O => \N__4433\,
            I => \N__4429\
        );

    \I__581\ : CascadeMux
    port map (
            O => \N__4432\,
            I => \N__4425\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4429\,
            I => \N__4421\
        );

    \I__579\ : InMux
    port map (
            O => \N__4428\,
            I => \N__4414\
        );

    \I__578\ : InMux
    port map (
            O => \N__4425\,
            I => \N__4414\
        );

    \I__577\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4414\
        );

    \I__576\ : Span4Mux_v
    port map (
            O => \N__4421\,
            I => \N__4411\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4414\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__574\ : Odrv4
    port map (
            O => \N__4411\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__573\ : InMux
    port map (
            O => \N__4406\,
            I => \N__4403\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4403\,
            I => \N__4398\
        );

    \I__571\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4393\
        );

    \I__570\ : InMux
    port map (
            O => \N__4401\,
            I => \N__4393\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__4398\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4393\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__4388\,
            I => \N__4384\
        );

    \I__566\ : CascadeMux
    port map (
            O => \N__4387\,
            I => \N__4381\
        );

    \I__565\ : InMux
    port map (
            O => \N__4384\,
            I => \N__4376\
        );

    \I__564\ : InMux
    port map (
            O => \N__4381\,
            I => \N__4376\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4376\,
            I => \U712_REG_SM.LDS_OUT_2_0_a2Z0Z_0\
        );

    \I__562\ : CascadeMux
    port map (
            O => \N__4373\,
            I => \N__4370\
        );

    \I__561\ : InMux
    port map (
            O => \N__4370\,
            I => \N__4367\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4367\,
            I => \N__4360\
        );

    \I__559\ : InMux
    port map (
            O => \N__4366\,
            I => \N__4357\
        );

    \I__558\ : InMux
    port map (
            O => \N__4365\,
            I => \N__4350\
        );

    \I__557\ : InMux
    port map (
            O => \N__4364\,
            I => \N__4350\
        );

    \I__556\ : InMux
    port map (
            O => \N__4363\,
            I => \N__4350\
        );

    \I__555\ : Odrv4
    port map (
            O => \N__4360\,
            I => \U712_REG_SM.N_342\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__4357\,
            I => \U712_REG_SM.N_342\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__4350\,
            I => \U712_REG_SM.N_342\
        );

    \I__552\ : InMux
    port map (
            O => \N__4343\,
            I => \N__4339\
        );

    \I__551\ : InMux
    port map (
            O => \N__4342\,
            I => \N__4336\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4339\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4336\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__548\ : IoInMux
    port map (
            O => \N__4331\,
            I => \N__4328\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4328\,
            I => \N__4325\
        );

    \I__546\ : IoSpan4Mux
    port map (
            O => \N__4325\,
            I => \N__4322\
        );

    \I__545\ : Span4Mux_s3_v
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__544\ : Span4Mux_h
    port map (
            O => \N__4319\,
            I => \N__4316\
        );

    \I__543\ : Sp12to4
    port map (
            O => \N__4316\,
            I => \N__4313\
        );

    \I__542\ : Span12Mux_v
    port map (
            O => \N__4313\,
            I => \N__4310\
        );

    \I__541\ : Odrv12
    port map (
            O => \N__4310\,
            I => \U712_REG_SM_un1_LDSn_i\
        );

    \I__540\ : InMux
    port map (
            O => \N__4307\,
            I => \N__4304\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__4304\,
            I => \N__4300\
        );

    \I__538\ : InMux
    port map (
            O => \N__4303\,
            I => \N__4297\
        );

    \I__537\ : Odrv4
    port map (
            O => \N__4300\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4297\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__535\ : InMux
    port map (
            O => \N__4292\,
            I => \N__4288\
        );

    \I__534\ : InMux
    port map (
            O => \N__4291\,
            I => \N__4285\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__4288\,
            I => \N__4281\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__4285\,
            I => \N__4278\
        );

    \I__531\ : InMux
    port map (
            O => \N__4284\,
            I => \N__4275\
        );

    \I__530\ : Odrv12
    port map (
            O => \N__4281\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__529\ : Odrv4
    port map (
            O => \N__4278\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__4275\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__527\ : IoInMux
    port map (
            O => \N__4268\,
            I => \N__4265\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4265\,
            I => \N__4262\
        );

    \I__525\ : IoSpan4Mux
    port map (
            O => \N__4262\,
            I => \N__4259\
        );

    \I__524\ : IoSpan4Mux
    port map (
            O => \N__4259\,
            I => \N__4256\
        );

    \I__523\ : Sp12to4
    port map (
            O => \N__4256\,
            I => \N__4253\
        );

    \I__522\ : Span12Mux_v
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__521\ : Odrv12
    port map (
            O => \N__4250\,
            I => \U712_REG_SM_un1_UDSn_i\
        );

    \I__520\ : CascadeMux
    port map (
            O => \N__4247\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_\
        );

    \I__519\ : CascadeMux
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__518\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4238\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4238\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6\
        );

    \I__516\ : InMux
    port map (
            O => \N__4235\,
            I => \N__4231\
        );

    \I__515\ : InMux
    port map (
            O => \N__4234\,
            I => \N__4228\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__4231\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4228\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__512\ : InMux
    port map (
            O => \N__4223\,
            I => \N__4218\
        );

    \I__511\ : InMux
    port map (
            O => \N__4222\,
            I => \N__4215\
        );

    \I__510\ : InMux
    port map (
            O => \N__4221\,
            I => \N__4212\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4218\,
            I => \N__4209\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4215\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__4212\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__506\ : Odrv4
    port map (
            O => \N__4209\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__505\ : CascadeMux
    port map (
            O => \N__4202\,
            I => \N__4197\
        );

    \I__504\ : InMux
    port map (
            O => \N__4201\,
            I => \N__4192\
        );

    \I__503\ : InMux
    port map (
            O => \N__4200\,
            I => \N__4192\
        );

    \I__502\ : InMux
    port map (
            O => \N__4197\,
            I => \N__4189\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__4192\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4189\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__4184\,
            I => \N__4181\
        );

    \I__498\ : InMux
    port map (
            O => \N__4181\,
            I => \N__4175\
        );

    \I__497\ : InMux
    port map (
            O => \N__4180\,
            I => \N__4172\
        );

    \I__496\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4169\
        );

    \I__495\ : InMux
    port map (
            O => \N__4178\,
            I => \N__4166\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4175\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__4172\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__4169\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4166\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__489\ : InMux
    port map (
            O => \N__4154\,
            I => \N__4150\
        );

    \I__488\ : InMux
    port map (
            O => \N__4153\,
            I => \N__4147\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4150\,
            I => \REG_TACK\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__4147\,
            I => \REG_TACK\
        );

    \I__485\ : InMux
    port map (
            O => \N__4142\,
            I => \N__4139\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4139\,
            I => \N__4135\
        );

    \I__483\ : InMux
    port map (
            O => \N__4138\,
            I => \N__4132\
        );

    \I__482\ : Span4Mux_v
    port map (
            O => \N__4135\,
            I => \N__4127\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4132\,
            I => \N__4127\
        );

    \I__480\ : Span4Mux_v
    port map (
            O => \N__4127\,
            I => \N__4124\
        );

    \I__479\ : Span4Mux_v
    port map (
            O => \N__4124\,
            I => \N__4121\
        );

    \I__478\ : Sp12to4
    port map (
            O => \N__4121\,
            I => \N__4118\
        );

    \I__477\ : Span12Mux_h
    port map (
            O => \N__4118\,
            I => \N__4115\
        );

    \I__476\ : Odrv12
    port map (
            O => \N__4115\,
            I => \TSn_c\
        );

    \I__475\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4109\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4109\,
            I => \N__4106\
        );

    \I__473\ : Span4Mux_v
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__472\ : Sp12to4
    port map (
            O => \N__4103\,
            I => \N__4100\
        );

    \I__471\ : Span12Mux_h
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__470\ : Span12Mux_v
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__469\ : Odrv12
    port map (
            O => \N__4094\,
            I => \REGSPACEn_c\
        );

    \I__468\ : InMux
    port map (
            O => \N__4091\,
            I => \N__4085\
        );

    \I__467\ : InMux
    port map (
            O => \N__4090\,
            I => \N__4085\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4085\,
            I => \U712_REG_SM.REG_CYCLE_GOZ0\
        );

    \I__465\ : InMux
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4079\,
            I => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1\
        );

    \I__463\ : CascadeMux
    port map (
            O => \N__4076\,
            I => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__4073\,
            I => \N__4070\
        );

    \I__461\ : InMux
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4067\,
            I => \N__4064\
        );

    \I__459\ : Span4Mux_v
    port map (
            O => \N__4064\,
            I => \N__4061\
        );

    \I__458\ : Sp12to4
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__457\ : Span12Mux_h
    port map (
            O => \N__4058\,
            I => \N__4055\
        );

    \I__456\ : Span12Mux_v
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__455\ : Odrv12
    port map (
            O => \N__4052\,
            I => \RAMSPACEn_c\
        );

    \I__454\ : InMux
    port map (
            O => \N__4049\,
            I => \N__4046\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__4046\,
            I => \N__4043\
        );

    \I__452\ : Span4Mux_v
    port map (
            O => \N__4043\,
            I => \N__4040\
        );

    \I__451\ : Sp12to4
    port map (
            O => \N__4040\,
            I => \N__4037\
        );

    \I__450\ : Span12Mux_h
    port map (
            O => \N__4037\,
            I => \N__4034\
        );

    \I__449\ : Span12Mux_v
    port map (
            O => \N__4034\,
            I => \N__4031\
        );

    \I__448\ : Odrv12
    port map (
            O => \N__4031\,
            I => \DBRn_c\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__4028\,
            I => \U712_CHIP_RAM.N_287_cascade_\
        );

    \I__446\ : InMux
    port map (
            O => \N__4025\,
            I => \N__4022\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4022\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_1_0\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__4019\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_cascade_\
        );

    \I__443\ : CascadeMux
    port map (
            O => \N__4016\,
            I => \N__4013\
        );

    \I__442\ : InMux
    port map (
            O => \N__4013\,
            I => \N__4006\
        );

    \I__441\ : InMux
    port map (
            O => \N__4012\,
            I => \N__4006\
        );

    \I__440\ : InMux
    port map (
            O => \N__4011\,
            I => \N__4003\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4006\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__4003\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__437\ : InMux
    port map (
            O => \N__3998\,
            I => \N__3994\
        );

    \I__436\ : InMux
    port map (
            O => \N__3997\,
            I => \N__3991\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__3994\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3991\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__433\ : InMux
    port map (
            O => \N__3986\,
            I => \N__3983\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__3983\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__431\ : CascadeMux
    port map (
            O => \N__3980\,
            I => \U712_CYCLE_TERM.N_307_i_0_en_cascade_\
        );

    \I__430\ : InMux
    port map (
            O => \N__3977\,
            I => \N__3972\
        );

    \I__429\ : InMux
    port map (
            O => \N__3976\,
            I => \N__3967\
        );

    \I__428\ : InMux
    port map (
            O => \N__3975\,
            I => \N__3967\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3972\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__3967\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__3962\,
            I => \N__3958\
        );

    \I__424\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3955\
        );

    \I__423\ : InMux
    port map (
            O => \N__3958\,
            I => \N__3951\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3955\,
            I => \N__3948\
        );

    \I__421\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3945\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3951\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__419\ : Odrv4
    port map (
            O => \N__3948\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3945\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__417\ : InMux
    port map (
            O => \N__3938\,
            I => \N__3935\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3935\,
            I => \N__3932\
        );

    \I__415\ : Sp12to4
    port map (
            O => \N__3932\,
            I => \N__3929\
        );

    \I__414\ : Odrv12
    port map (
            O => \N__3929\,
            I => \TACK_EN_i_ess\
        );

    \I__413\ : CEMux
    port map (
            O => \N__3926\,
            I => \N__3923\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__3923\,
            I => \N__3920\
        );

    \I__411\ : Odrv12
    port map (
            O => \N__3920\,
            I => \U712_CYCLE_TERM.N_307_i_0_en_0\
        );

    \I__410\ : IoInMux
    port map (
            O => \N__3917\,
            I => \N__3914\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3914\,
            I => \N__3911\
        );

    \I__408\ : Span12Mux_s2_v
    port map (
            O => \N__3911\,
            I => \N__3908\
        );

    \I__407\ : Odrv12
    port map (
            O => \N__3908\,
            I => \VBENn_c\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__3905\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3_cascade_\
        );

    \I__405\ : CascadeMux
    port map (
            O => \N__3902\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_\
        );

    \I__404\ : InMux
    port map (
            O => \N__3899\,
            I => \N__3896\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__3896\,
            I => \U712_CHIP_RAM.N_181\
        );

    \I__402\ : InMux
    port map (
            O => \N__3893\,
            I => \N__3883\
        );

    \I__401\ : InMux
    port map (
            O => \N__3892\,
            I => \N__3883\
        );

    \I__400\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3883\
        );

    \I__399\ : InMux
    port map (
            O => \N__3890\,
            I => \N__3880\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3883\,
            I => \N__3877\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__3880\,
            I => \N__3872\
        );

    \I__396\ : Span4Mux_v
    port map (
            O => \N__3877\,
            I => \N__3872\
        );

    \I__395\ : Span4Mux_v
    port map (
            O => \N__3872\,
            I => \N__3869\
        );

    \I__394\ : Sp12to4
    port map (
            O => \N__3869\,
            I => \N__3866\
        );

    \I__393\ : Span12Mux_h
    port map (
            O => \N__3866\,
            I => \N__3863\
        );

    \I__392\ : Odrv12
    port map (
            O => \N__3863\,
            I => \CLK40_OUT_i\
        );

    \I__391\ : IoInMux
    port map (
            O => \N__3860\,
            I => \N__3857\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3857\,
            I => \N__3854\
        );

    \I__389\ : Span12Mux_s8_h
    port map (
            O => \N__3854\,
            I => \N__3851\
        );

    \I__388\ : Span12Mux_v
    port map (
            O => \N__3851\,
            I => \N__3847\
        );

    \I__387\ : InMux
    port map (
            O => \N__3850\,
            I => \N__3844\
        );

    \I__386\ : Odrv12
    port map (
            O => \N__3847\,
            I => \TACK_OUTn\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__3844\,
            I => \TACK_OUTn\
        );

    \I__384\ : InMux
    port map (
            O => \N__3839\,
            I => \N__3827\
        );

    \I__383\ : InMux
    port map (
            O => \N__3838\,
            I => \N__3827\
        );

    \I__382\ : InMux
    port map (
            O => \N__3837\,
            I => \N__3827\
        );

    \I__381\ : InMux
    port map (
            O => \N__3836\,
            I => \N__3827\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__3827\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__379\ : InMux
    port map (
            O => \N__3824\,
            I => \N__3820\
        );

    \I__378\ : InMux
    port map (
            O => \N__3823\,
            I => \N__3817\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__3820\,
            I => \CPU_TACKm\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__3817\,
            I => \CPU_TACKm\
        );

    \I__375\ : CascadeMux
    port map (
            O => \N__3812\,
            I => \N__3809\
        );

    \I__374\ : InMux
    port map (
            O => \N__3809\,
            I => \N__3805\
        );

    \I__373\ : InMux
    port map (
            O => \N__3808\,
            I => \N__3802\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3805\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__3802\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__370\ : CascadeMux
    port map (
            O => \N__3797\,
            I => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\
        );

    \I__369\ : InMux
    port map (
            O => \N__3794\,
            I => \N__3791\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3791\,
            I => \N__3788\
        );

    \I__367\ : Span4Mux_v
    port map (
            O => \N__3788\,
            I => \N__3785\
        );

    \I__366\ : Sp12to4
    port map (
            O => \N__3785\,
            I => \N__3782\
        );

    \I__365\ : Odrv12
    port map (
            O => \N__3782\,
            I => \A_c_13\
        );

    \I__364\ : CascadeMux
    port map (
            O => \N__3779\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4_cascade_\
        );

    \I__363\ : InMux
    port map (
            O => \N__3776\,
            I => \N__3773\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__3773\,
            I => \N__3770\
        );

    \I__361\ : Span4Mux_h
    port map (
            O => \N__3770\,
            I => \N__3767\
        );

    \I__360\ : Sp12to4
    port map (
            O => \N__3767\,
            I => \N__3764\
        );

    \I__359\ : Span12Mux_v
    port map (
            O => \N__3764\,
            I => \N__3761\
        );

    \I__358\ : Odrv12
    port map (
            O => \N__3761\,
            I => \A_c_6\
        );

    \I__357\ : IoInMux
    port map (
            O => \N__3758\,
            I => \N__3755\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__3755\,
            I => \N__3752\
        );

    \I__355\ : Span12Mux_s9_h
    port map (
            O => \N__3752\,
            I => \N__3749\
        );

    \I__354\ : Span12Mux_h
    port map (
            O => \N__3749\,
            I => \N__3746\
        );

    \I__353\ : Odrv12
    port map (
            O => \N__3746\,
            I => \CMA_c_3\
        );

    \I__352\ : InMux
    port map (
            O => \N__3743\,
            I => \N__3740\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__3740\,
            I => \U712_CHIP_RAM.N_319\
        );

    \I__350\ : IoInMux
    port map (
            O => \N__3737\,
            I => \N__3734\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__3734\,
            I => \N__3731\
        );

    \I__348\ : Span4Mux_s2_h
    port map (
            O => \N__3731\,
            I => \N__3728\
        );

    \I__347\ : Span4Mux_v
    port map (
            O => \N__3728\,
            I => \N__3725\
        );

    \I__346\ : Span4Mux_v
    port map (
            O => \N__3725\,
            I => \N__3722\
        );

    \I__345\ : Sp12to4
    port map (
            O => \N__3722\,
            I => \N__3719\
        );

    \I__344\ : Span12Mux_s11_h
    port map (
            O => \N__3719\,
            I => \N__3716\
        );

    \I__343\ : Odrv12
    port map (
            O => \N__3716\,
            I => \CMA_c_4\
        );

    \I__342\ : InMux
    port map (
            O => \N__3713\,
            I => \N__3710\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__3710\,
            I => \N__3707\
        );

    \I__340\ : Span4Mux_v
    port map (
            O => \N__3707\,
            I => \N__3704\
        );

    \I__339\ : Sp12to4
    port map (
            O => \N__3704\,
            I => \N__3701\
        );

    \I__338\ : Odrv12
    port map (
            O => \N__3701\,
            I => \A_c_12\
        );

    \I__337\ : CascadeMux
    port map (
            O => \N__3698\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_\
        );

    \I__336\ : InMux
    port map (
            O => \N__3695\,
            I => \N__3692\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__3692\,
            I => \N__3689\
        );

    \I__334\ : Sp12to4
    port map (
            O => \N__3689\,
            I => \N__3686\
        );

    \I__333\ : Span12Mux_v
    port map (
            O => \N__3686\,
            I => \N__3683\
        );

    \I__332\ : Odrv12
    port map (
            O => \N__3683\,
            I => \A_c_5\
        );

    \I__331\ : InMux
    port map (
            O => \N__3680\,
            I => \N__3677\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__3677\,
            I => \U712_CHIP_RAM.N_318\
        );

    \I__329\ : IoInMux
    port map (
            O => \N__3674\,
            I => \N__3671\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__3671\,
            I => \N__3668\
        );

    \I__327\ : Span4Mux_s3_h
    port map (
            O => \N__3668\,
            I => \N__3665\
        );

    \I__326\ : Span4Mux_h
    port map (
            O => \N__3665\,
            I => \N__3662\
        );

    \I__325\ : Span4Mux_v
    port map (
            O => \N__3662\,
            I => \N__3659\
        );

    \I__324\ : Odrv4
    port map (
            O => \N__3659\,
            I => \CLK40_OUT_i_i\
        );

    \I__323\ : CascadeMux
    port map (
            O => \N__3656\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_0_a2_i_0_cascade_\
        );

    \I__322\ : IoInMux
    port map (
            O => \N__3653\,
            I => \N__3650\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__3650\,
            I => \N__3647\
        );

    \I__320\ : IoSpan4Mux
    port map (
            O => \N__3647\,
            I => \N__3644\
        );

    \I__319\ : Span4Mux_s2_v
    port map (
            O => \N__3644\,
            I => \N__3641\
        );

    \I__318\ : Span4Mux_v
    port map (
            O => \N__3641\,
            I => \N__3638\
        );

    \I__317\ : Odrv4
    port map (
            O => \N__3638\,
            I => \CLK80_OUT_i_i\
        );

    \I__316\ : IoInMux
    port map (
            O => \N__3635\,
            I => \N__3632\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__3632\,
            I => \N__3629\
        );

    \I__314\ : IoSpan4Mux
    port map (
            O => \N__3629\,
            I => \N__3626\
        );

    \I__313\ : Span4Mux_s3_h
    port map (
            O => \N__3626\,
            I => \N__3623\
        );

    \I__312\ : Span4Mux_h
    port map (
            O => \N__3623\,
            I => \N__3620\
        );

    \I__311\ : Odrv4
    port map (
            O => \N__3620\,
            I => \N_839_i\
        );

    \I__310\ : IoInMux
    port map (
            O => \N__3617\,
            I => \N__3614\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__3614\,
            I => \N__3611\
        );

    \I__308\ : IoSpan4Mux
    port map (
            O => \N__3611\,
            I => \N__3608\
        );

    \I__307\ : Span4Mux_s2_v
    port map (
            O => \N__3608\,
            I => \N__3605\
        );

    \I__306\ : Sp12to4
    port map (
            O => \N__3605\,
            I => \N__3602\
        );

    \I__305\ : Span12Mux_v
    port map (
            O => \N__3602\,
            I => \N__3599\
        );

    \I__304\ : Odrv12
    port map (
            O => \N__3599\,
            I => \CLK40_IN_c\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_8_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7634\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6169\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9248\,
            lcout => \CLK80_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3938\,
            lcout => \N_839_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010011"
        )
    port map (
            in0 => \N__7583\,
            in1 => \N__6818\,
            in2 => \N__8521\,
            in3 => \N__8134\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8135\,
            in1 => \N__3794\,
            in2 => \N__3779\,
            in3 => \N__3776\,
            lcout => \U712_CHIP_RAM.N_319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__3680\,
            in1 => \_gnd_net_\,
            in2 => \N__8641\,
            in3 => \N__8756\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9231\,
            ce => \N__7967\,
            sr => \N__9046\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__8755\,
            in1 => \N__8631\,
            in2 => \_gnd_net_\,
            in3 => \N__3743\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9231\,
            ce => \N__7967\,
            sr => \N__9046\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__8507\,
            in1 => \N__7880\,
            in2 => \N__8169\,
            in3 => \N__7466\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8158\,
            in1 => \N__3713\,
            in2 => \N__3698\,
            in3 => \N__3695\,
            lcout => \U712_CHIP_RAM.N_318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK40C_obuf_RNO_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3890\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110111011"
        )
    port map (
            in0 => \N__5800\,
            in1 => \N__5656\,
            in2 => \_gnd_net_\,
            in3 => \N__5349\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_0_a2_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5267\,
            in1 => \N__7203\,
            in2 => \N__3656\,
            in3 => \N__5096\,
            lcout => \U712_CHIP_RAM.N_181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__3837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3893\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9239\,
            ce => 'H',
            sr => \N__9019\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000110000"
        )
    port map (
            in0 => \N__3891\,
            in1 => \N__3976\,
            in2 => \N__3962\,
            in3 => \N__3839\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9239\,
            ce => 'H',
            sr => \N__9019\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3998\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9239\,
            ce => 'H',
            sr => \N__9019\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__3824\,
            in1 => \N__5801\,
            in2 => \N__8174\,
            in3 => \N__3899\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9239\,
            ce => 'H',
            sr => \N__9019\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4012\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9239\,
            ce => 'H',
            sr => \N__9019\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110011110100"
        )
    port map (
            in0 => \N__3838\,
            in1 => \N__3850\,
            in2 => \N__4016\,
            in3 => \N__3892\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9239\,
            ce => 'H',
            sr => \N__9019\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__3986\,
            in1 => \N__3975\,
            in2 => \N__3812\,
            in3 => \N__3836\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9239\,
            ce => 'H',
            sr => \N__9019\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4153\,
            in2 => \_gnd_net_\,
            in3 => \N__3823\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__7701\,
            in1 => \N__3808\,
            in2 => \N__3797\,
            in3 => \N__3954\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_307_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9083\,
            in1 => \_gnd_net_\,
            in2 => \N__3980\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.N_307_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__7691\,
            in1 => \N__3977\,
            in2 => \_gnd_net_\,
            in3 => \N__3961\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9243\,
            ce => \N__3926\,
            sr => \N__9004\
        );

    \U712_REG_SM.LDS_OUT_2_0_a2_0_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6058\,
            in2 => \_gnd_net_\,
            in3 => \N__4997\,
            lcout => \U712_REG_SM.LDS_OUT_2_0_a2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__4457\,
            in1 => \N__9089\,
            in2 => \N__4184\,
            in3 => \N__5090\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4745\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8137\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__5731\,
            in1 => \N__5325\,
            in2 => \_gnd_net_\,
            in3 => \N__5605\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5606\,
            in1 => \N__5334\,
            in2 => \_gnd_net_\,
            in3 => \N__5732\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__4222\,
            in1 => \N__4180\,
            in2 => \N__3905\,
            in3 => \N__5089\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3902\,
            in3 => \N__9086\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__4533\,
            in1 => \N__4558\,
            in2 => \N__5446\,
            in3 => \N__5406\,
            lcout => \U712_CHIP_RAM.N_272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101011"
        )
    port map (
            in0 => \N__5442\,
            in1 => \N__4142\,
            in2 => \N__4073\,
            in3 => \N__8162\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9232\,
            ce => 'H',
            sr => \N__9030\
        );

    \U712_CHIP_RAM.DBR_SYNC_0_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4049\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM_DBR_SYNC_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9232\,
            ce => 'H',
            sr => \N__9030\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__4557\,
            in1 => \N__4532\,
            in2 => \_gnd_net_\,
            in3 => \N__5438\,
            lcout => \U712_CHIP_RAM.N_287\,
            ltout => \U712_CHIP_RAM.N_287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRB433_1_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5614\,
            in1 => \N__4439\,
            in2 => \N__4028\,
            in3 => \N__5736\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVNIQ6_3_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4025\,
            in1 => \N__7177\,
            in2 => \N__4019\,
            in3 => \N__5081\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4537\,
            lcout => \U712_REG_SM_DBR_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9234\,
            ce => 'H',
            sr => \N__9024\
        );

    \U712_CHIP_RAM.DBDIR_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000001110100"
        )
    port map (
            in0 => \N__4489\,
            in1 => \N__7000\,
            in2 => \N__4614\,
            in3 => \N__6976\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9234\,
            ce => 'H',
            sr => \N__9024\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4011\,
            in2 => \_gnd_net_\,
            in3 => \N__3997\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101010000"
        )
    port map (
            in0 => \N__4832\,
            in1 => \N__4800\,
            in2 => \N__4157\,
            in3 => \N__4782\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9240\,
            ce => 'H',
            sr => \N__9005\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110011"
        )
    port map (
            in0 => \N__4091\,
            in1 => \N__4138\,
            in2 => \N__4432\,
            in3 => \N__4112\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9240\,
            ce => 'H',
            sr => \N__9005\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__4945\,
            in1 => \N__4366\,
            in2 => \_gnd_net_\,
            in3 => \N__6322\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9240\,
            ce => 'H',
            sr => \N__9005\
        );

    \U712_REG_SM.DS_EN_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__4284\,
            in1 => \N__4928\,
            in2 => \N__4955\,
            in3 => \N__4082\,
            lcout => \U712_REG_SM.DS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9240\,
            ce => 'H',
            sr => \N__9005\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__4424\,
            in1 => \N__4402\,
            in2 => \N__5018\,
            in3 => \N__6373\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9240\,
            ce => 'H',
            sr => \N__9005\
        );

    \U712_REG_SM.REG_CYCLE_GO_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__4401\,
            in1 => \N__4090\,
            in2 => \N__4373\,
            in3 => \N__4428\,
            lcout => \U712_REG_SM.REG_CYCLE_GOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9240\,
            ce => 'H',
            sr => \N__9005\
        );

    \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000001"
        )
    port map (
            in0 => \N__6387\,
            in1 => \N__4678\,
            in2 => \N__6374\,
            in3 => \N__5014\,
            lcout => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1\,
            ltout => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_1_ess_RNO_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4076\,
            in3 => \N__9081\,
            lcout => \U712_REG_SM.N_186_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4679\,
            in1 => \N__6371\,
            in2 => \_gnd_net_\,
            in3 => \N__6388\,
            lcout => \U712_REG_SM.N_342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDS_OUT_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101111"
        )
    port map (
            in0 => \N__6203\,
            in1 => \N__4342\,
            in2 => \N__4387\,
            in3 => \N__4364\,
            lcout => \U712_REG_SM.LDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9244\,
            ce => 'H',
            sr => \N__8994\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__4363\,
            in1 => \N__4433\,
            in2 => \N__4694\,
            in3 => \N__4406\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9244\,
            ce => 'H',
            sr => \N__8994\
        );

    \U712_REG_SM.UDS_OUT_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011111"
        )
    port map (
            in0 => \N__6204\,
            in1 => \N__4303\,
            in2 => \N__4388\,
            in3 => \N__4365\,
            lcout => \U712_REG_SM.UDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9244\,
            ce => 'H',
            sr => \N__8994\
        );

    \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4291\,
            in2 => \_gnd_net_\,
            in3 => \N__4343\,
            lcout => \U712_REG_SM_un1_LDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_RNIUP9B_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__4307\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4292\,
            lcout => \U712_REG_SM_un1_UDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__5637\,
            in1 => \N__5339\,
            in2 => \N__5799\,
            in3 => \N__5160\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4221\,
            in1 => \N__4179\,
            in2 => \N__5095\,
            in3 => \N__4455\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__9087\,
            in1 => \_gnd_net_\,
            in2 => \N__4247\,
            in3 => \N__4201\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__4200\,
            in1 => \N__9088\,
            in2 => \N__4244\,
            in3 => \N__4235\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4234\,
            in1 => \N__4223\,
            in2 => \N__4202\,
            in3 => \N__4178\,
            lcout => \U712_CHIP_RAM.N_276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5798\,
            in1 => \N__5642\,
            in2 => \_gnd_net_\,
            in3 => \N__5161\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__5261\,
            in1 => \N__5402\,
            in2 => \_gnd_net_\,
            in3 => \N__4469\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100111"
        )
    port map (
            in0 => \N__6962\,
            in1 => \N__5742\,
            in2 => \N__4463\,
            in3 => \N__5171\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5323\,
            in2 => \_gnd_net_\,
            in3 => \N__5074\,
            lcout => \U712_CHIP_RAM.N_273\,
            ltout => \U712_CHIP_RAM.N_273_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINN5O1_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5741\,
            in2 => \N__4460\,
            in3 => \N__7127\,
            lcout => \U712_CHIP_RAM.N_296_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5162\,
            in1 => \N__4456\,
            in2 => \_gnd_net_\,
            in3 => \N__5075\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICGJU_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5324\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5391\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000100"
        )
    port map (
            in0 => \N__5616\,
            in1 => \N__7114\,
            in2 => \N__5781\,
            in3 => \N__5817\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_0_a2_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7178\,
            in2 => \_gnd_net_\,
            in3 => \N__7708\,
            lcout => \U712_CHIP_RAM.N_347\,
            ltout => \U712_CHIP_RAM.N_347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHBQU6_0_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__5737\,
            in1 => \N__7216\,
            in2 => \N__4514\,
            in3 => \N__5465\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_378_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI8KLPE_0_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__5262\,
            in1 => \N__7709\,
            in2 => \N__4511\,
            in3 => \N__4508\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__7179\,
            in1 => \_gnd_net_\,
            in2 => \N__5541\,
            in3 => \N__4502\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011111010"
        )
    port map (
            in0 => \N__5110\,
            in1 => \_gnd_net_\,
            in2 => \N__4496\,
            in3 => \N__6975\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9228\,
            ce => 'H',
            sr => \N__9025\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5419\,
            in2 => \_gnd_net_\,
            in3 => \N__5109\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER50\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER50_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__7113\,
            in1 => \N__5615\,
            in2 => \N__4493\,
            in3 => \N__5531\,
            lcout => \U712_CHIP_RAM.N_424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_3_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011111111"
        )
    port map (
            in0 => \N__5792\,
            in1 => \N__7129\,
            in2 => \N__5658\,
            in3 => \N__4657\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000101101"
        )
    port map (
            in0 => \N__7128\,
            in1 => \N__5819\,
            in2 => \N__5657\,
            in3 => \N__5793\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__5003\,
            in1 => \N__4490\,
            in2 => \_gnd_net_\,
            in3 => \N__5395\,
            lcout => \U712_CHIP_RAM.N_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_sbtinv_3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5492\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5263\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5196\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100011111111"
        )
    port map (
            in0 => \N__5794\,
            in1 => \N__7130\,
            in2 => \N__5659\,
            in3 => \N__4658\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_e_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000110010"
        )
    port map (
            in0 => \N__5850\,
            in1 => \N__5493\,
            in2 => \N__4646\,
            in3 => \N__8717\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9233\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_3_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__5851\,
            in1 => \N__5660\,
            in2 => \N__4643\,
            in3 => \N__5510\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9235\,
            ce => \N__4634\,
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__4783\,
            in1 => \N__6350\,
            in2 => \N__4807\,
            in3 => \N__4834\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9236\,
            ce => 'H',
            sr => \N__9006\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101010000"
        )
    port map (
            in0 => \N__4667\,
            in1 => \N__6349\,
            in2 => \N__4922\,
            in3 => \N__4833\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9236\,
            ce => 'H',
            sr => \N__9006\
        );

    \U712_BUFFERS.DRDDIR_i_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__4737\,
            in1 => \N__5982\,
            in2 => \N__4621\,
            in3 => \N__4999\,
            lcout => \N_188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__6337\,
            in1 => \N__6577\,
            in2 => \_gnd_net_\,
            in3 => \N__6532\,
            lcout => \U712_REG_SM.N_288\,
            ltout => \U712_REG_SM.N_288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4565\,
            in2 => \N__4544\,
            in3 => \N__4541\,
            lcout => \U712_REG_SM.N_301\,
            ltout => \U712_REG_SM.N_301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001100"
        )
    port map (
            in0 => \N__4835\,
            in1 => \N__4756\,
            in2 => \N__4811\,
            in3 => \N__4736\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9237\,
            ce => 'H',
            sr => \N__8998\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__4766\,
            in1 => \N__4784\,
            in2 => \N__4808\,
            in3 => \N__4757\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9237\,
            ce => 'H',
            sr => \N__8998\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000000000"
        )
    port map (
            in0 => \N__4755\,
            in1 => \N__4946\,
            in2 => \N__6323\,
            in3 => \N__4765\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9237\,
            ce => 'H',
            sr => \N__8998\
        );

    \U712_BUFFERS.un1_DRDENn_0_a2_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5983\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4738\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__6575\,
            in1 => \_gnd_net_\,
            in2 => \N__6531\,
            in3 => \N__4690\,
            lcout => \U712_REG_SM.N_341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__6552\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6125\,
            lcout => \U712_REG_SM.N_294\,
            ltout => \U712_REG_SM.N_294_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6405\,
            in1 => \N__6606\,
            in2 => \N__4670\,
            in3 => \N__6640\,
            lcout => \U712_REG_SM.N_373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6574\,
            in2 => \_gnd_net_\,
            in3 => \N__6519\,
            lcout => \U712_REG_SM.N_292\,
            ltout => \U712_REG_SM.N_292_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4920\,
            in1 => \N__6605\,
            in2 => \N__5021\,
            in3 => \N__6639\,
            lcout => \U712_REG_SM.N_507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__6553\,
            in1 => \N__6644\,
            in2 => \_gnd_net_\,
            in3 => \N__4998\,
            lcout => \U712_REG_SM.N_104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6604\,
            in2 => \_gnd_net_\,
            in3 => \N__6638\,
            lcout => \U712_REG_SM.N_298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4944\,
            in1 => \N__6576\,
            in2 => \N__6341\,
            in3 => \N__6523\,
            lcout => \U712_REG_SM.N_372\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_1_ess_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4921\,
            in1 => \N__6645\,
            in2 => \N__6410\,
            in3 => \N__6607\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9242\,
            ce => \N__4856\,
            sr => \N__8992\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__5259\,
            in1 => \N__6955\,
            in2 => \N__4844\,
            in3 => \N__5204\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__8063\,
            in1 => \N__6963\,
            in2 => \N__4850\,
            in3 => \N__5408\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9210\,
            ce => 'H',
            sr => \N__9031\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNO_2_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5613\,
            in1 => \N__5746\,
            in2 => \N__5353\,
            in3 => \N__8062\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNO_1_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5085\,
            in1 => \N__5257\,
            in2 => \N__4847\,
            in3 => \N__7189\,
            lcout => \U712_CHIP_RAM.N_393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJV8G1_2_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100000010000"
        )
    port map (
            in0 => \N__5611\,
            in1 => \N__5327\,
            in2 => \N__5091\,
            in3 => \N__8061\,
            lcout => \U712_CHIP_RAM.N_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6IFV8_0_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__7181\,
            in1 => \N__9084\,
            in2 => \N__5783\,
            in3 => \N__5453\,
            lcout => \U712_CHIP_RAM.N_310\,
            ltout => \U712_CHIP_RAM.N_310_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIDCLTE_0_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111110"
        )
    port map (
            in0 => \N__5258\,
            in1 => \N__5203\,
            in2 => \N__5165\,
            in3 => \N__6954\,
            lcout => \U712_CHIP_RAM.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_10_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7180\,
            in1 => \N__5612\,
            in2 => \N__5782\,
            in3 => \N__5535\,
            lcout => \U712_CHIP_RAM.N_293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111110"
        )
    port map (
            in0 => \N__5247\,
            in1 => \N__5734\,
            in2 => \N__5638\,
            in3 => \N__5338\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_3_0_a2_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7193\,
            in2 => \N__5147\,
            in3 => \N__5077\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_179_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010110010101111"
        )
    port map (
            in0 => \N__5122\,
            in1 => \N__6914\,
            in2 => \N__5144\,
            in3 => \N__5735\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9215\,
            ce => 'H',
            sr => \N__9026\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__7097\,
            in1 => \N__5420\,
            in2 => \_gnd_net_\,
            in3 => \N__5111\,
            lcout => \U712_CHIP_RAM.N_284\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5607\,
            in2 => \_gnd_net_\,
            in3 => \N__5076\,
            lcout => \U712_CHIP_RAM.N_438\,
            ltout => \U712_CHIP_RAM.N_438_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNILE372_2_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5326\,
            in1 => \N__7098\,
            in2 => \N__5024\,
            in3 => \N__5733\,
            lcout => \U712_CHIP_RAM.N_425\,
            ltout => \U712_CHIP_RAM.N_425_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI94U46_2_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__5474\,
            in1 => \N__5246\,
            in2 => \N__5468\,
            in3 => \N__5464\,
            lcout => \U712_CHIP_RAM.N_302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001100"
        )
    port map (
            in0 => \N__5958\,
            in1 => \N__8786\,
            in2 => \N__8813\,
            in3 => \N__5401\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9224\,
            ce => 'H',
            sr => \N__9020\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNO_0_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5397\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5447\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH_CYCLE_START_2_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5959\,
            in1 => \N__6875\,
            in2 => \N__5423\,
            in3 => \N__8132\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9224\,
            ce => 'H',
            sr => \N__9020\
        );

    \U712_CHIP_RAM.DMA_CYCLE_1_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__6965\,
            in1 => \N__5957\,
            in2 => \N__5407\,
            in3 => \N__5177\,
            lcout => \RAMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9224\,
            ce => 'H',
            sr => \N__9020\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7916\,
            in2 => \_gnd_net_\,
            in3 => \N__5396\,
            lcout => \U712_CHIP_RAM.DBENn_7_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5787\,
            in1 => \N__7188\,
            in2 => \N__5354\,
            in3 => \N__5273\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIB6KL9_2_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010000"
        )
    port map (
            in0 => \N__5260\,
            in1 => \N__6964\,
            in2 => \N__5207\,
            in3 => \N__5202\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010110011111100"
        )
    port map (
            in0 => \N__5788\,
            in1 => \N__6014\,
            in2 => \N__5864\,
            in3 => \N__5861\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9224\,
            ce => 'H',
            sr => \N__9020\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110110"
        )
    port map (
            in0 => \N__5790\,
            in1 => \N__5542\,
            in2 => \N__5855\,
            in3 => \N__7112\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111100"
        )
    port map (
            in0 => \N__8480\,
            in1 => \N__5828\,
            in2 => \N__5822\,
            in3 => \N__5494\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVS9V_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__5789\,
            in1 => \N__7108\,
            in2 => \_gnd_net_\,
            in3 => \N__5818\,
            lcout => \U712_CHIP_RAM.N_305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__6913\,
            in1 => \N__5791\,
            in2 => \N__7126\,
            in3 => \N__5646\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__7205\,
            in1 => \N__5543\,
            in2 => \N__5513\,
            in3 => \N__7702\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111100"
        )
    port map (
            in0 => \N__8569\,
            in1 => \N__5509\,
            in2 => \N__5498\,
            in3 => \N__5495\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNITDMK_3_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8718\,
            in1 => \N__8568\,
            in2 => \N__8470\,
            in3 => \N__7043\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => \U712_CHIP_RAM.REFRESH_RST_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI9T531_3_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__8696\,
            in1 => \N__8471\,
            in2 => \N__5477\,
            in3 => \N__7044\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__5972\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6024\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0\,
            ltout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_192_i_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100011"
        )
    port map (
            in0 => \N__8858\,
            in1 => \N__5914\,
            in2 => \N__6113\,
            in3 => \N__5870\,
            lcout => \N_192_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_194_i_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__5915\,
            in1 => \N__6089\,
            in2 => \N__8900\,
            in3 => \N__6275\,
            lcout => \N_194_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__6065\,
            in1 => \N__6304\,
            in2 => \_gnd_net_\,
            in3 => \N__8150\,
            lcout => \U712_BYTE_ENABLE.N_404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_0_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6025\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5973\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0\,
            ltout => \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_196_i_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__5912\,
            in1 => \N__6179\,
            in2 => \N__5936\,
            in3 => \N__8853\,
            lcout => \N_196_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__8148\,
            in1 => \N__6265\,
            in2 => \N__6305\,
            in3 => \N__6232\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_198_i_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__5913\,
            in1 => \N__5897\,
            in2 => \N__5891\,
            in3 => \N__8893\,
            lcout => \N_198_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_0_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__8149\,
            in1 => \N__6233\,
            in2 => \_gnd_net_\,
            in3 => \N__6266\,
            lcout => \U712_BYTE_ENABLE.N_405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__6406\,
            in1 => \N__6389\,
            in2 => \_gnd_net_\,
            in3 => \N__6372\,
            lcout => \U712_REG_SM.N_309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__6124\,
            in1 => \N__6603\,
            in2 => \N__6647\,
            in3 => \N__6551\,
            lcout => \U712_REG_SM.N_282\,
            ltout => \U712_REG_SM.N_282_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6578\,
            in2 => \N__6326\,
            in3 => \N__6533\,
            lcout => \U712_REG_SM.N_306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__6300\,
            in1 => \N__6264\,
            in2 => \N__8168\,
            in3 => \N__6231\,
            lcout => \U712_BYTE_ENABLE.N_407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6263\,
            in1 => \N__6230\,
            in2 => \_gnd_net_\,
            in3 => \N__8151\,
            lcout => \U712_BYTE_ENABLE.N_409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_0_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6173\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9238\,
            ce => 'H',
            sr => \N__8993\
        );

    \U712_REG_SM.C3_SYNC_0_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6140\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9238\,
            ce => 'H',
            sr => \N__8993\
        );

    \U712_REG_SM.C1_SYNC_2_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6608\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9238\,
            ce => 'H',
            sr => \N__8993\
        );

    \U712_REG_SM.C1_SYNC_1_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6646\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9238\,
            ce => 'H',
            sr => \N__8993\
        );

    \U712_REG_SM.C3_SYNC_2_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6530\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9238\,
            ce => 'H',
            sr => \N__8993\
        );

    \U712_REG_SM.C3_SYNC_1_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6554\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9241\,
            ce => 'H',
            sr => \N__8991\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__6416\,
            in1 => \_gnd_net_\,
            in2 => \N__8639\,
            in3 => \N__8759\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9203\,
            ce => \N__7964\,
            sr => \N__9036\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011010001"
        )
    port map (
            in0 => \N__8518\,
            in1 => \N__8620\,
            in2 => \N__6659\,
            in3 => \N__8758\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9203\,
            ce => \N__7964\,
            sr => \N__9036\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8757\,
            in1 => \N__8519\,
            in2 => \N__8638\,
            in3 => \N__7061\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9203\,
            ce => \N__7964\,
            sr => \N__9036\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__7325\,
            in1 => \N__8092\,
            in2 => \N__7421\,
            in3 => \N__8520\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8093\,
            in1 => \N__6458\,
            in2 => \N__6440\,
            in3 => \N__6437\,
            lcout => \U712_CHIP_RAM.N_317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111110101"
        )
    port map (
            in0 => \N__7235\,
            in1 => \N__7592\,
            in2 => \N__8146\,
            in3 => \N__8503\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8106\,
            in1 => \N__6857\,
            in2 => \N__6839\,
            in3 => \N__6836\,
            lcout => \U712_CHIP_RAM.N_320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7622\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9207\,
            ce => \N__7837\,
            sr => \N__9027\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__7241\,
            in1 => \N__8502\,
            in2 => \N__8147\,
            in3 => \N__7538\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8107\,
            in1 => \N__6809\,
            in2 => \N__6791\,
            in3 => \N__6788\,
            lcout => \U712_CHIP_RAM.N_321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__8496\,
            in1 => \N__7229\,
            in2 => \N__8133\,
            in3 => \N__9257\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__6767\,
            in1 => \N__6746\,
            in2 => \N__6725\,
            in3 => \N__8080\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__8753\,
            in1 => \_gnd_net_\,
            in2 => \N__6722\,
            in3 => \N__8619\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9211\,
            ce => \N__7951\,
            sr => \N__9021\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7223\,
            in1 => \N__8076\,
            in2 => \N__8514\,
            in3 => \N__7499\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__6701\,
            in1 => \N__6680\,
            in2 => \N__6662\,
            in3 => \N__8099\,
            lcout => \U712_CHIP_RAM.N_316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__7125\,
            in1 => \N__7217\,
            in2 => \_gnd_net_\,
            in3 => \N__7204\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9216\,
            ce => 'H',
            sr => \N__9013\
        );

    \U712_CHIP_RAM.CRCSn_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7060\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9216\,
            ce => 'H',
            sr => \N__9013\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__6912\,
            in1 => \N__7004\,
            in2 => \N__6989\,
            in3 => \N__6977\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9225\,
            ce => 'H',
            sr => \N__9007\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIV62J1_3_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9082\,
            in2 => \_gnd_net_\,
            in3 => \N__6893\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__7363\,
            in1 => \N__7743\,
            in2 => \N__7346\,
            in3 => \N__7795\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_0_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7393\,
            in2 => \N__6887\,
            in3 => \N__6865\,
            lcout => \U712_CHIP_RAM.REFRESHZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9230\,
            ce => 'H',
            sr => \N__8999\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7794\,
            in1 => \N__7341\,
            in2 => \_gnd_net_\,
            in3 => \N__7362\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH9lt7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_1_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__6866\,
            in1 => \N__6884\,
            in2 => \N__6878\,
            in3 => \N__7744\,
            lcout => \U712_CHIP_RAM.REFRESHZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9230\,
            ce => 'H',
            sr => \N__8999\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_RNILI9L_5_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7762\,
            in2 => \_gnd_net_\,
            in3 => \N__7777\,
            lcout => \U712_CHIP_RAM.REFRESH9lto7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7489\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9202\,
            ce => \N__7833\,
            sr => \N__9023\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__8627\,
            in1 => \_gnd_net_\,
            in2 => \N__8767\,
            in3 => \N__7319\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9205\,
            ce => \N__7965\,
            sr => \N__9018\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100000001"
        )
    port map (
            in0 => \N__8760\,
            in1 => \N__8506\,
            in2 => \N__8640\,
            in3 => \N__7292\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9205\,
            ce => \N__7965\,
            sr => \N__9018\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__7271\,
            in1 => \N__8204\,
            in2 => \N__7574\,
            in3 => \N__8136\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9205\,
            ce => \N__7965\,
            sr => \N__9018\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8309\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9206\,
            ce => \N__7832\,
            sr => \N__9012\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7564\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9206\,
            ce => \N__7832\,
            sr => \N__9012\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7529\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9206\,
            ce => \N__7832\,
            sr => \N__9012\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7453\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9206\,
            ce => \N__7832\,
            sr => \N__9012\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7525\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9209\,
            ce => \N__9116\,
            sr => \N__9003\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7493\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9209\,
            ce => \N__9116\,
            sr => \N__9003\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7457\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9209\,
            ce => \N__9116\,
            sr => \N__9003\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__9080\,
            in1 => \N__8779\,
            in2 => \_gnd_net_\,
            in3 => \N__8802\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7382\,
            in2 => \_gnd_net_\,
            in3 => \N__7376\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__7721\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7373\,
            in2 => \_gnd_net_\,
            in3 => \N__7367\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__7721\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7364\,
            in2 => \_gnd_net_\,
            in3 => \N__7349\,
            lcout => \U712_CHIP_RAM.REFRESH9lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__7721\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7345\,
            in2 => \_gnd_net_\,
            in3 => \N__7328\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__7721\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7796\,
            in2 => \_gnd_net_\,
            in3 => \N__7781\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__7721\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7778\,
            in2 => \_gnd_net_\,
            in3 => \N__7766\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__7721\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7763\,
            in2 => \_gnd_net_\,
            in3 => \N__7751\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__7721\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7745\,
            in2 => \_gnd_net_\,
            in3 => \N__7748\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__7721\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7685\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7618\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9208\,
            ce => \N__9108\,
            sr => \N__9028\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7907\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9208\,
            ce => \N__9108\,
            sr => \N__9028\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7871\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9208\,
            ce => \N__9108\,
            sr => \N__9028\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7565\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9208\,
            ce => \N__9108\,
            sr => \N__9028\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__7844\,
            in1 => \N__8505\,
            in2 => \N__8173\,
            in3 => \N__8273\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__8166\,
            in1 => \N__8267\,
            in2 => \N__8249\,
            in3 => \N__8246\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__8615\,
            in1 => \_gnd_net_\,
            in2 => \N__8228\,
            in3 => \N__8754\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9212\,
            ce => \N__7966\,
            sr => \N__9022\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__8504\,
            in1 => \N__8749\,
            in2 => \_gnd_net_\,
            in3 => \N__8614\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_8\,
            ltout => \U712_CHIP_RAM.CMA_5_i_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__8198\,
            in1 => \N__8377\,
            in2 => \N__8177\,
            in3 => \N__8167\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9212\,
            ce => \N__7966\,
            sr => \N__9022\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9295\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9217\,
            ce => \N__7838\,
            sr => \N__9014\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7906\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9217\,
            ce => \N__7838\,
            sr => \N__9014\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7867\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9217\,
            ce => \N__7838\,
            sr => \N__9014\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8892\,
            in2 => \_gnd_net_\,
            in3 => \N__8857\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9226\,
            ce => 'H',
            sr => \N__9008\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8806\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9226\,
            ce => 'H',
            sr => \N__9008\
        );

    \U712_CHIP_RAM.RASn_LC_14_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8768\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9204\,
            ce => 'H',
            sr => \N__9050\
        );

    \U712_CHIP_RAM.WEn_LC_14_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8642\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9204\,
            ce => 'H',
            sr => \N__9050\
        );

    \U712_CHIP_RAM.CASn_LC_14_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8522\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9204\,
            ce => 'H',
            sr => \N__9050\
        );

    \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_14_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__9085\,
            in1 => \N__8326\,
            in2 => \_gnd_net_\,
            in3 => \N__8315\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8378\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8342\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9213\,
            ce => 'H',
            sr => \N__9032\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8327\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9213\,
            ce => 'H',
            sr => \N__9032\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8308\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9218\,
            ce => \N__9112\,
            sr => \N__9029\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9296\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9218\,
            ce => \N__9112\,
            sr => \N__9029\
        );
end \INTERFACE\;

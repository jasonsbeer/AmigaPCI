-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 7 2025 17:55:14

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    DRA : in std_logic_vector(8 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RAMENn : out std_logic;
    RASn : out std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__10415\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_OUT_i_i\ : std_logic;
signal \CLK40_OUT_i_i\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_GOZ0\ : std_logic;
signal \U712_REG_SM.UDS_OUT_2_0_a2_0_a3_0\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.LDS_OUT_2_0_a2_0_a3_0\ : std_logic;
signal \U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1\ : std_logic;
signal \N_944_i\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_cascade_\ : std_logic;
signal \N_41_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_273\ : std_logic;
signal \N_43_i\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_275_cascade_\ : std_logic;
signal \N_42_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_271_cascade_\ : std_logic;
signal \N_44_i\ : std_logic;
signal \A_c_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \U712_BYTE_ENABLE.N_277\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_270\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_266_cascade_\ : std_logic;
signal \U712_REG_SM.N_215\ : std_logic;
signal \U712_REG_SM.N_215_cascade_\ : std_logic;
signal \U712_REG_SM.N_200_cascade_\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \U712_REG_SM.N_200\ : std_logic;
signal \U712_REG_SM.N_219\ : std_logic;
signal \U712_REG_SM.N_325_cascade_\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_198\ : std_logic;
signal \U712_REG_SM.N_212\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_198_cascade_\ : std_logic;
signal \U712_REG_SM.DS_EN_RNOZ0Z_0_cascade_\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.LDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_LDSn_i\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.N_325\ : std_logic;
signal \U712_REG_SM.N_201\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_RNOZ0Z_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_265\ : std_logic;
signal \U712_REG_SM.N_183\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_1\ : std_logic;
signal \U712_CHIP_RAM.DBR_SYNCZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_177_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_197\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_307_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_cascade_\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_0\ : std_logic;
signal \U712_REG_SM.DS_ENZ0\ : std_logic;
signal \U712_REG_SM.UDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_UDSn_i\ : std_logic;
signal \RnW_c\ : std_logic;
signal \DRDDIR_i_m4_i_m2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_209\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.N_323_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a2_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a3_3_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_242_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_188_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_306\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_238\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_323\ : std_logic;
signal \U712_CHIP_RAM.N_240\ : std_logic;
signal \U712_CHIP_RAM.N_10_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER16_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_328\ : std_logic;
signal \U712_CHIP_RAM.N_307\ : std_logic;
signal \U712_CHIP_RAM.N_328_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_177\ : std_logic;
signal \U712_CHIP_RAM.N_251_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_cascade_\ : std_logic;
signal \bfn_10_14_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA30_0_i_cascade_\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_10\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_66_0_i_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNI9MVM2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_222\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_9_0_cascade_\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_3_0\ : std_logic;
signal \U712_CHIP_RAM.N_305_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_221\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\ : std_logic;
signal \U712_CHIP_RAM.N_305\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_10\ : std_logic;
signal \U712_CHIP_RAM.N_260\ : std_logic;
signal \U712_CYCLE_TERM.N_214_i_0_en_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_3\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \A_c_19\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_316_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_3_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_180\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a3_2_1_0\ : std_logic;
signal \U712_CHIP_RAM.N_254_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_0\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.N_187\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_5\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a3_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.N_96\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER16\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_0_a3_0\ : std_logic;
signal \U712_CYCLE_TERM.N_214_i_0_en\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_312\ : std_logic;
signal \U712_CHIP_RAM.N_243\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \CLK40_OUT_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \CASn_c\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA30_0_i_0\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_8C_net\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(8 downto 0);
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    LDSn <= \LDSn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_OUT_i\,
            REFERENCECLK => \N__3691\,
            RESETB => \N__6424\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_OUT\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10415\,
            DIN => \N__10414\,
            DOUT => \N__10413\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10415\,
            PADOUT => \N__10414\,
            PADIN => \N__10413\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5890\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10406\,
            DIN => \N__10405\,
            DOUT => \N__10404\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10406\,
            PADOUT => \N__10405\,
            PADIN => \N__10404\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10397\,
            DIN => \N__10396\,
            DOUT => \N__10395\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10397\,
            PADOUT => \N__10396\,
            PADIN => \N__10395\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8977\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10388\,
            DIN => \N__10387\,
            DOUT => \N__10386\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10388\,
            PADOUT => \N__10387\,
            PADIN => \N__10386\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4927\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10379\,
            DIN => \N__10378\,
            DOUT => \N__10377\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10379\,
            PADOUT => \N__10378\,
            PADIN => \N__10377\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10370\,
            DIN => \N__10369\,
            DOUT => \N__10368\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10370\,
            PADOUT => \N__10369\,
            PADIN => \N__10368\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10361\,
            DIN => \N__10360\,
            DOUT => \N__10359\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10361\,
            PADOUT => \N__10360\,
            PADIN => \N__10359\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10352\,
            DIN => \N__10351\,
            DOUT => \N__10350\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10352\,
            PADOUT => \N__10351\,
            PADIN => \N__10350\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10343\,
            DIN => \N__10342\,
            DOUT => \N__10341\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10343\,
            PADOUT => \N__10342\,
            PADIN => \N__10341\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10334\,
            DIN => \N__10333\,
            DOUT => \N__10332\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10334\,
            PADOUT => \N__10333\,
            PADIN => \N__10332\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6553\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10325\,
            DIN => \N__10324\,
            DOUT => \N__10323\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10325\,
            PADOUT => \N__10324\,
            PADIN => \N__10323\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7759\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10316\,
            DIN => \N__10315\,
            DOUT => \N__10314\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10316\,
            PADOUT => \N__10315\,
            PADIN => \N__10314\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10307\,
            DIN => \N__10306\,
            DOUT => \N__10305\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10307\,
            PADOUT => \N__10306\,
            PADIN => \N__10305\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10298\,
            DIN => \N__10297\,
            DOUT => \N__10296\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10298\,
            PADOUT => \N__10297\,
            PADIN => \N__10296\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3907\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10289\,
            DIN => \N__10288\,
            DOUT => \N__10287\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10289\,
            PADOUT => \N__10288\,
            PADIN => \N__10287\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10280\,
            DIN => \N__10279\,
            DOUT => \N__10278\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10280\,
            PADOUT => \N__10279\,
            PADIN => \N__10278\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10271\,
            DIN => \N__10270\,
            DOUT => \N__10269\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10271\,
            PADOUT => \N__10270\,
            PADIN => \N__10269\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7627\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10262\,
            DIN => \N__10261\,
            DOUT => \N__10260\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10262\,
            PADOUT => \N__10261\,
            PADIN => \N__10260\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10253\,
            DIN => \N__10252\,
            DOUT => \N__10251\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10253\,
            PADOUT => \N__10252\,
            PADIN => \N__10251\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6409\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10244\,
            DIN => \N__10243\,
            DOUT => \N__10242\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10244\,
            PADOUT => \N__10243\,
            PADIN => \N__10242\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10235\,
            DIN => \N__10234\,
            DOUT => \N__10233\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10235\,
            PADOUT => \N__10234\,
            PADIN => \N__10233\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10226\,
            DIN => \N__10225\,
            DOUT => \N__10224\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10226\,
            PADOUT => \N__10225\,
            PADIN => \N__10224\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10217\,
            DIN => \N__10216\,
            DOUT => \N__10215\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10217\,
            PADOUT => \N__10216\,
            PADIN => \N__10215\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10208\,
            DIN => \N__10207\,
            DOUT => \N__10206\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10208\,
            PADOUT => \N__10207\,
            PADIN => \N__10206\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10199\,
            DIN => \N__10198\,
            DOUT => \N__10197\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10199\,
            PADOUT => \N__10198\,
            PADIN => \N__10197\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10190\,
            DIN => \N__10189\,
            DOUT => \N__10188\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10190\,
            PADOUT => \N__10189\,
            PADIN => \N__10188\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10181\,
            DIN => \N__10180\,
            DOUT => \N__10179\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10181\,
            PADOUT => \N__10180\,
            PADIN => \N__10179\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10172\,
            DIN => \N__10171\,
            DOUT => \N__10170\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10172\,
            PADOUT => \N__10171\,
            PADIN => \N__10170\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10163\,
            DIN => \N__10162\,
            DOUT => \N__10161\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10163\,
            PADOUT => \N__10162\,
            PADIN => \N__10161\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6271\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10154\,
            DIN => \N__10153\,
            DOUT => \N__10152\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10154\,
            PADOUT => \N__10153\,
            PADIN => \N__10152\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10145\,
            DIN => \N__10144\,
            DOUT => \N__10143\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10145\,
            PADOUT => \N__10144\,
            PADIN => \N__10143\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10136\,
            DIN => \N__10135\,
            DOUT => \N__10134\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10136\,
            PADOUT => \N__10135\,
            PADIN => \N__10134\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10127\,
            DIN => \N__10126\,
            DOUT => \N__10125\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10127\,
            PADOUT => \N__10126\,
            PADIN => \N__10125\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10118\,
            DIN => \N__10117\,
            DOUT => \N__10116\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10118\,
            PADOUT => \N__10117\,
            PADIN => \N__10116\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3724\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10109\,
            DIN => \N__10108\,
            DOUT => \N__10107\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10109\,
            PADOUT => \N__10108\,
            PADIN => \N__10107\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4363\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10100\,
            DIN => \N__10099\,
            DOUT => \N__10098\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10100\,
            PADOUT => \N__10099\,
            PADIN => \N__10098\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10091\,
            DIN => \N__10090\,
            DOUT => \N__10089\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10091\,
            PADOUT => \N__10090\,
            PADIN => \N__10089\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8989\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10082\,
            DIN => \N__10081\,
            DOUT => \N__10080\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10082\,
            PADOUT => \N__10081\,
            PADIN => \N__10080\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10073\,
            DIN => \N__10072\,
            DOUT => \N__10071\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10073\,
            PADOUT => \N__10072\,
            PADIN => \N__10071\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10064\,
            DIN => \N__10063\,
            DOUT => \N__10062\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10064\,
            PADOUT => \N__10063\,
            PADIN => \N__10062\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3739\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10055\,
            DIN => \N__10054\,
            DOUT => \N__10053\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10055\,
            PADOUT => \N__10054\,
            PADIN => \N__10053\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10046\,
            DIN => \N__10045\,
            DOUT => \N__10044\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10046\,
            PADOUT => \N__10045\,
            PADIN => \N__10044\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3982\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10037\,
            DIN => \N__10036\,
            DOUT => \N__10035\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10037\,
            PADOUT => \N__10036\,
            PADIN => \N__10035\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5647\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10028\,
            DIN => \N__10027\,
            DOUT => \N__10026\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10028\,
            PADOUT => \N__10027\,
            PADIN => \N__10026\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10019\,
            DIN => \N__10018\,
            DOUT => \N__10017\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10019\,
            PADOUT => \N__10018\,
            PADIN => \N__10017\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__10010\,
            DIN => \N__10009\,
            DOUT => \N__10008\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10010\,
            PADOUT => \N__10009\,
            PADIN => \N__10008\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10001\,
            DIN => \N__10000\,
            DOUT => \N__9999\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10001\,
            PADOUT => \N__10000\,
            PADIN => \N__9999\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6151\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9992\,
            DIN => \N__9991\,
            DOUT => \N__9990\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9992\,
            PADOUT => \N__9991\,
            PADIN => \N__9990\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9983\,
            DIN => \N__9982\,
            DOUT => \N__9981\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9983\,
            PADOUT => \N__9982\,
            PADIN => \N__9981\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8809\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9974\,
            DIN => \N__9973\,
            DOUT => \N__9972\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9974\,
            PADOUT => \N__9973\,
            PADIN => \N__9972\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7654\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9965\,
            DIN => \N__9964\,
            DOUT => \N__9963\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9965\,
            PADOUT => \N__9964\,
            PADIN => \N__9963\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3892\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9956\,
            DIN => \N__9955\,
            DOUT => \N__9954\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9956\,
            PADOUT => \N__9955\,
            PADIN => \N__9954\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6331\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9947\,
            DIN => \N__9946\,
            DOUT => \N__9945\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9947\,
            PADOUT => \N__9946\,
            PADIN => \N__9945\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3978\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9938\,
            DIN => \N__9937\,
            DOUT => \N__9936\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9938\,
            PADOUT => \N__9937\,
            PADIN => \N__9936\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9929\,
            DIN => \N__9928\,
            DOUT => \N__9927\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9929\,
            PADOUT => \N__9928\,
            PADIN => \N__9927\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9920\,
            DIN => \N__9919\,
            DOUT => \N__9918\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9920\,
            PADOUT => \N__9919\,
            PADIN => \N__9918\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3844\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9911\,
            DIN => \N__9910\,
            DOUT => \N__9909\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9911\,
            PADOUT => \N__9910\,
            PADIN => \N__9909\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6388\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9902\,
            DIN => \N__9901\,
            DOUT => \N__9900\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9902\,
            PADOUT => \N__9901\,
            PADIN => \N__9900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5230\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9893\,
            DIN => \N__9892\,
            DOUT => \N__9891\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9893\,
            PADOUT => \N__9892\,
            PADIN => \N__9891\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3871\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9884\,
            DIN => \N__9883\,
            DOUT => \N__9882\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9884\,
            PADOUT => \N__9883\,
            PADIN => \N__9882\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9875\,
            DIN => \N__9874\,
            DOUT => \N__9873\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9875\,
            PADOUT => \N__9874\,
            PADIN => \N__9873\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9866\,
            DIN => \N__9865\,
            DOUT => \N__9864\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9866\,
            PADOUT => \N__9865\,
            PADIN => \N__9864\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9857\,
            DIN => \N__9856\,
            DOUT => \N__9855\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9857\,
            PADOUT => \N__9856\,
            PADIN => \N__9855\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9848\,
            DIN => \N__9847\,
            DOUT => \N__9846\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9848\,
            PADOUT => \N__9847\,
            PADIN => \N__9846\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6463\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9839\,
            DIN => \N__9838\,
            DOUT => \N__9837\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9839\,
            PADOUT => \N__9838\,
            PADIN => \N__9837\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9830\,
            DIN => \N__9829\,
            DOUT => \N__9828\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9830\,
            PADOUT => \N__9829\,
            PADIN => \N__9828\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4165\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9821\,
            DIN => \N__9820\,
            DOUT => \N__9819\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9821\,
            PADOUT => \N__9820\,
            PADIN => \N__9819\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3928\,
            DIN0 => OPEN,
            DOUT0 => \N__8014\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9812\,
            DIN => \N__9811\,
            DOUT => \N__9810\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9812\,
            PADOUT => \N__9811\,
            PADIN => \N__9810\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5659\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9803\,
            DIN => \N__9802\,
            DOUT => \N__9801\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9803\,
            PADOUT => \N__9802\,
            PADIN => \N__9801\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9794\,
            DIN => \N__9793\,
            DOUT => \N__9792\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9794\,
            PADOUT => \N__9793\,
            PADIN => \N__9792\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9785\,
            DIN => \N__9784\,
            DOUT => \N__9783\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9785\,
            PADOUT => \N__9784\,
            PADIN => \N__9783\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6295\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9776\,
            DIN => \N__9775\,
            DOUT => \N__9774\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9776\,
            PADOUT => \N__9775\,
            PADIN => \N__9774\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9767\,
            DIN => \N__9766\,
            DOUT => \N__9765\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9767\,
            PADOUT => \N__9766\,
            PADIN => \N__9765\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9758\,
            DIN => \N__9757\,
            DOUT => \N__9756\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9758\,
            PADOUT => \N__9757\,
            PADIN => \N__9756\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9749\,
            DIN => \N__9748\,
            DOUT => \N__9747\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9749\,
            PADOUT => \N__9748\,
            PADIN => \N__9747\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9740\,
            DIN => \N__9739\,
            DOUT => \N__9738\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9740\,
            PADOUT => \N__9739\,
            PADIN => \N__9738\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6796\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9731\,
            DIN => \N__9730\,
            DOUT => \N__9729\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9731\,
            PADOUT => \N__9730\,
            PADIN => \N__9729\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5002\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9722\,
            DIN => \N__9721\,
            DOUT => \N__9720\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9722\,
            PADOUT => \N__9721\,
            PADIN => \N__9720\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6046\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9713\,
            DIN => \N__9712\,
            DOUT => \N__9711\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9713\,
            PADOUT => \N__9712\,
            PADIN => \N__9711\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2323\ : CEMux
    port map (
            O => \N__9694\,
            I => \N__9688\
        );

    \I__2322\ : CEMux
    port map (
            O => \N__9693\,
            I => \N__9685\
        );

    \I__2321\ : CEMux
    port map (
            O => \N__9692\,
            I => \N__9682\
        );

    \I__2320\ : CEMux
    port map (
            O => \N__9691\,
            I => \N__9679\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__9688\,
            I => \N__9675\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__9685\,
            I => \N__9672\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__9682\,
            I => \N__9669\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__9679\,
            I => \N__9664\
        );

    \I__2315\ : CEMux
    port map (
            O => \N__9678\,
            I => \N__9661\
        );

    \I__2314\ : Span4Mux_v
    port map (
            O => \N__9675\,
            I => \N__9658\
        );

    \I__2313\ : Span4Mux_h
    port map (
            O => \N__9672\,
            I => \N__9653\
        );

    \I__2312\ : Span4Mux_h
    port map (
            O => \N__9669\,
            I => \N__9653\
        );

    \I__2311\ : CEMux
    port map (
            O => \N__9668\,
            I => \N__9650\
        );

    \I__2310\ : CEMux
    port map (
            O => \N__9667\,
            I => \N__9647\
        );

    \I__2309\ : Sp12to4
    port map (
            O => \N__9664\,
            I => \N__9642\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__9661\,
            I => \N__9642\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__9658\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__9653\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__9650\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__9647\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__2303\ : Odrv12
    port map (
            O => \N__9642\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__2302\ : InMux
    port map (
            O => \N__9631\,
            I => \N__9627\
        );

    \I__2301\ : InMux
    port map (
            O => \N__9630\,
            I => \N__9624\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__9627\,
            I => \N__9621\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__9624\,
            I => \N__9618\
        );

    \I__2298\ : Span4Mux_h
    port map (
            O => \N__9621\,
            I => \N__9615\
        );

    \I__2297\ : Span4Mux_v
    port map (
            O => \N__9618\,
            I => \N__9612\
        );

    \I__2296\ : Sp12to4
    port map (
            O => \N__9615\,
            I => \N__9609\
        );

    \I__2295\ : Span4Mux_v
    port map (
            O => \N__9612\,
            I => \N__9606\
        );

    \I__2294\ : Span12Mux_v
    port map (
            O => \N__9609\,
            I => \N__9601\
        );

    \I__2293\ : Sp12to4
    port map (
            O => \N__9606\,
            I => \N__9601\
        );

    \I__2292\ : Odrv12
    port map (
            O => \N__9601\,
            I => \DRA_c_4\
        );

    \I__2291\ : InMux
    port map (
            O => \N__9598\,
            I => \N__9595\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__9595\,
            I => \N__9592\
        );

    \I__2289\ : Odrv12
    port map (
            O => \N__9592\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2288\ : CEMux
    port map (
            O => \N__9589\,
            I => \N__9582\
        );

    \I__2287\ : CEMux
    port map (
            O => \N__9588\,
            I => \N__9579\
        );

    \I__2286\ : CEMux
    port map (
            O => \N__9587\,
            I => \N__9575\
        );

    \I__2285\ : CEMux
    port map (
            O => \N__9586\,
            I => \N__9572\
        );

    \I__2284\ : CEMux
    port map (
            O => \N__9585\,
            I => \N__9569\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__9582\,
            I => \N__9566\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__9579\,
            I => \N__9563\
        );

    \I__2281\ : CEMux
    port map (
            O => \N__9578\,
            I => \N__9560\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__9575\,
            I => \N__9557\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__9572\,
            I => \N__9554\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__9569\,
            I => \N__9551\
        );

    \I__2277\ : Span4Mux_h
    port map (
            O => \N__9566\,
            I => \N__9544\
        );

    \I__2276\ : Span4Mux_v
    port map (
            O => \N__9563\,
            I => \N__9544\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__9560\,
            I => \N__9544\
        );

    \I__2274\ : Span4Mux_h
    port map (
            O => \N__9557\,
            I => \N__9541\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__9554\,
            I => \N__9536\
        );

    \I__2272\ : Span4Mux_h
    port map (
            O => \N__9551\,
            I => \N__9536\
        );

    \I__2271\ : Sp12to4
    port map (
            O => \N__9544\,
            I => \N__9533\
        );

    \I__2270\ : Odrv4
    port map (
            O => \N__9541\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__9536\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__2268\ : Odrv12
    port map (
            O => \N__9533\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__2267\ : InMux
    port map (
            O => \N__9526\,
            I => \N__9518\
        );

    \I__2266\ : InMux
    port map (
            O => \N__9525\,
            I => \N__9515\
        );

    \I__2265\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9512\
        );

    \I__2264\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9509\
        );

    \I__2263\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9506\
        );

    \I__2262\ : InMux
    port map (
            O => \N__9521\,
            I => \N__9503\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__9518\,
            I => \N__9479\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__9515\,
            I => \N__9464\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__9512\,
            I => \N__9461\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__9509\,
            I => \N__9457\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__9506\,
            I => \N__9454\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__9503\,
            I => \N__9442\
        );

    \I__2255\ : SRMux
    port map (
            O => \N__9502\,
            I => \N__9343\
        );

    \I__2254\ : SRMux
    port map (
            O => \N__9501\,
            I => \N__9343\
        );

    \I__2253\ : SRMux
    port map (
            O => \N__9500\,
            I => \N__9343\
        );

    \I__2252\ : SRMux
    port map (
            O => \N__9499\,
            I => \N__9343\
        );

    \I__2251\ : SRMux
    port map (
            O => \N__9498\,
            I => \N__9343\
        );

    \I__2250\ : SRMux
    port map (
            O => \N__9497\,
            I => \N__9343\
        );

    \I__2249\ : SRMux
    port map (
            O => \N__9496\,
            I => \N__9343\
        );

    \I__2248\ : SRMux
    port map (
            O => \N__9495\,
            I => \N__9343\
        );

    \I__2247\ : SRMux
    port map (
            O => \N__9494\,
            I => \N__9343\
        );

    \I__2246\ : SRMux
    port map (
            O => \N__9493\,
            I => \N__9343\
        );

    \I__2245\ : SRMux
    port map (
            O => \N__9492\,
            I => \N__9343\
        );

    \I__2244\ : SRMux
    port map (
            O => \N__9491\,
            I => \N__9343\
        );

    \I__2243\ : SRMux
    port map (
            O => \N__9490\,
            I => \N__9343\
        );

    \I__2242\ : SRMux
    port map (
            O => \N__9489\,
            I => \N__9343\
        );

    \I__2241\ : SRMux
    port map (
            O => \N__9488\,
            I => \N__9343\
        );

    \I__2240\ : SRMux
    port map (
            O => \N__9487\,
            I => \N__9343\
        );

    \I__2239\ : SRMux
    port map (
            O => \N__9486\,
            I => \N__9343\
        );

    \I__2238\ : SRMux
    port map (
            O => \N__9485\,
            I => \N__9343\
        );

    \I__2237\ : SRMux
    port map (
            O => \N__9484\,
            I => \N__9343\
        );

    \I__2236\ : SRMux
    port map (
            O => \N__9483\,
            I => \N__9343\
        );

    \I__2235\ : SRMux
    port map (
            O => \N__9482\,
            I => \N__9343\
        );

    \I__2234\ : Glb2LocalMux
    port map (
            O => \N__9479\,
            I => \N__9343\
        );

    \I__2233\ : SRMux
    port map (
            O => \N__9478\,
            I => \N__9343\
        );

    \I__2232\ : SRMux
    port map (
            O => \N__9477\,
            I => \N__9343\
        );

    \I__2231\ : SRMux
    port map (
            O => \N__9476\,
            I => \N__9343\
        );

    \I__2230\ : SRMux
    port map (
            O => \N__9475\,
            I => \N__9343\
        );

    \I__2229\ : SRMux
    port map (
            O => \N__9474\,
            I => \N__9343\
        );

    \I__2228\ : SRMux
    port map (
            O => \N__9473\,
            I => \N__9343\
        );

    \I__2227\ : SRMux
    port map (
            O => \N__9472\,
            I => \N__9343\
        );

    \I__2226\ : SRMux
    port map (
            O => \N__9471\,
            I => \N__9343\
        );

    \I__2225\ : SRMux
    port map (
            O => \N__9470\,
            I => \N__9343\
        );

    \I__2224\ : SRMux
    port map (
            O => \N__9469\,
            I => \N__9343\
        );

    \I__2223\ : SRMux
    port map (
            O => \N__9468\,
            I => \N__9343\
        );

    \I__2222\ : SRMux
    port map (
            O => \N__9467\,
            I => \N__9343\
        );

    \I__2221\ : Glb2LocalMux
    port map (
            O => \N__9464\,
            I => \N__9343\
        );

    \I__2220\ : Glb2LocalMux
    port map (
            O => \N__9461\,
            I => \N__9343\
        );

    \I__2219\ : SRMux
    port map (
            O => \N__9460\,
            I => \N__9343\
        );

    \I__2218\ : Glb2LocalMux
    port map (
            O => \N__9457\,
            I => \N__9343\
        );

    \I__2217\ : Glb2LocalMux
    port map (
            O => \N__9454\,
            I => \N__9343\
        );

    \I__2216\ : SRMux
    port map (
            O => \N__9453\,
            I => \N__9343\
        );

    \I__2215\ : SRMux
    port map (
            O => \N__9452\,
            I => \N__9343\
        );

    \I__2214\ : SRMux
    port map (
            O => \N__9451\,
            I => \N__9343\
        );

    \I__2213\ : SRMux
    port map (
            O => \N__9450\,
            I => \N__9343\
        );

    \I__2212\ : SRMux
    port map (
            O => \N__9449\,
            I => \N__9343\
        );

    \I__2211\ : SRMux
    port map (
            O => \N__9448\,
            I => \N__9343\
        );

    \I__2210\ : SRMux
    port map (
            O => \N__9447\,
            I => \N__9343\
        );

    \I__2209\ : SRMux
    port map (
            O => \N__9446\,
            I => \N__9343\
        );

    \I__2208\ : SRMux
    port map (
            O => \N__9445\,
            I => \N__9343\
        );

    \I__2207\ : Glb2LocalMux
    port map (
            O => \N__9442\,
            I => \N__9343\
        );

    \I__2206\ : GlobalMux
    port map (
            O => \N__9343\,
            I => \N__9340\
        );

    \I__2205\ : gio2CtrlBuf
    port map (
            O => \N__9340\,
            I => \RESETn_c_i_g\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__9337\,
            I => \N__9334\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9331\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__9331\,
            I => \N__9328\
        );

    \I__2201\ : Span4Mux_h
    port map (
            O => \N__9328\,
            I => \N__9325\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__9325\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2199\ : InMux
    port map (
            O => \N__9322\,
            I => \N__9319\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__9319\,
            I => \N__9316\
        );

    \I__2197\ : Odrv4
    port map (
            O => \N__9316\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2196\ : InMux
    port map (
            O => \N__9313\,
            I => \N__9310\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__9310\,
            I => \N__9300\
        );

    \I__2194\ : ClkMux
    port map (
            O => \N__9309\,
            I => \N__9283\
        );

    \I__2193\ : ClkMux
    port map (
            O => \N__9308\,
            I => \N__9283\
        );

    \I__2192\ : ClkMux
    port map (
            O => \N__9307\,
            I => \N__9283\
        );

    \I__2191\ : ClkMux
    port map (
            O => \N__9306\,
            I => \N__9283\
        );

    \I__2190\ : ClkMux
    port map (
            O => \N__9305\,
            I => \N__9283\
        );

    \I__2189\ : ClkMux
    port map (
            O => \N__9304\,
            I => \N__9283\
        );

    \I__2188\ : ClkMux
    port map (
            O => \N__9303\,
            I => \N__9283\
        );

    \I__2187\ : Glb2LocalMux
    port map (
            O => \N__9300\,
            I => \N__9283\
        );

    \I__2186\ : GlobalMux
    port map (
            O => \N__9283\,
            I => \N__9280\
        );

    \I__2185\ : gio2CtrlBuf
    port map (
            O => \N__9280\,
            I => \C1_c_g\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9277\,
            I => \N__9272\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9276\,
            I => \N__9269\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9275\,
            I => \N__9266\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9272\,
            I => \N__9263\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__9269\,
            I => \N__9260\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9266\,
            I => \N__9257\
        );

    \I__2178\ : Sp12to4
    port map (
            O => \N__9263\,
            I => \N__9254\
        );

    \I__2177\ : Sp12to4
    port map (
            O => \N__9260\,
            I => \N__9251\
        );

    \I__2176\ : Span4Mux_v
    port map (
            O => \N__9257\,
            I => \N__9248\
        );

    \I__2175\ : Span12Mux_v
    port map (
            O => \N__9254\,
            I => \N__9245\
        );

    \I__2174\ : Span12Mux_h
    port map (
            O => \N__9251\,
            I => \N__9242\
        );

    \I__2173\ : Sp12to4
    port map (
            O => \N__9248\,
            I => \N__9239\
        );

    \I__2172\ : Span12Mux_h
    port map (
            O => \N__9245\,
            I => \N__9234\
        );

    \I__2171\ : Span12Mux_v
    port map (
            O => \N__9242\,
            I => \N__9234\
        );

    \I__2170\ : Span12Mux_h
    port map (
            O => \N__9239\,
            I => \N__9231\
        );

    \I__2169\ : Odrv12
    port map (
            O => \N__9234\,
            I => \DBRn_c\
        );

    \I__2168\ : Odrv12
    port map (
            O => \N__9231\,
            I => \DBRn_c\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9226\,
            I => \N__9223\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__9223\,
            I => \N__9220\
        );

    \I__2165\ : Odrv12
    port map (
            O => \N__9220\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9214\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__9214\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9211\,
            I => \N__9208\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__9208\,
            I => \N__9205\
        );

    \I__2160\ : Span4Mux_v
    port map (
            O => \N__9205\,
            I => \N__9201\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9204\,
            I => \N__9198\
        );

    \I__2158\ : Sp12to4
    port map (
            O => \N__9201\,
            I => \N__9193\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9198\,
            I => \N__9193\
        );

    \I__2156\ : Span12Mux_h
    port map (
            O => \N__9193\,
            I => \N__9190\
        );

    \I__2155\ : Odrv12
    port map (
            O => \N__9190\,
            I => \DRA_c_7\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9187\,
            I => \N__9184\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__9184\,
            I => \N__9181\
        );

    \I__2152\ : Span4Mux_h
    port map (
            O => \N__9181\,
            I => \N__9178\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__9178\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9175\,
            I => \N__9171\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9174\,
            I => \N__9168\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9171\,
            I => \N__9163\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__9168\,
            I => \N__9163\
        );

    \I__2146\ : Span4Mux_h
    port map (
            O => \N__9163\,
            I => \N__9160\
        );

    \I__2145\ : Sp12to4
    port map (
            O => \N__9160\,
            I => \N__9157\
        );

    \I__2144\ : Span12Mux_v
    port map (
            O => \N__9157\,
            I => \N__9154\
        );

    \I__2143\ : Odrv12
    port map (
            O => \N__9154\,
            I => \DRA_c_8\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9151\,
            I => \N__9148\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__9148\,
            I => \N__9145\
        );

    \I__2140\ : Span4Mux_h
    port map (
            O => \N__9145\,
            I => \N__9142\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__9142\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9139\,
            I => \N__9135\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9138\,
            I => \N__9132\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9135\,
            I => \N__9127\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__9132\,
            I => \N__9127\
        );

    \I__2134\ : Span4Mux_v
    port map (
            O => \N__9127\,
            I => \N__9124\
        );

    \I__2133\ : Sp12to4
    port map (
            O => \N__9124\,
            I => \N__9121\
        );

    \I__2132\ : Span12Mux_h
    port map (
            O => \N__9121\,
            I => \N__9118\
        );

    \I__2131\ : Odrv12
    port map (
            O => \N__9118\,
            I => \DRA_c_5\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9115\,
            I => \N__9109\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9114\,
            I => \N__9109\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__9109\,
            I => \N__9106\
        );

    \I__2127\ : Span4Mux_h
    port map (
            O => \N__9106\,
            I => \N__9103\
        );

    \I__2126\ : Odrv4
    port map (
            O => \N__9103\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9100\,
            I => \N__9097\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9097\,
            I => \N__9087\
        );

    \I__2123\ : ClkMux
    port map (
            O => \N__9096\,
            I => \N__9070\
        );

    \I__2122\ : ClkMux
    port map (
            O => \N__9095\,
            I => \N__9070\
        );

    \I__2121\ : ClkMux
    port map (
            O => \N__9094\,
            I => \N__9070\
        );

    \I__2120\ : ClkMux
    port map (
            O => \N__9093\,
            I => \N__9070\
        );

    \I__2119\ : ClkMux
    port map (
            O => \N__9092\,
            I => \N__9070\
        );

    \I__2118\ : ClkMux
    port map (
            O => \N__9091\,
            I => \N__9070\
        );

    \I__2117\ : ClkMux
    port map (
            O => \N__9090\,
            I => \N__9070\
        );

    \I__2116\ : Glb2LocalMux
    port map (
            O => \N__9087\,
            I => \N__9070\
        );

    \I__2115\ : GlobalMux
    port map (
            O => \N__9070\,
            I => \N__9067\
        );

    \I__2114\ : gio2CtrlBuf
    port map (
            O => \N__9067\,
            I => \C3_c_g\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9064\,
            I => \N__9059\
        );

    \I__2112\ : InMux
    port map (
            O => \N__9063\,
            I => \N__9054\
        );

    \I__2111\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9054\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9059\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__9054\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__2108\ : CascadeMux
    port map (
            O => \N__9049\,
            I => \N__9045\
        );

    \I__2107\ : InMux
    port map (
            O => \N__9048\,
            I => \N__9042\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9045\,
            I => \N__9039\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__9042\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9039\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__2103\ : InMux
    port map (
            O => \N__9034\,
            I => \N__9030\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9033\,
            I => \N__9027\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9030\,
            I => \N__9022\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__9027\,
            I => \N__9017\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9026\,
            I => \N__9014\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9025\,
            I => \N__9011\
        );

    \I__2097\ : Span12Mux_v
    port map (
            O => \N__9022\,
            I => \N__9008\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9021\,
            I => \N__9003\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9020\,
            I => \N__9003\
        );

    \I__2094\ : Span4Mux_h
    port map (
            O => \N__9017\,
            I => \N__8996\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__9014\,
            I => \N__8996\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__9011\,
            I => \N__8996\
        );

    \I__2091\ : Odrv12
    port map (
            O => \N__9008\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9003\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__8996\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2088\ : IoInMux
    port map (
            O => \N__8989\,
            I => \N__8986\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__8986\,
            I => \N__8983\
        );

    \I__2086\ : Span12Mux_s8_v
    port map (
            O => \N__8983\,
            I => \N__8980\
        );

    \I__2085\ : Odrv12
    port map (
            O => \N__8980\,
            I => \RASn_c\
        );

    \I__2084\ : IoInMux
    port map (
            O => \N__8977\,
            I => \N__8974\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__8974\,
            I => \N__8971\
        );

    \I__2082\ : IoSpan4Mux
    port map (
            O => \N__8971\,
            I => \N__8968\
        );

    \I__2081\ : Span4Mux_s2_v
    port map (
            O => \N__8968\,
            I => \N__8965\
        );

    \I__2080\ : Sp12to4
    port map (
            O => \N__8965\,
            I => \N__8962\
        );

    \I__2079\ : Span12Mux_s10_v
    port map (
            O => \N__8962\,
            I => \N__8959\
        );

    \I__2078\ : Odrv12
    port map (
            O => \N__8959\,
            I => \CASn_c\
        );

    \I__2077\ : InMux
    port map (
            O => \N__8956\,
            I => \N__8953\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__8953\,
            I => \N__8950\
        );

    \I__2075\ : Span4Mux_v
    port map (
            O => \N__8950\,
            I => \N__8946\
        );

    \I__2074\ : InMux
    port map (
            O => \N__8949\,
            I => \N__8943\
        );

    \I__2073\ : Sp12to4
    port map (
            O => \N__8946\,
            I => \N__8938\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__8943\,
            I => \N__8938\
        );

    \I__2071\ : Span12Mux_h
    port map (
            O => \N__8938\,
            I => \N__8935\
        );

    \I__2070\ : Odrv12
    port map (
            O => \N__8935\,
            I => \DRA_c_6\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__8932\,
            I => \N__8929\
        );

    \I__2068\ : InMux
    port map (
            O => \N__8929\,
            I => \N__8926\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__8926\,
            I => \N__8923\
        );

    \I__2066\ : Odrv4
    port map (
            O => \N__8923\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2065\ : InMux
    port map (
            O => \N__8920\,
            I => \N__8916\
        );

    \I__2064\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8913\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__8916\,
            I => \N__8906\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__8913\,
            I => \N__8903\
        );

    \I__2061\ : InMux
    port map (
            O => \N__8912\,
            I => \N__8900\
        );

    \I__2060\ : InMux
    port map (
            O => \N__8911\,
            I => \N__8897\
        );

    \I__2059\ : InMux
    port map (
            O => \N__8910\,
            I => \N__8894\
        );

    \I__2058\ : InMux
    port map (
            O => \N__8909\,
            I => \N__8891\
        );

    \I__2057\ : Span4Mux_h
    port map (
            O => \N__8906\,
            I => \N__8885\
        );

    \I__2056\ : Span4Mux_v
    port map (
            O => \N__8903\,
            I => \N__8882\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__8900\,
            I => \N__8877\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__8897\,
            I => \N__8877\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__8894\,
            I => \N__8872\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__8891\,
            I => \N__8872\
        );

    \I__2051\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8867\
        );

    \I__2050\ : InMux
    port map (
            O => \N__8889\,
            I => \N__8867\
        );

    \I__2049\ : InMux
    port map (
            O => \N__8888\,
            I => \N__8864\
        );

    \I__2048\ : Odrv4
    port map (
            O => \N__8885\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2047\ : Odrv4
    port map (
            O => \N__8882\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__8877\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__8872\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__8867\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__8864\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__8851\,
            I => \N__8846\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__8850\,
            I => \N__8841\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__8849\,
            I => \N__8837\
        );

    \I__2039\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8834\
        );

    \I__2038\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8831\
        );

    \I__2037\ : InMux
    port map (
            O => \N__8844\,
            I => \N__8826\
        );

    \I__2036\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8826\
        );

    \I__2035\ : InMux
    port map (
            O => \N__8840\,
            I => \N__8821\
        );

    \I__2034\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8821\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__8834\,
            I => \N__8818\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__8831\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__8826\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__8821\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__8818\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2028\ : IoInMux
    port map (
            O => \N__8809\,
            I => \N__8806\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__8806\,
            I => \N__8803\
        );

    \I__2026\ : IoSpan4Mux
    port map (
            O => \N__8803\,
            I => \N__8800\
        );

    \I__2025\ : Sp12to4
    port map (
            O => \N__8800\,
            I => \N__8797\
        );

    \I__2024\ : Span12Mux_s9_h
    port map (
            O => \N__8797\,
            I => \N__8794\
        );

    \I__2023\ : Span12Mux_v
    port map (
            O => \N__8794\,
            I => \N__8791\
        );

    \I__2022\ : Odrv12
    port map (
            O => \N__8791\,
            I => \CMA_c_4\
        );

    \I__2021\ : InMux
    port map (
            O => \N__8788\,
            I => \N__8785\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__8785\,
            I => \N__8755\
        );

    \I__2019\ : ClkMux
    port map (
            O => \N__8784\,
            I => \N__8674\
        );

    \I__2018\ : ClkMux
    port map (
            O => \N__8783\,
            I => \N__8674\
        );

    \I__2017\ : ClkMux
    port map (
            O => \N__8782\,
            I => \N__8674\
        );

    \I__2016\ : ClkMux
    port map (
            O => \N__8781\,
            I => \N__8674\
        );

    \I__2015\ : ClkMux
    port map (
            O => \N__8780\,
            I => \N__8674\
        );

    \I__2014\ : ClkMux
    port map (
            O => \N__8779\,
            I => \N__8674\
        );

    \I__2013\ : ClkMux
    port map (
            O => \N__8778\,
            I => \N__8674\
        );

    \I__2012\ : ClkMux
    port map (
            O => \N__8777\,
            I => \N__8674\
        );

    \I__2011\ : ClkMux
    port map (
            O => \N__8776\,
            I => \N__8674\
        );

    \I__2010\ : ClkMux
    port map (
            O => \N__8775\,
            I => \N__8674\
        );

    \I__2009\ : ClkMux
    port map (
            O => \N__8774\,
            I => \N__8674\
        );

    \I__2008\ : ClkMux
    port map (
            O => \N__8773\,
            I => \N__8674\
        );

    \I__2007\ : ClkMux
    port map (
            O => \N__8772\,
            I => \N__8674\
        );

    \I__2006\ : ClkMux
    port map (
            O => \N__8771\,
            I => \N__8674\
        );

    \I__2005\ : ClkMux
    port map (
            O => \N__8770\,
            I => \N__8674\
        );

    \I__2004\ : ClkMux
    port map (
            O => \N__8769\,
            I => \N__8674\
        );

    \I__2003\ : ClkMux
    port map (
            O => \N__8768\,
            I => \N__8674\
        );

    \I__2002\ : ClkMux
    port map (
            O => \N__8767\,
            I => \N__8674\
        );

    \I__2001\ : ClkMux
    port map (
            O => \N__8766\,
            I => \N__8674\
        );

    \I__2000\ : ClkMux
    port map (
            O => \N__8765\,
            I => \N__8674\
        );

    \I__1999\ : ClkMux
    port map (
            O => \N__8764\,
            I => \N__8674\
        );

    \I__1998\ : ClkMux
    port map (
            O => \N__8763\,
            I => \N__8674\
        );

    \I__1997\ : ClkMux
    port map (
            O => \N__8762\,
            I => \N__8674\
        );

    \I__1996\ : ClkMux
    port map (
            O => \N__8761\,
            I => \N__8674\
        );

    \I__1995\ : ClkMux
    port map (
            O => \N__8760\,
            I => \N__8674\
        );

    \I__1994\ : ClkMux
    port map (
            O => \N__8759\,
            I => \N__8674\
        );

    \I__1993\ : ClkMux
    port map (
            O => \N__8758\,
            I => \N__8674\
        );

    \I__1992\ : Glb2LocalMux
    port map (
            O => \N__8755\,
            I => \N__8674\
        );

    \I__1991\ : ClkMux
    port map (
            O => \N__8754\,
            I => \N__8674\
        );

    \I__1990\ : ClkMux
    port map (
            O => \N__8753\,
            I => \N__8674\
        );

    \I__1989\ : ClkMux
    port map (
            O => \N__8752\,
            I => \N__8674\
        );

    \I__1988\ : ClkMux
    port map (
            O => \N__8751\,
            I => \N__8674\
        );

    \I__1987\ : ClkMux
    port map (
            O => \N__8750\,
            I => \N__8674\
        );

    \I__1986\ : ClkMux
    port map (
            O => \N__8749\,
            I => \N__8674\
        );

    \I__1985\ : ClkMux
    port map (
            O => \N__8748\,
            I => \N__8674\
        );

    \I__1984\ : ClkMux
    port map (
            O => \N__8747\,
            I => \N__8674\
        );

    \I__1983\ : GlobalMux
    port map (
            O => \N__8674\,
            I => \CLK80_OUT\
        );

    \I__1982\ : CEMux
    port map (
            O => \N__8671\,
            I => \N__8665\
        );

    \I__1981\ : CEMux
    port map (
            O => \N__8670\,
            I => \N__8661\
        );

    \I__1980\ : CEMux
    port map (
            O => \N__8669\,
            I => \N__8658\
        );

    \I__1979\ : CEMux
    port map (
            O => \N__8668\,
            I => \N__8655\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__8665\,
            I => \N__8651\
        );

    \I__1977\ : CEMux
    port map (
            O => \N__8664\,
            I => \N__8648\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__8661\,
            I => \N__8645\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__8658\,
            I => \N__8642\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__8655\,
            I => \N__8639\
        );

    \I__1973\ : CEMux
    port map (
            O => \N__8654\,
            I => \N__8636\
        );

    \I__1972\ : Span4Mux_h
    port map (
            O => \N__8651\,
            I => \N__8631\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__8648\,
            I => \N__8631\
        );

    \I__1970\ : Span4Mux_v
    port map (
            O => \N__8645\,
            I => \N__8628\
        );

    \I__1969\ : Span4Mux_v
    port map (
            O => \N__8642\,
            I => \N__8625\
        );

    \I__1968\ : Span4Mux_h
    port map (
            O => \N__8639\,
            I => \N__8620\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__8636\,
            I => \N__8620\
        );

    \I__1966\ : Span4Mux_v
    port map (
            O => \N__8631\,
            I => \N__8617\
        );

    \I__1965\ : Odrv4
    port map (
            O => \N__8628\,
            I => \U712_CHIP_RAM.un1_CMA30_0_i_0\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__8625\,
            I => \U712_CHIP_RAM.un1_CMA30_0_i_0\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__8620\,
            I => \U712_CHIP_RAM.un1_CMA30_0_i_0\
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__8617\,
            I => \U712_CHIP_RAM.un1_CMA30_0_i_0\
        );

    \I__1961\ : InMux
    port map (
            O => \N__8608\,
            I => \N__8605\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__8605\,
            I => \N__8602\
        );

    \I__1959\ : Span4Mux_v
    port map (
            O => \N__8602\,
            I => \N__8599\
        );

    \I__1958\ : Sp12to4
    port map (
            O => \N__8599\,
            I => \N__8596\
        );

    \I__1957\ : Span12Mux_h
    port map (
            O => \N__8596\,
            I => \N__8593\
        );

    \I__1956\ : Odrv12
    port map (
            O => \N__8593\,
            I => \A_c_13\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8587\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__8587\,
            I => \N__8584\
        );

    \I__1953\ : Span4Mux_v
    port map (
            O => \N__8584\,
            I => \N__8581\
        );

    \I__1952\ : Sp12to4
    port map (
            O => \N__8581\,
            I => \N__8578\
        );

    \I__1951\ : Span12Mux_h
    port map (
            O => \N__8578\,
            I => \N__8575\
        );

    \I__1950\ : Odrv12
    port map (
            O => \N__8575\,
            I => \A_c_6\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__8572\,
            I => \N__8566\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__8571\,
            I => \N__8558\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__8570\,
            I => \N__8555\
        );

    \I__1946\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8549\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8566\,
            I => \N__8542\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8565\,
            I => \N__8539\
        );

    \I__1943\ : InMux
    port map (
            O => \N__8564\,
            I => \N__8536\
        );

    \I__1942\ : InMux
    port map (
            O => \N__8563\,
            I => \N__8529\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8529\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8561\,
            I => \N__8529\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8516\
        );

    \I__1938\ : InMux
    port map (
            O => \N__8555\,
            I => \N__8516\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8554\,
            I => \N__8516\
        );

    \I__1936\ : InMux
    port map (
            O => \N__8553\,
            I => \N__8511\
        );

    \I__1935\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8511\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__8549\,
            I => \N__8508\
        );

    \I__1933\ : InMux
    port map (
            O => \N__8548\,
            I => \N__8505\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8547\,
            I => \N__8500\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8546\,
            I => \N__8500\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8545\,
            I => \N__8496\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__8542\,
            I => \N__8487\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__8539\,
            I => \N__8487\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__8536\,
            I => \N__8487\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__8529\,
            I => \N__8487\
        );

    \I__1925\ : InMux
    port map (
            O => \N__8528\,
            I => \N__8484\
        );

    \I__1924\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8473\
        );

    \I__1923\ : InMux
    port map (
            O => \N__8526\,
            I => \N__8473\
        );

    \I__1922\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8473\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8473\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8523\,
            I => \N__8473\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__8516\,
            I => \N__8468\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__8511\,
            I => \N__8468\
        );

    \I__1917\ : Span4Mux_h
    port map (
            O => \N__8508\,
            I => \N__8461\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__8505\,
            I => \N__8461\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__8500\,
            I => \N__8461\
        );

    \I__1914\ : InMux
    port map (
            O => \N__8499\,
            I => \N__8458\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__8496\,
            I => \N__8455\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__8487\,
            I => \N__8452\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__8484\,
            I => \N__8447\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__8473\,
            I => \N__8447\
        );

    \I__1909\ : Span4Mux_h
    port map (
            O => \N__8468\,
            I => \N__8438\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__8461\,
            I => \N__8438\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8458\,
            I => \N__8438\
        );

    \I__1906\ : Span4Mux_h
    port map (
            O => \N__8455\,
            I => \N__8438\
        );

    \I__1905\ : Odrv4
    port map (
            O => \N__8452\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1904\ : Odrv12
    port map (
            O => \N__8447\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__8438\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8431\,
            I => \N__8424\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8424\
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__8429\,
            I => \N__8412\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__8424\,
            I => \N__8409\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8406\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__8422\,
            I => \N__8403\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8397\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8391\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__8419\,
            I => \N__8384\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8418\,
            I => \N__8381\
        );

    \I__1892\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8378\
        );

    \I__1891\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8371\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8415\,
            I => \N__8371\
        );

    \I__1889\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8371\
        );

    \I__1888\ : Span4Mux_v
    port map (
            O => \N__8409\,
            I => \N__8366\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8406\,
            I => \N__8366\
        );

    \I__1886\ : InMux
    port map (
            O => \N__8403\,
            I => \N__8359\
        );

    \I__1885\ : InMux
    port map (
            O => \N__8402\,
            I => \N__8359\
        );

    \I__1884\ : InMux
    port map (
            O => \N__8401\,
            I => \N__8359\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8400\,
            I => \N__8356\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__8397\,
            I => \N__8353\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8396\,
            I => \N__8346\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8395\,
            I => \N__8346\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8394\,
            I => \N__8346\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8391\,
            I => \N__8343\
        );

    \I__1877\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8336\
        );

    \I__1876\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8336\
        );

    \I__1875\ : InMux
    port map (
            O => \N__8388\,
            I => \N__8336\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8331\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8384\,
            I => \N__8331\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8381\,
            I => \N__8327\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8378\,
            I => \N__8318\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8371\,
            I => \N__8318\
        );

    \I__1869\ : Span4Mux_h
    port map (
            O => \N__8366\,
            I => \N__8318\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8359\,
            I => \N__8318\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8356\,
            I => \N__8311\
        );

    \I__1866\ : Span4Mux_v
    port map (
            O => \N__8353\,
            I => \N__8311\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8346\,
            I => \N__8311\
        );

    \I__1864\ : Span4Mux_v
    port map (
            O => \N__8343\,
            I => \N__8304\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__8336\,
            I => \N__8304\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8331\,
            I => \N__8304\
        );

    \I__1861\ : InMux
    port map (
            O => \N__8330\,
            I => \N__8301\
        );

    \I__1860\ : Span4Mux_v
    port map (
            O => \N__8327\,
            I => \N__8296\
        );

    \I__1859\ : Span4Mux_v
    port map (
            O => \N__8318\,
            I => \N__8296\
        );

    \I__1858\ : Span4Mux_h
    port map (
            O => \N__8311\,
            I => \N__8293\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__8304\,
            I => \CPU_CYCLEm\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8301\,
            I => \CPU_CYCLEm\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__8296\,
            I => \CPU_CYCLEm\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__8293\,
            I => \CPU_CYCLEm\
        );

    \I__1853\ : CascadeMux
    port map (
            O => \N__8284\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\
        );

    \I__1852\ : InMux
    port map (
            O => \N__8281\,
            I => \N__8278\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__8278\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1850\ : InMux
    port map (
            O => \N__8275\,
            I => \N__8272\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8272\,
            I => \N__8269\
        );

    \I__1848\ : Span4Mux_v
    port map (
            O => \N__8269\,
            I => \N__8265\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8268\,
            I => \N__8262\
        );

    \I__1846\ : Sp12to4
    port map (
            O => \N__8265\,
            I => \N__8259\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8262\,
            I => \N__8256\
        );

    \I__1844\ : Span12Mux_h
    port map (
            O => \N__8259\,
            I => \N__8253\
        );

    \I__1843\ : Span12Mux_v
    port map (
            O => \N__8256\,
            I => \N__8250\
        );

    \I__1842\ : Span12Mux_v
    port map (
            O => \N__8253\,
            I => \N__8245\
        );

    \I__1841\ : Span12Mux_h
    port map (
            O => \N__8250\,
            I => \N__8245\
        );

    \I__1840\ : Odrv12
    port map (
            O => \N__8245\,
            I => \DRA_c_0\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__8242\,
            I => \N__8239\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8239\,
            I => \N__8236\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__8236\,
            I => \N__8233\
        );

    \I__1836\ : Span4Mux_h
    port map (
            O => \N__8233\,
            I => \N__8230\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__8230\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8227\,
            I => \N__8223\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8226\,
            I => \N__8220\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8223\,
            I => \N__8215\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__8220\,
            I => \N__8215\
        );

    \I__1830\ : Span4Mux_v
    port map (
            O => \N__8215\,
            I => \N__8212\
        );

    \I__1829\ : Span4Mux_v
    port map (
            O => \N__8212\,
            I => \N__8209\
        );

    \I__1828\ : Sp12to4
    port map (
            O => \N__8209\,
            I => \N__8206\
        );

    \I__1827\ : Span12Mux_h
    port map (
            O => \N__8206\,
            I => \N__8203\
        );

    \I__1826\ : Odrv12
    port map (
            O => \N__8203\,
            I => \DRA_c_3\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8197\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__8197\,
            I => \N__8194\
        );

    \I__1823\ : Span4Mux_v
    port map (
            O => \N__8194\,
            I => \N__8191\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__8191\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8188\,
            I => \N__8185\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8185\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8182\,
            I => \N__8179\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__8179\,
            I => \N__8175\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8178\,
            I => \N__8172\
        );

    \I__1816\ : Span4Mux_h
    port map (
            O => \N__8175\,
            I => \N__8167\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__8172\,
            I => \N__8167\
        );

    \I__1814\ : Sp12to4
    port map (
            O => \N__8167\,
            I => \N__8164\
        );

    \I__1813\ : Span12Mux_v
    port map (
            O => \N__8164\,
            I => \N__8161\
        );

    \I__1812\ : Span12Mux_h
    port map (
            O => \N__8161\,
            I => \N__8158\
        );

    \I__1811\ : Odrv12
    port map (
            O => \N__8158\,
            I => \DRA_c_1\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8149\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8154\,
            I => \N__8149\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8149\,
            I => \N__8146\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__8146\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__8143\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0_cascade_\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8140\,
            I => \N__8137\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__8137\,
            I => \N__8131\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8136\,
            I => \N__8128\
        );

    \I__1802\ : InMux
    port map (
            O => \N__8135\,
            I => \N__8125\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8134\,
            I => \N__8122\
        );

    \I__1800\ : Span4Mux_h
    port map (
            O => \N__8131\,
            I => \N__8117\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8128\,
            I => \N__8117\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8125\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8122\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1796\ : Odrv4
    port map (
            O => \N__8117\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8110\,
            I => \N__8107\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__8107\,
            I => \N__8104\
        );

    \I__1793\ : Span4Mux_v
    port map (
            O => \N__8104\,
            I => \N__8100\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8096\
        );

    \I__1791\ : Span4Mux_h
    port map (
            O => \N__8100\,
            I => \N__8093\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8090\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__8096\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1788\ : Odrv4
    port map (
            O => \N__8093\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__8090\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8083\,
            I => \N__8077\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8082\,
            I => \N__8077\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8077\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1783\ : InMux
    port map (
            O => \N__8074\,
            I => \N__8071\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8071\,
            I => \N__8068\
        );

    \I__1781\ : Span4Mux_v
    port map (
            O => \N__8068\,
            I => \N__8065\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__8065\,
            I => \N__8059\
        );

    \I__1779\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8054\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8063\,
            I => \N__8054\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8062\,
            I => \N__8051\
        );

    \I__1776\ : Sp12to4
    port map (
            O => \N__8059\,
            I => \N__8048\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__8054\,
            I => \N__8043\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__8051\,
            I => \N__8043\
        );

    \I__1773\ : Span12Mux_h
    port map (
            O => \N__8048\,
            I => \N__8038\
        );

    \I__1772\ : Span12Mux_v
    port map (
            O => \N__8043\,
            I => \N__8038\
        );

    \I__1771\ : Odrv12
    port map (
            O => \N__8038\,
            I => \CLK40_OUT_i\
        );

    \I__1770\ : CascadeMux
    port map (
            O => \N__8035\,
            I => \N__8032\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8032\,
            I => \N__8026\
        );

    \I__1768\ : InMux
    port map (
            O => \N__8031\,
            I => \N__8019\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8030\,
            I => \N__8019\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8029\,
            I => \N__8019\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__8026\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8019\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1763\ : IoInMux
    port map (
            O => \N__8014\,
            I => \N__8011\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__8011\,
            I => \N__8008\
        );

    \I__1761\ : Span4Mux_s3_h
    port map (
            O => \N__8008\,
            I => \N__8005\
        );

    \I__1760\ : Span4Mux_v
    port map (
            O => \N__8005\,
            I => \N__8002\
        );

    \I__1759\ : Span4Mux_v
    port map (
            O => \N__8002\,
            I => \N__7999\
        );

    \I__1758\ : Sp12to4
    port map (
            O => \N__7999\,
            I => \N__7995\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__7998\,
            I => \N__7992\
        );

    \I__1756\ : Span12Mux_h
    port map (
            O => \N__7995\,
            I => \N__7989\
        );

    \I__1755\ : InMux
    port map (
            O => \N__7992\,
            I => \N__7986\
        );

    \I__1754\ : Odrv12
    port map (
            O => \N__7989\,
            I => \TACK_OUTn\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__7986\,
            I => \TACK_OUTn\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__7981\,
            I => \N__7974\
        );

    \I__1751\ : InMux
    port map (
            O => \N__7980\,
            I => \N__7971\
        );

    \I__1750\ : InMux
    port map (
            O => \N__7979\,
            I => \N__7966\
        );

    \I__1749\ : InMux
    port map (
            O => \N__7978\,
            I => \N__7966\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__7977\,
            I => \N__7962\
        );

    \I__1747\ : InMux
    port map (
            O => \N__7974\,
            I => \N__7955\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__7971\,
            I => \N__7952\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__7966\,
            I => \N__7949\
        );

    \I__1744\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7946\
        );

    \I__1743\ : InMux
    port map (
            O => \N__7962\,
            I => \N__7943\
        );

    \I__1742\ : InMux
    port map (
            O => \N__7961\,
            I => \N__7938\
        );

    \I__1741\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7938\
        );

    \I__1740\ : InMux
    port map (
            O => \N__7959\,
            I => \N__7934\
        );

    \I__1739\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7931\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__7955\,
            I => \N__7928\
        );

    \I__1737\ : Span4Mux_h
    port map (
            O => \N__7952\,
            I => \N__7925\
        );

    \I__1736\ : Span4Mux_h
    port map (
            O => \N__7949\,
            I => \N__7920\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__7946\,
            I => \N__7920\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__7943\,
            I => \N__7915\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__7938\,
            I => \N__7915\
        );

    \I__1732\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7912\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__7934\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__7931\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1729\ : Odrv4
    port map (
            O => \N__7928\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1728\ : Odrv4
    port map (
            O => \N__7925\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__7920\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1726\ : Odrv12
    port map (
            O => \N__7915\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__7912\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__7897\,
            I => \N__7893\
        );

    \I__1723\ : InMux
    port map (
            O => \N__7896\,
            I => \N__7889\
        );

    \I__1722\ : InMux
    port map (
            O => \N__7893\,
            I => \N__7886\
        );

    \I__1721\ : InMux
    port map (
            O => \N__7892\,
            I => \N__7880\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__7889\,
            I => \N__7875\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__7886\,
            I => \N__7875\
        );

    \I__1718\ : InMux
    port map (
            O => \N__7885\,
            I => \N__7872\
        );

    \I__1717\ : InMux
    port map (
            O => \N__7884\,
            I => \N__7867\
        );

    \I__1716\ : InMux
    port map (
            O => \N__7883\,
            I => \N__7867\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__7880\,
            I => \U712_CHIP_RAM.N_312\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__7875\,
            I => \U712_CHIP_RAM.N_312\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__7872\,
            I => \U712_CHIP_RAM.N_312\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__7867\,
            I => \U712_CHIP_RAM.N_312\
        );

    \I__1711\ : InMux
    port map (
            O => \N__7858\,
            I => \N__7855\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__7855\,
            I => \N__7852\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__7852\,
            I => \U712_CHIP_RAM.N_243\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__7849\,
            I => \N__7846\
        );

    \I__1707\ : InMux
    port map (
            O => \N__7846\,
            I => \N__7838\
        );

    \I__1706\ : InMux
    port map (
            O => \N__7845\,
            I => \N__7835\
        );

    \I__1705\ : InMux
    port map (
            O => \N__7844\,
            I => \N__7832\
        );

    \I__1704\ : InMux
    port map (
            O => \N__7843\,
            I => \N__7825\
        );

    \I__1703\ : InMux
    port map (
            O => \N__7842\,
            I => \N__7825\
        );

    \I__1702\ : InMux
    port map (
            O => \N__7841\,
            I => \N__7825\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__7838\,
            I => \N__7812\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__7835\,
            I => \N__7812\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__7832\,
            I => \N__7812\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__7825\,
            I => \N__7812\
        );

    \I__1697\ : InMux
    port map (
            O => \N__7824\,
            I => \N__7809\
        );

    \I__1696\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7806\
        );

    \I__1695\ : InMux
    port map (
            O => \N__7822\,
            I => \N__7803\
        );

    \I__1694\ : InMux
    port map (
            O => \N__7821\,
            I => \N__7800\
        );

    \I__1693\ : Span4Mux_v
    port map (
            O => \N__7812\,
            I => \N__7797\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__7809\,
            I => \N__7788\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__7806\,
            I => \N__7788\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__7803\,
            I => \N__7788\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__7800\,
            I => \N__7788\
        );

    \I__1688\ : Sp12to4
    port map (
            O => \N__7797\,
            I => \N__7785\
        );

    \I__1687\ : Span12Mux_v
    port map (
            O => \N__7788\,
            I => \N__7782\
        );

    \I__1686\ : Span12Mux_h
    port map (
            O => \N__7785\,
            I => \N__7779\
        );

    \I__1685\ : Span12Mux_h
    port map (
            O => \N__7782\,
            I => \N__7776\
        );

    \I__1684\ : Odrv12
    port map (
            O => \N__7779\,
            I => \RESETn_c\
        );

    \I__1683\ : Odrv12
    port map (
            O => \N__7776\,
            I => \RESETn_c\
        );

    \I__1682\ : IoInMux
    port map (
            O => \N__7771\,
            I => \N__7768\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__7768\,
            I => \N__7765\
        );

    \I__1680\ : Span12Mux_s1_v
    port map (
            O => \N__7765\,
            I => \N__7762\
        );

    \I__1679\ : Odrv12
    port map (
            O => \N__7762\,
            I => \RESETn_c_i\
        );

    \I__1678\ : IoInMux
    port map (
            O => \N__7759\,
            I => \N__7756\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__7756\,
            I => \N__7753\
        );

    \I__1676\ : IoSpan4Mux
    port map (
            O => \N__7753\,
            I => \N__7750\
        );

    \I__1675\ : IoSpan4Mux
    port map (
            O => \N__7750\,
            I => \N__7747\
        );

    \I__1674\ : Span4Mux_s2_v
    port map (
            O => \N__7747\,
            I => \N__7743\
        );

    \I__1673\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7740\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__7743\,
            I => \N__7734\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__7740\,
            I => \N__7734\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__7739\,
            I => \N__7729\
        );

    \I__1669\ : Span4Mux_h
    port map (
            O => \N__7734\,
            I => \N__7725\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7722\
        );

    \I__1667\ : InMux
    port map (
            O => \N__7732\,
            I => \N__7719\
        );

    \I__1666\ : InMux
    port map (
            O => \N__7729\,
            I => \N__7716\
        );

    \I__1665\ : InMux
    port map (
            O => \N__7728\,
            I => \N__7713\
        );

    \I__1664\ : Span4Mux_v
    port map (
            O => \N__7725\,
            I => \N__7710\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__7722\,
            I => \N__7705\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7719\,
            I => \N__7705\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__7716\,
            I => \N__7702\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7713\,
            I => \N__7699\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__7710\,
            I => \N__7692\
        );

    \I__1658\ : Span4Mux_h
    port map (
            O => \N__7705\,
            I => \N__7692\
        );

    \I__1657\ : Span4Mux_h
    port map (
            O => \N__7702\,
            I => \N__7692\
        );

    \I__1656\ : Odrv12
    port map (
            O => \N__7699\,
            I => \RAMENn_c\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__7692\,
            I => \RAMENn_c\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7687\,
            I => \N__7684\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__7684\,
            I => \N__7680\
        );

    \I__1652\ : InMux
    port map (
            O => \N__7683\,
            I => \N__7677\
        );

    \I__1651\ : Span4Mux_v
    port map (
            O => \N__7680\,
            I => \N__7674\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__7677\,
            I => \N__7671\
        );

    \I__1649\ : Span4Mux_v
    port map (
            O => \N__7674\,
            I => \N__7667\
        );

    \I__1648\ : Span4Mux_h
    port map (
            O => \N__7671\,
            I => \N__7664\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7670\,
            I => \N__7661\
        );

    \I__1646\ : Odrv4
    port map (
            O => \N__7667\,
            I => \REG_CYCLEm\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__7664\,
            I => \REG_CYCLEm\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7661\,
            I => \REG_CYCLEm\
        );

    \I__1643\ : IoInMux
    port map (
            O => \N__7654\,
            I => \N__7651\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__7651\,
            I => \N__7648\
        );

    \I__1641\ : IoSpan4Mux
    port map (
            O => \N__7648\,
            I => \N__7645\
        );

    \I__1640\ : Sp12to4
    port map (
            O => \N__7645\,
            I => \N__7642\
        );

    \I__1639\ : Span12Mux_s6_v
    port map (
            O => \N__7642\,
            I => \N__7639\
        );

    \I__1638\ : Span12Mux_h
    port map (
            O => \N__7639\,
            I => \N__7636\
        );

    \I__1637\ : Odrv12
    port map (
            O => \N__7636\,
            I => \DRDENn_c\
        );

    \I__1636\ : InMux
    port map (
            O => \N__7633\,
            I => \N__7630\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__7630\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1634\ : IoInMux
    port map (
            O => \N__7627\,
            I => \N__7624\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7624\,
            I => \N__7621\
        );

    \I__1632\ : Span12Mux_s0_v
    port map (
            O => \N__7621\,
            I => \N__7618\
        );

    \I__1631\ : Span12Mux_v
    port map (
            O => \N__7618\,
            I => \N__7615\
        );

    \I__1630\ : Odrv12
    port map (
            O => \N__7615\,
            I => \CMA_c_0\
        );

    \I__1629\ : CascadeMux
    port map (
            O => \N__7612\,
            I => \N__7609\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7609\,
            I => \N__7606\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__7606\,
            I => \N__7603\
        );

    \I__1626\ : Odrv12
    port map (
            O => \N__7603\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1625\ : InMux
    port map (
            O => \N__7600\,
            I => \N__7597\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7597\,
            I => \N__7594\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__7594\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1622\ : InMux
    port map (
            O => \N__7591\,
            I => \N__7587\
        );

    \I__1621\ : InMux
    port map (
            O => \N__7590\,
            I => \N__7584\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__7587\,
            I => \N__7579\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7584\,
            I => \N__7579\
        );

    \I__1618\ : Sp12to4
    port map (
            O => \N__7579\,
            I => \N__7576\
        );

    \I__1617\ : Span12Mux_v
    port map (
            O => \N__7576\,
            I => \N__7573\
        );

    \I__1616\ : Span12Mux_h
    port map (
            O => \N__7573\,
            I => \N__7570\
        );

    \I__1615\ : Odrv12
    port map (
            O => \N__7570\,
            I => \DRA_c_2\
        );

    \I__1614\ : InMux
    port map (
            O => \N__7567\,
            I => \N__7564\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__7564\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__7561\,
            I => \N__7558\
        );

    \I__1611\ : InMux
    port map (
            O => \N__7558\,
            I => \N__7555\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__7555\,
            I => \N__7552\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__7552\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1608\ : InMux
    port map (
            O => \N__7549\,
            I => \N__7546\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__7546\,
            I => \N__7543\
        );

    \I__1606\ : Span4Mux_h
    port map (
            O => \N__7543\,
            I => \N__7540\
        );

    \I__1605\ : Odrv4
    port map (
            O => \N__7540\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1604\ : InMux
    port map (
            O => \N__7537\,
            I => \N__7531\
        );

    \I__1603\ : InMux
    port map (
            O => \N__7536\,
            I => \N__7528\
        );

    \I__1602\ : InMux
    port map (
            O => \N__7535\,
            I => \N__7517\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7534\,
            I => \N__7517\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7531\,
            I => \N__7513\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__7528\,
            I => \N__7510\
        );

    \I__1598\ : InMux
    port map (
            O => \N__7527\,
            I => \N__7506\
        );

    \I__1597\ : InMux
    port map (
            O => \N__7526\,
            I => \N__7500\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7525\,
            I => \N__7493\
        );

    \I__1595\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7493\
        );

    \I__1594\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7493\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7522\,
            I => \N__7490\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__7517\,
            I => \N__7487\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7484\
        );

    \I__1590\ : Span4Mux_v
    port map (
            O => \N__7513\,
            I => \N__7479\
        );

    \I__1589\ : Span4Mux_h
    port map (
            O => \N__7510\,
            I => \N__7479\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7509\,
            I => \N__7476\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__7506\,
            I => \N__7473\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7505\,
            I => \N__7468\
        );

    \I__1585\ : InMux
    port map (
            O => \N__7504\,
            I => \N__7468\
        );

    \I__1584\ : InMux
    port map (
            O => \N__7503\,
            I => \N__7465\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__7500\,
            I => \N__7460\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7493\,
            I => \N__7460\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__7490\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__7487\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__7484\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1578\ : Odrv4
    port map (
            O => \N__7479\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7476\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__7473\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7468\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__7465\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1573\ : Odrv4
    port map (
            O => \N__7460\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7437\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7440\,
            I => \N__7434\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__7437\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1Z0Z_1\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7434\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1Z0Z_1\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7429\,
            I => \N__7426\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__7426\,
            I => \N__7423\
        );

    \I__1566\ : Odrv12
    port map (
            O => \N__7423\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_0\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7420\,
            I => \N__7416\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7413\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__7416\,
            I => \CPU_TACKm\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__7413\,
            I => \CPU_TACKm\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7408\,
            I => \N__7404\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__7407\,
            I => \N__7400\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7404\,
            I => \N__7397\
        );

    \I__1558\ : InMux
    port map (
            O => \N__7403\,
            I => \N__7394\
        );

    \I__1557\ : InMux
    port map (
            O => \N__7400\,
            I => \N__7391\
        );

    \I__1556\ : Span4Mux_v
    port map (
            O => \N__7397\,
            I => \N__7388\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7394\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__7391\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__7388\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1552\ : CascadeMux
    port map (
            O => \N__7381\,
            I => \N__7378\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7378\,
            I => \N__7375\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7375\,
            I => \N__7370\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7366\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7373\,
            I => \N__7363\
        );

    \I__1547\ : Span4Mux_h
    port map (
            O => \N__7370\,
            I => \N__7360\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7369\,
            I => \N__7357\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7366\,
            I => \U712_REG_SM.N_187\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7363\,
            I => \U712_REG_SM.N_187\
        );

    \I__1543\ : Odrv4
    port map (
            O => \N__7360\,
            I => \U712_REG_SM.N_187\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__7357\,
            I => \U712_REG_SM.N_187\
        );

    \I__1541\ : CascadeMux
    port map (
            O => \N__7348\,
            I => \N__7345\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7345\,
            I => \N__7341\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7344\,
            I => \N__7338\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7341\,
            I => \N__7333\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__7338\,
            I => \N__7330\
        );

    \I__1536\ : InMux
    port map (
            O => \N__7337\,
            I => \N__7325\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7336\,
            I => \N__7325\
        );

    \I__1534\ : Span4Mux_h
    port map (
            O => \N__7333\,
            I => \N__7322\
        );

    \I__1533\ : Span4Mux_v
    port map (
            O => \N__7330\,
            I => \N__7319\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__7325\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1531\ : Odrv4
    port map (
            O => \N__7322\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1530\ : Odrv4
    port map (
            O => \N__7319\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7312\,
            I => \N__7306\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7311\,
            I => \N__7306\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7306\,
            I => \REG_TACK\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7303\,
            I => \N__7300\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7300\,
            I => \N__7297\
        );

    \I__1524\ : Odrv4
    port map (
            O => \N__7297\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_0_a3_0\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7291\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7291\,
            I => \N__7288\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__7288\,
            I => \N__7285\
        );

    \I__1520\ : Odrv4
    port map (
            O => \N__7285\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__1519\ : InMux
    port map (
            O => \N__7282\,
            I => \N__7279\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7279\,
            I => \N__7276\
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__7276\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a3_0_a3_0\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7273\,
            I => \N__7259\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7272\,
            I => \N__7259\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7259\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7270\,
            I => \N__7254\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7269\,
            I => \N__7254\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7268\,
            I => \N__7247\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7267\,
            I => \N__7247\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7266\,
            I => \N__7247\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7259\,
            I => \U712_CHIP_RAM.N_96\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7254\,
            I => \U712_CHIP_RAM.N_96\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7247\,
            I => \U712_CHIP_RAM.N_96\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__7240\,
            I => \N__7235\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__7239\,
            I => \N__7232\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7229\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7235\,
            I => \N__7224\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7232\,
            I => \N__7224\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7229\,
            I => \N__7221\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__7224\,
            I => \N__7213\
        );

    \I__1498\ : Span4Mux_v
    port map (
            O => \N__7221\,
            I => \N__7213\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7220\,
            I => \N__7210\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7219\,
            I => \N__7207\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7218\,
            I => \N__7204\
        );

    \I__1494\ : Odrv4
    port map (
            O => \N__7213\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER16\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__7210\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER16\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7207\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER16\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7204\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER16\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7195\,
            I => \N__7192\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7192\,
            I => \N__7189\
        );

    \I__1488\ : Span4Mux_h
    port map (
            O => \N__7189\,
            I => \N__7186\
        );

    \I__1487\ : Odrv4
    port map (
            O => \N__7186\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__1486\ : CEMux
    port map (
            O => \N__7183\,
            I => \N__7179\
        );

    \I__1485\ : CEMux
    port map (
            O => \N__7182\,
            I => \N__7176\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7179\,
            I => \N__7173\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7176\,
            I => \N__7170\
        );

    \I__1482\ : Span4Mux_h
    port map (
            O => \N__7173\,
            I => \N__7167\
        );

    \I__1481\ : Odrv12
    port map (
            O => \N__7170\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__1480\ : Odrv4
    port map (
            O => \N__7167\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__1479\ : CascadeMux
    port map (
            O => \N__7162\,
            I => \N__7158\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__7161\,
            I => \N__7152\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7158\,
            I => \N__7146\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7157\,
            I => \N__7146\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7141\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7155\,
            I => \N__7141\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7152\,
            I => \N__7125\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7151\,
            I => \N__7125\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7146\,
            I => \N__7122\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7141\,
            I => \N__7119\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7110\
        );

    \I__1468\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7110\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7138\,
            I => \N__7110\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7137\,
            I => \N__7110\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7107\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7104\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7134\,
            I => \N__7099\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7133\,
            I => \N__7099\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7132\,
            I => \N__7096\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7131\,
            I => \N__7091\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7091\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7125\,
            I => \N__7086\
        );

    \I__1457\ : Span4Mux_h
    port map (
            O => \N__7122\,
            I => \N__7086\
        );

    \I__1456\ : Span4Mux_h
    port map (
            O => \N__7119\,
            I => \N__7083\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7110\,
            I => \N__7080\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7107\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7104\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__7099\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7096\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7091\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__7086\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__7083\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1447\ : Odrv12
    port map (
            O => \N__7080\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1446\ : InMux
    port map (
            O => \N__7063\,
            I => \N__7060\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7060\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_0_a3_0\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7057\,
            I => \N__7054\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7054\,
            I => \U712_CYCLE_TERM.N_214_i_0_en\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7051\,
            I => \N__7034\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7050\,
            I => \N__7034\
        );

    \I__1440\ : InMux
    port map (
            O => \N__7049\,
            I => \N__7031\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7048\,
            I => \N__7025\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7047\,
            I => \N__7022\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7046\,
            I => \N__7013\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7045\,
            I => \N__7013\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7044\,
            I => \N__7013\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7043\,
            I => \N__7013\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7042\,
            I => \N__7008\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7008\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__7040\,
            I => \N__7004\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__7039\,
            I => \N__6995\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7034\,
            I => \N__6988\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__7031\,
            I => \N__6985\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7030\,
            I => \N__6978\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7029\,
            I => \N__6978\
        );

    \I__1425\ : InMux
    port map (
            O => \N__7028\,
            I => \N__6978\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__7025\,
            I => \N__6975\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__7022\,
            I => \N__6968\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7013\,
            I => \N__6968\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7008\,
            I => \N__6968\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7007\,
            I => \N__6965\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7004\,
            I => \N__6962\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7003\,
            I => \N__6959\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7002\,
            I => \N__6954\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7001\,
            I => \N__6954\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6949\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6999\,
            I => \N__6949\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6998\,
            I => \N__6944\
        );

    \I__1412\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6944\
        );

    \I__1411\ : InMux
    port map (
            O => \N__6994\,
            I => \N__6941\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6993\,
            I => \N__6934\
        );

    \I__1409\ : InMux
    port map (
            O => \N__6992\,
            I => \N__6934\
        );

    \I__1408\ : InMux
    port map (
            O => \N__6991\,
            I => \N__6934\
        );

    \I__1407\ : Span4Mux_v
    port map (
            O => \N__6988\,
            I => \N__6927\
        );

    \I__1406\ : Span4Mux_v
    port map (
            O => \N__6985\,
            I => \N__6927\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__6978\,
            I => \N__6927\
        );

    \I__1404\ : Span4Mux_h
    port map (
            O => \N__6975\,
            I => \N__6922\
        );

    \I__1403\ : Span4Mux_h
    port map (
            O => \N__6968\,
            I => \N__6922\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__6965\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__6962\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__6959\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__6954\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6949\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__6944\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__6941\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__6934\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__6927\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__6922\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1392\ : CascadeMux
    port map (
            O => \N__6901\,
            I => \N__6894\
        );

    \I__1391\ : CascadeMux
    port map (
            O => \N__6900\,
            I => \N__6890\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__6899\,
            I => \N__6886\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__6898\,
            I => \N__6882\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__6897\,
            I => \N__6876\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6894\,
            I => \N__6873\
        );

    \I__1386\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6870\
        );

    \I__1385\ : InMux
    port map (
            O => \N__6890\,
            I => \N__6866\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6889\,
            I => \N__6861\
        );

    \I__1383\ : InMux
    port map (
            O => \N__6886\,
            I => \N__6861\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6885\,
            I => \N__6856\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6882\,
            I => \N__6856\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6849\
        );

    \I__1379\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6849\
        );

    \I__1378\ : InMux
    port map (
            O => \N__6879\,
            I => \N__6849\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6876\,
            I => \N__6846\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__6873\,
            I => \N__6839\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__6870\,
            I => \N__6839\
        );

    \I__1374\ : InMux
    port map (
            O => \N__6869\,
            I => \N__6836\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__6866\,
            I => \N__6829\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__6861\,
            I => \N__6829\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__6856\,
            I => \N__6829\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__6849\,
            I => \N__6823\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__6846\,
            I => \N__6823\
        );

    \I__1368\ : InMux
    port map (
            O => \N__6845\,
            I => \N__6820\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6844\,
            I => \N__6817\
        );

    \I__1366\ : Span4Mux_v
    port map (
            O => \N__6839\,
            I => \N__6810\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__6836\,
            I => \N__6810\
        );

    \I__1364\ : Span4Mux_v
    port map (
            O => \N__6829\,
            I => \N__6810\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6828\,
            I => \N__6807\
        );

    \I__1362\ : Odrv4
    port map (
            O => \N__6823\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6820\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__6817\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1359\ : Odrv4
    port map (
            O => \N__6810\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__6807\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1357\ : IoInMux
    port map (
            O => \N__6796\,
            I => \N__6793\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__6793\,
            I => \N__6790\
        );

    \I__1355\ : Span4Mux_s3_h
    port map (
            O => \N__6790\,
            I => \N__6787\
        );

    \I__1354\ : Sp12to4
    port map (
            O => \N__6787\,
            I => \N__6784\
        );

    \I__1353\ : Span12Mux_v
    port map (
            O => \N__6784\,
            I => \N__6781\
        );

    \I__1352\ : Span12Mux_h
    port map (
            O => \N__6781\,
            I => \N__6778\
        );

    \I__1351\ : Odrv12
    port map (
            O => \N__6778\,
            I => \CMA_c_5\
        );

    \I__1350\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6772\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6772\,
            I => \N__6769\
        );

    \I__1348\ : Span4Mux_v
    port map (
            O => \N__6769\,
            I => \N__6766\
        );

    \I__1347\ : Sp12to4
    port map (
            O => \N__6766\,
            I => \N__6763\
        );

    \I__1346\ : Span12Mux_h
    port map (
            O => \N__6763\,
            I => \N__6760\
        );

    \I__1345\ : Odrv12
    port map (
            O => \N__6760\,
            I => \A_c_7\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__6757\,
            I => \U712_CHIP_RAM.N_316_cascade_\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6754\,
            I => \N__6751\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6751\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6748\,
            I => \N__6745\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__6745\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6742\,
            I => \N__6736\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6741\,
            I => \N__6736\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6736\,
            I => \N__6733\
        );

    \I__1336\ : Span4Mux_h
    port map (
            O => \N__6733\,
            I => \N__6728\
        );

    \I__1335\ : InMux
    port map (
            O => \N__6732\,
            I => \N__6723\
        );

    \I__1334\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6723\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__6728\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6723\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__6718\,
            I => \N__6715\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6715\,
            I => \N__6709\
        );

    \I__1329\ : InMux
    port map (
            O => \N__6714\,
            I => \N__6709\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__6709\,
            I => \N__6706\
        );

    \I__1327\ : Span4Mux_h
    port map (
            O => \N__6706\,
            I => \N__6703\
        );

    \I__1326\ : Sp12to4
    port map (
            O => \N__6703\,
            I => \N__6700\
        );

    \I__1325\ : Span12Mux_v
    port map (
            O => \N__6700\,
            I => \N__6697\
        );

    \I__1324\ : Span12Mux_h
    port map (
            O => \N__6697\,
            I => \N__6694\
        );

    \I__1323\ : Odrv12
    port map (
            O => \N__6694\,
            I => \A_c_14\
        );

    \I__1322\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6688\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6688\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6685\,
            I => \N__6682\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6682\,
            I => \N__6679\
        );

    \I__1318\ : Span4Mux_h
    port map (
            O => \N__6679\,
            I => \N__6670\
        );

    \I__1317\ : InMux
    port map (
            O => \N__6678\,
            I => \N__6667\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6677\,
            I => \N__6662\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6676\,
            I => \N__6662\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6659\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6656\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6673\,
            I => \N__6653\
        );

    \I__1311\ : Odrv4
    port map (
            O => \N__6670\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__6667\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6662\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__6659\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__6656\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__6653\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1305\ : CEMux
    port map (
            O => \N__6640\,
            I => \N__6637\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__6637\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_3_0_0\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6634\,
            I => \N__6631\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__6631\,
            I => \N__6627\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6630\,
            I => \N__6623\
        );

    \I__1300\ : Span4Mux_v
    port map (
            O => \N__6627\,
            I => \N__6618\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6626\,
            I => \N__6615\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6623\,
            I => \N__6612\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6622\,
            I => \N__6609\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6621\,
            I => \N__6606\
        );

    \I__1295\ : Odrv4
    port map (
            O => \N__6618\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6615\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1293\ : Odrv4
    port map (
            O => \N__6612\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__6609\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__6606\,
            I => \U712_CHIP_RAM.N_180\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6592\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6592\,
            I => \N__6589\
        );

    \I__1288\ : Span4Mux_v
    port map (
            O => \N__6589\,
            I => \N__6586\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__6586\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a3_2_1_0\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6578\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__6582\,
            I => \N__6575\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6581\,
            I => \N__6572\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6578\,
            I => \N__6569\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6575\,
            I => \N__6566\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6572\,
            I => \U712_CHIP_RAM.N_254_2\
        );

    \I__1280\ : Odrv4
    port map (
            O => \N__6569\,
            I => \U712_CHIP_RAM.N_254_2\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6566\,
            I => \U712_CHIP_RAM.N_254_2\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6559\,
            I => \N__6556\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6556\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1276\ : IoInMux
    port map (
            O => \N__6553\,
            I => \N__6550\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6550\,
            I => \N__6547\
        );

    \I__1274\ : IoSpan4Mux
    port map (
            O => \N__6547\,
            I => \N__6544\
        );

    \I__1273\ : Span4Mux_s2_h
    port map (
            O => \N__6544\,
            I => \N__6541\
        );

    \I__1272\ : Sp12to4
    port map (
            O => \N__6541\,
            I => \N__6538\
        );

    \I__1271\ : Span12Mux_h
    port map (
            O => \N__6538\,
            I => \N__6535\
        );

    \I__1270\ : Odrv12
    port map (
            O => \N__6535\,
            I => \CMA_c_7\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6532\,
            I => \N__6529\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6529\,
            I => \N__6526\
        );

    \I__1267\ : Span12Mux_v
    port map (
            O => \N__6526\,
            I => \N__6523\
        );

    \I__1266\ : Span12Mux_h
    port map (
            O => \N__6523\,
            I => \N__6520\
        );

    \I__1265\ : Odrv12
    port map (
            O => \N__6520\,
            I => \A_c_15\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6517\,
            I => \N__6514\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__6514\,
            I => \N__6511\
        );

    \I__1262\ : Span4Mux_v
    port map (
            O => \N__6511\,
            I => \N__6508\
        );

    \I__1261\ : Sp12to4
    port map (
            O => \N__6508\,
            I => \N__6505\
        );

    \I__1260\ : Span12Mux_h
    port map (
            O => \N__6505\,
            I => \N__6502\
        );

    \I__1259\ : Odrv12
    port map (
            O => \N__6502\,
            I => \A_c_8\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__6499\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6493\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__6493\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6490\,
            I => \N__6487\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6487\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6481\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__6481\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6475\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6475\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__6472\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6469\,
            I => \N__6466\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6466\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1246\ : IoInMux
    port map (
            O => \N__6463\,
            I => \N__6460\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6460\,
            I => \N__6457\
        );

    \I__1244\ : Span12Mux_s7_v
    port map (
            O => \N__6457\,
            I => \N__6454\
        );

    \I__1243\ : Odrv12
    port map (
            O => \N__6454\,
            I => \CMA_c_1\
        );

    \I__1242\ : CEMux
    port map (
            O => \N__6451\,
            I => \N__6448\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6448\,
            I => \N__6445\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__6445\,
            I => \U712_CYCLE_TERM.N_214_i_0_en_0\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6442\,
            I => \N__6439\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6439\,
            I => \N__6436\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__6436\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_1\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6433\,
            I => \N__6430\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6430\,
            I => \N__6427\
        );

    \I__1234\ : Odrv4
    port map (
            O => \N__6427\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_3\
        );

    \I__1233\ : IoInMux
    port map (
            O => \N__6424\,
            I => \N__6421\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6421\,
            I => \N__6418\
        );

    \I__1231\ : Span4Mux_s2_v
    port map (
            O => \N__6418\,
            I => \N__6415\
        );

    \I__1230\ : Span4Mux_v
    port map (
            O => \N__6415\,
            I => \N__6412\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__6412\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1228\ : IoInMux
    port map (
            O => \N__6409\,
            I => \N__6406\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6406\,
            I => \N__6403\
        );

    \I__1226\ : Span4Mux_s2_v
    port map (
            O => \N__6403\,
            I => \N__6400\
        );

    \I__1225\ : Span4Mux_v
    port map (
            O => \N__6400\,
            I => \N__6397\
        );

    \I__1224\ : Span4Mux_v
    port map (
            O => \N__6397\,
            I => \N__6394\
        );

    \I__1223\ : Span4Mux_h
    port map (
            O => \N__6394\,
            I => \N__6391\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__6391\,
            I => \CRCSn_c\
        );

    \I__1221\ : IoInMux
    port map (
            O => \N__6388\,
            I => \N__6385\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6385\,
            I => \N__6382\
        );

    \I__1219\ : Span4Mux_s0_h
    port map (
            O => \N__6382\,
            I => \N__6379\
        );

    \I__1218\ : Span4Mux_h
    port map (
            O => \N__6379\,
            I => \N__6376\
        );

    \I__1217\ : Sp12to4
    port map (
            O => \N__6376\,
            I => \N__6373\
        );

    \I__1216\ : Span12Mux_s9_v
    port map (
            O => \N__6373\,
            I => \N__6370\
        );

    \I__1215\ : Span12Mux_h
    port map (
            O => \N__6370\,
            I => \N__6367\
        );

    \I__1214\ : Odrv12
    port map (
            O => \N__6367\,
            I => \WEn_c\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6364\,
            I => \N__6361\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6361\,
            I => \N__6358\
        );

    \I__1211\ : Span12Mux_v
    port map (
            O => \N__6358\,
            I => \N__6355\
        );

    \I__1210\ : Span12Mux_h
    port map (
            O => \N__6355\,
            I => \N__6352\
        );

    \I__1209\ : Odrv12
    port map (
            O => \N__6352\,
            I => \A_c_19\
        );

    \I__1208\ : CascadeMux
    port map (
            O => \N__6349\,
            I => \N__6346\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6346\,
            I => \N__6343\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__6343\,
            I => \N__6340\
        );

    \I__1205\ : Span12Mux_v
    port map (
            O => \N__6340\,
            I => \N__6337\
        );

    \I__1204\ : Span12Mux_h
    port map (
            O => \N__6337\,
            I => \N__6334\
        );

    \I__1203\ : Odrv12
    port map (
            O => \N__6334\,
            I => \RAS0n_c\
        );

    \I__1202\ : IoInMux
    port map (
            O => \N__6331\,
            I => \N__6328\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6328\,
            I => \N__6325\
        );

    \I__1200\ : IoSpan4Mux
    port map (
            O => \N__6325\,
            I => \N__6322\
        );

    \I__1199\ : Span4Mux_s2_h
    port map (
            O => \N__6322\,
            I => \N__6319\
        );

    \I__1198\ : Sp12to4
    port map (
            O => \N__6319\,
            I => \N__6316\
        );

    \I__1197\ : Span12Mux_h
    port map (
            O => \N__6316\,
            I => \N__6313\
        );

    \I__1196\ : Odrv12
    port map (
            O => \N__6313\,
            I => \CMA_c_9\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6307\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__6307\,
            I => \N__6304\
        );

    \I__1193\ : Span12Mux_v
    port map (
            O => \N__6304\,
            I => \N__6301\
        );

    \I__1192\ : Span12Mux_h
    port map (
            O => \N__6301\,
            I => \N__6298\
        );

    \I__1191\ : Odrv12
    port map (
            O => \N__6298\,
            I => \A_c_17\
        );

    \I__1190\ : IoInMux
    port map (
            O => \N__6295\,
            I => \N__6292\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__6292\,
            I => \N__6289\
        );

    \I__1188\ : IoSpan4Mux
    port map (
            O => \N__6289\,
            I => \N__6286\
        );

    \I__1187\ : Span4Mux_s3_h
    port map (
            O => \N__6286\,
            I => \N__6283\
        );

    \I__1186\ : Span4Mux_v
    port map (
            O => \N__6283\,
            I => \N__6280\
        );

    \I__1185\ : Span4Mux_h
    port map (
            O => \N__6280\,
            I => \N__6277\
        );

    \I__1184\ : Sp12to4
    port map (
            O => \N__6277\,
            I => \N__6274\
        );

    \I__1183\ : Odrv12
    port map (
            O => \N__6274\,
            I => \CMA_c_8\
        );

    \I__1182\ : IoInMux
    port map (
            O => \N__6271\,
            I => \N__6268\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6268\,
            I => \N__6265\
        );

    \I__1180\ : IoSpan4Mux
    port map (
            O => \N__6265\,
            I => \N__6262\
        );

    \I__1179\ : Span4Mux_s3_h
    port map (
            O => \N__6262\,
            I => \N__6259\
        );

    \I__1178\ : Sp12to4
    port map (
            O => \N__6259\,
            I => \N__6256\
        );

    \I__1177\ : Span12Mux_s8_h
    port map (
            O => \N__6256\,
            I => \N__6253\
        );

    \I__1176\ : Span12Mux_v
    port map (
            O => \N__6253\,
            I => \N__6250\
        );

    \I__1175\ : Odrv12
    port map (
            O => \N__6250\,
            I => \CMA_c_6\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6242\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6239\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__6245\,
            I => \N__6236\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6242\,
            I => \N__6230\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6239\,
            I => \N__6230\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6236\,
            I => \N__6227\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6235\,
            I => \N__6224\
        );

    \I__1167\ : Span4Mux_v
    port map (
            O => \N__6230\,
            I => \N__6221\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6227\,
            I => \N__6216\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6224\,
            I => \N__6216\
        );

    \I__1164\ : Odrv4
    port map (
            O => \N__6221\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__6216\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6211\,
            I => \N__6207\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6210\,
            I => \N__6204\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__6207\,
            I => \N__6200\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6204\,
            I => \N__6197\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__6203\,
            I => \N__6193\
        );

    \I__1157\ : Span4Mux_v
    port map (
            O => \N__6200\,
            I => \N__6187\
        );

    \I__1156\ : Span4Mux_h
    port map (
            O => \N__6197\,
            I => \N__6187\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6196\,
            I => \N__6182\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6193\,
            I => \N__6179\
        );

    \I__1153\ : InMux
    port map (
            O => \N__6192\,
            I => \N__6176\
        );

    \I__1152\ : Span4Mux_v
    port map (
            O => \N__6187\,
            I => \N__6173\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6186\,
            I => \N__6168\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6168\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6182\,
            I => \N__6165\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6179\,
            I => \N__6162\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6176\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1146\ : Odrv4
    port map (
            O => \N__6173\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6168\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1144\ : Odrv4
    port map (
            O => \N__6165\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1143\ : Odrv4
    port map (
            O => \N__6162\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1142\ : IoInMux
    port map (
            O => \N__6151\,
            I => \N__6148\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__6148\,
            I => \N__6145\
        );

    \I__1140\ : Span4Mux_s1_v
    port map (
            O => \N__6145\,
            I => \N__6142\
        );

    \I__1139\ : Sp12to4
    port map (
            O => \N__6142\,
            I => \N__6139\
        );

    \I__1138\ : Span12Mux_h
    port map (
            O => \N__6139\,
            I => \N__6136\
        );

    \I__1137\ : Odrv12
    port map (
            O => \N__6136\,
            I => \CMA_c_10\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__6133\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_2_cascade_\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6130\,
            I => \N__6126\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6129\,
            I => \N__6123\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6126\,
            I => \U712_CHIP_RAM.N_221\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6123\,
            I => \U712_CHIP_RAM.N_221\
        );

    \I__1131\ : CEMux
    port map (
            O => \N__6118\,
            I => \N__6114\
        );

    \I__1130\ : CEMux
    port map (
            O => \N__6117\,
            I => \N__6111\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6114\,
            I => \N__6106\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6111\,
            I => \N__6106\
        );

    \I__1127\ : Span4Mux_v
    port map (
            O => \N__6106\,
            I => \N__6103\
        );

    \I__1126\ : Span4Mux_h
    port map (
            O => \N__6103\,
            I => \N__6100\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__6100\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6094\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6094\,
            I => \N__6088\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6085\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6080\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6091\,
            I => \N__6080\
        );

    \I__1119\ : Odrv12
    port map (
            O => \N__6088\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6085\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__6080\,
            I => \U712_CHIP_RAM.N_305\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__6073\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_cascade_\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6070\,
            I => \N__6067\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6067\,
            I => \N__6063\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6066\,
            I => \N__6059\
        );

    \I__1112\ : Span4Mux_v
    port map (
            O => \N__6063\,
            I => \N__6056\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6062\,
            I => \N__6053\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6059\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__6056\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6053\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1107\ : IoInMux
    port map (
            O => \N__6046\,
            I => \N__6043\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6043\,
            I => \N__6040\
        );

    \I__1105\ : IoSpan4Mux
    port map (
            O => \N__6040\,
            I => \N__6037\
        );

    \I__1104\ : Span4Mux_s3_h
    port map (
            O => \N__6037\,
            I => \N__6034\
        );

    \I__1103\ : Sp12to4
    port map (
            O => \N__6034\,
            I => \N__6031\
        );

    \I__1102\ : Span12Mux_h
    port map (
            O => \N__6031\,
            I => \N__6027\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6030\,
            I => \N__6024\
        );

    \I__1100\ : Odrv12
    port map (
            O => \N__6027\,
            I => \CLK_EN_c\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6024\,
            I => \CLK_EN_c\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__6019\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__6016\,
            I => \N__6013\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6013\,
            I => \N__6009\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__6012\,
            I => \N__6006\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6009\,
            I => \N__5998\
        );

    \I__1093\ : InMux
    port map (
            O => \N__6006\,
            I => \N__5995\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__6005\,
            I => \N__5992\
        );

    \I__1091\ : InMux
    port map (
            O => \N__6004\,
            I => \N__5980\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6003\,
            I => \N__5980\
        );

    \I__1089\ : InMux
    port map (
            O => \N__6002\,
            I => \N__5980\
        );

    \I__1088\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5980\
        );

    \I__1087\ : Span4Mux_h
    port map (
            O => \N__5998\,
            I => \N__5976\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5995\,
            I => \N__5973\
        );

    \I__1085\ : InMux
    port map (
            O => \N__5992\,
            I => \N__5970\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5991\,
            I => \N__5967\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5990\,
            I => \N__5964\
        );

    \I__1082\ : InMux
    port map (
            O => \N__5989\,
            I => \N__5961\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__5980\,
            I => \N__5958\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5979\,
            I => \N__5955\
        );

    \I__1079\ : Odrv4
    port map (
            O => \N__5976\,
            I => \U712_CHIP_RAM.N_10\
        );

    \I__1078\ : Odrv4
    port map (
            O => \N__5973\,
            I => \U712_CHIP_RAM.N_10\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5970\,
            I => \U712_CHIP_RAM.N_10\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5967\,
            I => \U712_CHIP_RAM.N_10\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__5964\,
            I => \U712_CHIP_RAM.N_10\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__5961\,
            I => \U712_CHIP_RAM.N_10\
        );

    \I__1073\ : Odrv4
    port map (
            O => \N__5958\,
            I => \U712_CHIP_RAM.N_10\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5955\,
            I => \U712_CHIP_RAM.N_10\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__5938\,
            I => \N__5935\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5935\,
            I => \N__5932\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5932\,
            I => \U712_CHIP_RAM.N_260\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__5929\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_66_0_i_1_cascade_\
        );

    \I__1067\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5920\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5920\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5920\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9MVM2Z0Z_1\
        );

    \I__1064\ : InMux
    port map (
            O => \N__5917\,
            I => \N__5914\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__5914\,
            I => \U712_CHIP_RAM.N_222\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__5911\,
            I => \N__5907\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5910\,
            I => \N__5904\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5907\,
            I => \N__5901\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5904\,
            I => \N__5898\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__5901\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa\
        );

    \I__1057\ : Odrv12
    port map (
            O => \N__5898\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__5893\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_9_0_cascade_\
        );

    \I__1055\ : IoInMux
    port map (
            O => \N__5890\,
            I => \N__5887\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5887\,
            I => \N__5884\
        );

    \I__1053\ : Span4Mux_s1_v
    port map (
            O => \N__5884\,
            I => \N__5881\
        );

    \I__1052\ : Span4Mux_v
    port map (
            O => \N__5881\,
            I => \N__5878\
        );

    \I__1051\ : Span4Mux_v
    port map (
            O => \N__5878\,
            I => \N__5875\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__5875\,
            I => \N__5870\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5867\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5864\
        );

    \I__1047\ : Span4Mux_h
    port map (
            O => \N__5870\,
            I => \N__5857\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__5867\,
            I => \N__5857\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5864\,
            I => \N__5857\
        );

    \I__1044\ : Span4Mux_h
    port map (
            O => \N__5857\,
            I => \N__5853\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5856\,
            I => \N__5850\
        );

    \I__1042\ : Odrv4
    port map (
            O => \N__5853\,
            I => \DBENn_c\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5850\,
            I => \DBENn_c\
        );

    \I__1040\ : InMux
    port map (
            O => \N__5845\,
            I => \N__5842\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__5842\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_3_0\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__5839\,
            I => \U712_CHIP_RAM.N_305_cascade_\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__5836\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_0_cascade_\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__5833\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5830\,
            I => \N__5827\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5827\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5824\,
            I => \N__5821\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5821\,
            I => \N__5818\
        );

    \I__1031\ : Span4Mux_v
    port map (
            O => \N__5818\,
            I => \N__5815\
        );

    \I__1030\ : Sp12to4
    port map (
            O => \N__5815\,
            I => \N__5812\
        );

    \I__1029\ : Span12Mux_h
    port map (
            O => \N__5812\,
            I => \N__5809\
        );

    \I__1028\ : Span12Mux_v
    port map (
            O => \N__5809\,
            I => \N__5806\
        );

    \I__1027\ : Odrv12
    port map (
            O => \N__5806\,
            I => \A_c_3\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5803\,
            I => \N__5800\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5800\,
            I => \N__5797\
        );

    \I__1024\ : Span4Mux_v
    port map (
            O => \N__5797\,
            I => \N__5794\
        );

    \I__1023\ : Sp12to4
    port map (
            O => \N__5794\,
            I => \N__5791\
        );

    \I__1022\ : Span12Mux_h
    port map (
            O => \N__5791\,
            I => \N__5788\
        );

    \I__1021\ : Odrv12
    port map (
            O => \N__5788\,
            I => \A_c_10\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5785\,
            I => \N__5782\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5782\,
            I => \N__5779\
        );

    \I__1018\ : Span4Mux_v
    port map (
            O => \N__5779\,
            I => \N__5776\
        );

    \I__1017\ : Sp12to4
    port map (
            O => \N__5776\,
            I => \N__5773\
        );

    \I__1016\ : Span12Mux_h
    port map (
            O => \N__5773\,
            I => \N__5770\
        );

    \I__1015\ : Odrv12
    port map (
            O => \N__5770\,
            I => \A_c_9\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5767\,
            I => \N__5764\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__5764\,
            I => \N__5761\
        );

    \I__1012\ : Span12Mux_h
    port map (
            O => \N__5761\,
            I => \N__5758\
        );

    \I__1011\ : Span12Mux_v
    port map (
            O => \N__5758\,
            I => \N__5755\
        );

    \I__1010\ : Odrv12
    port map (
            O => \N__5755\,
            I => \A_c_2\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5752\,
            I => \N__5749\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5749\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_0\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__5746\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_1_cascade_\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__5743\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_2_cascade_\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5740\,
            I => \N__5736\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5739\,
            I => \N__5733\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5736\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__5733\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5725\,
            I => \N__5722\
        );

    \I__999\ : Span4Mux_v
    port map (
            O => \N__5722\,
            I => \N__5719\
        );

    \I__998\ : Odrv4
    port map (
            O => \N__5719\,
            I => \TACK_EN_i_ess\
        );

    \I__997\ : InMux
    port map (
            O => \N__5716\,
            I => \N__5713\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5713\,
            I => \N__5710\
        );

    \I__995\ : Span4Mux_v
    port map (
            O => \N__5710\,
            I => \N__5707\
        );

    \I__994\ : Span4Mux_v
    port map (
            O => \N__5707\,
            I => \N__5704\
        );

    \I__993\ : Sp12to4
    port map (
            O => \N__5704\,
            I => \N__5701\
        );

    \I__992\ : Span12Mux_h
    port map (
            O => \N__5701\,
            I => \N__5698\
        );

    \I__991\ : Odrv12
    port map (
            O => \N__5698\,
            I => \A_c_18\
        );

    \I__990\ : InMux
    port map (
            O => \N__5695\,
            I => \N__5692\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__5692\,
            I => \N__5689\
        );

    \I__988\ : Span4Mux_v
    port map (
            O => \N__5689\,
            I => \N__5686\
        );

    \I__987\ : Span4Mux_v
    port map (
            O => \N__5686\,
            I => \N__5683\
        );

    \I__986\ : Sp12to4
    port map (
            O => \N__5683\,
            I => \N__5680\
        );

    \I__985\ : Span12Mux_h
    port map (
            O => \N__5680\,
            I => \N__5677\
        );

    \I__984\ : Odrv12
    port map (
            O => \N__5677\,
            I => \A_c_16\
        );

    \I__983\ : CascadeMux
    port map (
            O => \N__5674\,
            I => \N__5671\
        );

    \I__982\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5668\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5668\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__980\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5662\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__5662\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__978\ : IoInMux
    port map (
            O => \N__5659\,
            I => \N__5656\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5656\,
            I => \N__5653\
        );

    \I__976\ : Span12Mux_s5_v
    port map (
            O => \N__5653\,
            I => \N__5650\
        );

    \I__975\ : Odrv12
    port map (
            O => \N__5650\,
            I => \CMA_c_2\
        );

    \I__974\ : IoInMux
    port map (
            O => \N__5647\,
            I => \N__5644\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__5644\,
            I => \N__5641\
        );

    \I__972\ : Span12Mux_s8_h
    port map (
            O => \N__5641\,
            I => \N__5638\
        );

    \I__971\ : Span12Mux_v
    port map (
            O => \N__5638\,
            I => \N__5635\
        );

    \I__970\ : Odrv12
    port map (
            O => \N__5635\,
            I => \CMA_c_3\
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__5632\,
            I => \U712_CHIP_RAM.un1_CMA30_0_i_cascade_\
        );

    \I__968\ : InMux
    port map (
            O => \N__5629\,
            I => \N__5626\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__5626\,
            I => \N__5623\
        );

    \I__966\ : Sp12to4
    port map (
            O => \N__5623\,
            I => \N__5620\
        );

    \I__965\ : Span12Mux_v
    port map (
            O => \N__5620\,
            I => \N__5617\
        );

    \I__964\ : Span12Mux_h
    port map (
            O => \N__5617\,
            I => \N__5614\
        );

    \I__963\ : Odrv12
    port map (
            O => \N__5614\,
            I => \A_c_5\
        );

    \I__962\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5608\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__5608\,
            I => \N__5605\
        );

    \I__960\ : Span4Mux_v
    port map (
            O => \N__5605\,
            I => \N__5602\
        );

    \I__959\ : Sp12to4
    port map (
            O => \N__5602\,
            I => \N__5599\
        );

    \I__958\ : Span12Mux_h
    port map (
            O => \N__5599\,
            I => \N__5596\
        );

    \I__957\ : Odrv12
    port map (
            O => \N__5596\,
            I => \A_c_12\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__5593\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_cascade_\
        );

    \I__955\ : InMux
    port map (
            O => \N__5590\,
            I => \bfn_10_14_0_\
        );

    \I__954\ : InMux
    port map (
            O => \N__5587\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__953\ : InMux
    port map (
            O => \N__5584\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__952\ : InMux
    port map (
            O => \N__5581\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__5578\,
            I => \N__5575\
        );

    \I__950\ : InMux
    port map (
            O => \N__5575\,
            I => \N__5571\
        );

    \I__949\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5568\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5571\,
            I => \N__5565\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__5568\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__946\ : Odrv4
    port map (
            O => \N__5565\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__945\ : InMux
    port map (
            O => \N__5560\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__944\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5553\
        );

    \I__943\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5550\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5553\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5550\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__940\ : InMux
    port map (
            O => \N__5545\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__939\ : InMux
    port map (
            O => \N__5542\,
            I => \N__5538\
        );

    \I__938\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5535\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__5538\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5535\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__935\ : InMux
    port map (
            O => \N__5530\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__934\ : InMux
    port map (
            O => \N__5527\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__933\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5521\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__5521\,
            I => \U712_CHIP_RAM.N_323\
        );

    \I__931\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5515\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__5515\,
            I => \U712_CHIP_RAM.N_240\
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__5512\,
            I => \U712_CHIP_RAM.N_10_cascade_\
        );

    \I__928\ : CascadeMux
    port map (
            O => \N__5509\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER16_cascade_\
        );

    \I__927\ : InMux
    port map (
            O => \N__5506\,
            I => \N__5503\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5503\,
            I => \N__5500\
        );

    \I__925\ : Odrv4
    port map (
            O => \N__5500\,
            I => \U712_CHIP_RAM.N_328\
        );

    \I__924\ : InMux
    port map (
            O => \N__5497\,
            I => \N__5494\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5494\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__5491\,
            I => \U712_CHIP_RAM.N_328_cascade_\
        );

    \I__921\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5484\
        );

    \I__920\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5481\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__5484\,
            I => \U712_CHIP_RAM.N_177\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5481\,
            I => \U712_CHIP_RAM.N_177\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__5476\,
            I => \U712_CHIP_RAM.N_251_cascade_\
        );

    \I__916\ : InMux
    port map (
            O => \N__5473\,
            I => \N__5470\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__5470\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__5467\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a3_3_2_0_cascade_\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__5464\,
            I => \U712_CHIP_RAM.N_242_cascade_\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__5461\,
            I => \U712_CHIP_RAM.N_188_cascade_\
        );

    \I__911\ : CEMux
    port map (
            O => \N__5458\,
            I => \N__5455\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__5455\,
            I => \N__5452\
        );

    \I__909\ : Sp12to4
    port map (
            O => \N__5452\,
            I => \N__5449\
        );

    \I__908\ : Odrv12
    port map (
            O => \N__5449\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0_0\
        );

    \I__907\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5438\
        );

    \I__906\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5438\
        );

    \I__905\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5433\
        );

    \I__904\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5433\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5438\,
            I => \U712_CHIP_RAM.N_306\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5433\,
            I => \U712_CHIP_RAM.N_306\
        );

    \I__901\ : InMux
    port map (
            O => \N__5428\,
            I => \N__5423\
        );

    \I__900\ : InMux
    port map (
            O => \N__5427\,
            I => \N__5420\
        );

    \I__899\ : InMux
    port map (
            O => \N__5426\,
            I => \N__5417\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__5423\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5420\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5417\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__895\ : InMux
    port map (
            O => \N__5410\,
            I => \N__5407\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__5407\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0\
        );

    \I__893\ : InMux
    port map (
            O => \N__5404\,
            I => \N__5401\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5401\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0\
        );

    \I__891\ : InMux
    port map (
            O => \N__5398\,
            I => \N__5394\
        );

    \I__890\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5391\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__5394\,
            I => \U712_CHIP_RAM.N_238\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5391\,
            I => \U712_CHIP_RAM.N_238\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__5386\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_\
        );

    \I__886\ : InMux
    port map (
            O => \N__5383\,
            I => \N__5379\
        );

    \I__885\ : InMux
    port map (
            O => \N__5382\,
            I => \N__5376\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5379\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__5376\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__882\ : InMux
    port map (
            O => \N__5371\,
            I => \N__5368\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5368\,
            I => \N__5365\
        );

    \I__880\ : Span4Mux_v
    port map (
            O => \N__5365\,
            I => \N__5362\
        );

    \I__879\ : Odrv4
    port map (
            O => \N__5362\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__878\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5356\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5356\,
            I => \N__5353\
        );

    \I__876\ : Span12Mux_v
    port map (
            O => \N__5353\,
            I => \N__5350\
        );

    \I__875\ : Span12Mux_h
    port map (
            O => \N__5350\,
            I => \N__5347\
        );

    \I__874\ : Odrv12
    port map (
            O => \N__5347\,
            I => \A_c_4\
        );

    \I__873\ : InMux
    port map (
            O => \N__5344\,
            I => \N__5341\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5341\,
            I => \N__5338\
        );

    \I__871\ : Span4Mux_v
    port map (
            O => \N__5338\,
            I => \N__5335\
        );

    \I__870\ : Sp12to4
    port map (
            O => \N__5335\,
            I => \N__5332\
        );

    \I__869\ : Span12Mux_h
    port map (
            O => \N__5332\,
            I => \N__5329\
        );

    \I__868\ : Odrv12
    port map (
            O => \N__5329\,
            I => \A_c_11\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__5326\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\
        );

    \I__866\ : SRMux
    port map (
            O => \N__5323\,
            I => \N__5320\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5320\,
            I => \N__5317\
        );

    \I__864\ : Odrv12
    port map (
            O => \N__5317\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__5314\,
            I => \N__5311\
        );

    \I__862\ : InMux
    port map (
            O => \N__5311\,
            I => \N__5304\
        );

    \I__861\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5304\
        );

    \I__860\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5301\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5304\,
            I => \N__5296\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5301\,
            I => \N__5296\
        );

    \I__857\ : Odrv4
    port map (
            O => \N__5296\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__856\ : InMux
    port map (
            O => \N__5293\,
            I => \N__5286\
        );

    \I__855\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5286\
        );

    \I__854\ : InMux
    port map (
            O => \N__5291\,
            I => \N__5283\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5286\,
            I => \U712_REG_SM.N_209\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5283\,
            I => \U712_REG_SM.N_209\
        );

    \I__851\ : InMux
    port map (
            O => \N__5278\,
            I => \N__5275\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5275\,
            I => \N__5272\
        );

    \I__849\ : Span4Mux_v
    port map (
            O => \N__5272\,
            I => \N__5269\
        );

    \I__848\ : Span4Mux_v
    port map (
            O => \N__5269\,
            I => \N__5264\
        );

    \I__847\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5261\
        );

    \I__846\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5258\
        );

    \I__845\ : Span4Mux_v
    port map (
            O => \N__5264\,
            I => \N__5253\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5261\,
            I => \N__5253\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__5258\,
            I => \N__5250\
        );

    \I__842\ : Span4Mux_v
    port map (
            O => \N__5253\,
            I => \N__5247\
        );

    \I__841\ : Span12Mux_h
    port map (
            O => \N__5250\,
            I => \N__5244\
        );

    \I__840\ : IoSpan4Mux
    port map (
            O => \N__5247\,
            I => \N__5241\
        );

    \I__839\ : Span12Mux_v
    port map (
            O => \N__5244\,
            I => \N__5238\
        );

    \I__838\ : IoSpan4Mux
    port map (
            O => \N__5241\,
            I => \N__5235\
        );

    \I__837\ : Odrv12
    port map (
            O => \N__5238\,
            I => \AWEn_c\
        );

    \I__836\ : Odrv4
    port map (
            O => \N__5235\,
            I => \AWEn_c\
        );

    \I__835\ : IoInMux
    port map (
            O => \N__5230\,
            I => \N__5227\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5227\,
            I => \N__5224\
        );

    \I__833\ : IoSpan4Mux
    port map (
            O => \N__5224\,
            I => \N__5221\
        );

    \I__832\ : Span4Mux_s3_v
    port map (
            O => \N__5221\,
            I => \N__5218\
        );

    \I__831\ : Sp12to4
    port map (
            O => \N__5218\,
            I => \N__5214\
        );

    \I__830\ : InMux
    port map (
            O => \N__5217\,
            I => \N__5211\
        );

    \I__829\ : Odrv12
    port map (
            O => \N__5214\,
            I => \DBDIR_c\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5211\,
            I => \DBDIR_c\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__5206\,
            I => \U712_CHIP_RAM.N_323_cascade_\
        );

    \I__826\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5200\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5200\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a2_0_0_0\
        );

    \I__824\ : InMux
    port map (
            O => \N__5197\,
            I => \N__5193\
        );

    \I__823\ : InMux
    port map (
            O => \N__5196\,
            I => \N__5190\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5193\,
            I => \N__5187\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5190\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__820\ : Odrv12
    port map (
            O => \N__5187\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__819\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5178\
        );

    \I__818\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5175\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5178\,
            I => \N__5172\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5175\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__815\ : Odrv12
    port map (
            O => \N__5172\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__814\ : InMux
    port map (
            O => \N__5167\,
            I => \N__5164\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5164\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__5161\,
            I => \U712_CHIP_RAM.N_307_cascade_\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__5158\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_cascade_\
        );

    \I__810\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5149\
        );

    \I__809\ : InMux
    port map (
            O => \N__5154\,
            I => \N__5149\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5149\,
            I => \N__5146\
        );

    \I__807\ : Span4Mux_v
    port map (
            O => \N__5146\,
            I => \N__5142\
        );

    \I__806\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5139\
        );

    \I__805\ : Span4Mux_v
    port map (
            O => \N__5142\,
            I => \N__5134\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5139\,
            I => \N__5134\
        );

    \I__803\ : Span4Mux_h
    port map (
            O => \N__5134\,
            I => \N__5131\
        );

    \I__802\ : Sp12to4
    port map (
            O => \N__5131\,
            I => \N__5128\
        );

    \I__801\ : Span12Mux_v
    port map (
            O => \N__5128\,
            I => \N__5125\
        );

    \I__800\ : Span12Mux_h
    port map (
            O => \N__5125\,
            I => \N__5122\
        );

    \I__799\ : Odrv12
    port map (
            O => \N__5122\,
            I => \CASUn_c\
        );

    \I__798\ : CascadeMux
    port map (
            O => \N__5119\,
            I => \N__5116\
        );

    \I__797\ : InMux
    port map (
            O => \N__5116\,
            I => \N__5110\
        );

    \I__796\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5110\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__5110\,
            I => \N__5106\
        );

    \I__794\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5103\
        );

    \I__793\ : Span4Mux_v
    port map (
            O => \N__5106\,
            I => \N__5100\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5103\,
            I => \N__5097\
        );

    \I__791\ : Sp12to4
    port map (
            O => \N__5100\,
            I => \N__5094\
        );

    \I__790\ : Sp12to4
    port map (
            O => \N__5097\,
            I => \N__5091\
        );

    \I__789\ : Span12Mux_h
    port map (
            O => \N__5094\,
            I => \N__5088\
        );

    \I__788\ : Span12Mux_v
    port map (
            O => \N__5091\,
            I => \N__5085\
        );

    \I__787\ : Span12Mux_v
    port map (
            O => \N__5088\,
            I => \N__5082\
        );

    \I__786\ : Span12Mux_h
    port map (
            O => \N__5085\,
            I => \N__5079\
        );

    \I__785\ : Odrv12
    port map (
            O => \N__5082\,
            I => \CASLn_c\
        );

    \I__784\ : Odrv12
    port map (
            O => \N__5079\,
            I => \CASLn_c\
        );

    \I__783\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5068\
        );

    \I__782\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5068\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5068\,
            I => \N__5065\
        );

    \I__780\ : Odrv4
    port map (
            O => \N__5065\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__779\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5058\
        );

    \I__778\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5055\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5058\,
            I => \N__5052\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__5055\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__775\ : Odrv12
    port map (
            O => \N__5052\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__774\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5043\
        );

    \I__773\ : InMux
    port map (
            O => \N__5046\,
            I => \N__5040\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5043\,
            I => \N__5036\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5040\,
            I => \N__5033\
        );

    \I__770\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5030\
        );

    \I__769\ : Odrv4
    port map (
            O => \N__5036\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__768\ : Odrv4
    port map (
            O => \N__5033\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__5030\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__766\ : InMux
    port map (
            O => \N__5023\,
            I => \N__5020\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__5020\,
            I => \N__5016\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__5019\,
            I => \N__5013\
        );

    \I__763\ : Span4Mux_v
    port map (
            O => \N__5016\,
            I => \N__5010\
        );

    \I__762\ : InMux
    port map (
            O => \N__5013\,
            I => \N__5007\
        );

    \I__761\ : Odrv4
    port map (
            O => \N__5010\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__5007\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__759\ : IoInMux
    port map (
            O => \N__5002\,
            I => \N__4999\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4999\,
            I => \N__4996\
        );

    \I__757\ : Span12Mux_s11_v
    port map (
            O => \N__4996\,
            I => \N__4993\
        );

    \I__756\ : Span12Mux_h
    port map (
            O => \N__4993\,
            I => \N__4990\
        );

    \I__755\ : Odrv12
    port map (
            O => \N__4990\,
            I => \U712_REG_SM_un1_UDSn_i\
        );

    \I__754\ : InMux
    port map (
            O => \N__4987\,
            I => \N__4980\
        );

    \I__753\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4980\
        );

    \I__752\ : InMux
    port map (
            O => \N__4985\,
            I => \N__4977\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4980\,
            I => \N__4973\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__4977\,
            I => \N__4970\
        );

    \I__749\ : InMux
    port map (
            O => \N__4976\,
            I => \N__4966\
        );

    \I__748\ : Span4Mux_v
    port map (
            O => \N__4973\,
            I => \N__4963\
        );

    \I__747\ : Span4Mux_v
    port map (
            O => \N__4970\,
            I => \N__4960\
        );

    \I__746\ : InMux
    port map (
            O => \N__4969\,
            I => \N__4957\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4966\,
            I => \N__4954\
        );

    \I__744\ : Sp12to4
    port map (
            O => \N__4963\,
            I => \N__4947\
        );

    \I__743\ : Sp12to4
    port map (
            O => \N__4960\,
            I => \N__4947\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4957\,
            I => \N__4947\
        );

    \I__741\ : Span4Mux_v
    port map (
            O => \N__4954\,
            I => \N__4944\
        );

    \I__740\ : Span12Mux_h
    port map (
            O => \N__4947\,
            I => \N__4941\
        );

    \I__739\ : Sp12to4
    port map (
            O => \N__4944\,
            I => \N__4938\
        );

    \I__738\ : Span12Mux_v
    port map (
            O => \N__4941\,
            I => \N__4935\
        );

    \I__737\ : Span12Mux_h
    port map (
            O => \N__4938\,
            I => \N__4932\
        );

    \I__736\ : Odrv12
    port map (
            O => \N__4935\,
            I => \RnW_c\
        );

    \I__735\ : Odrv12
    port map (
            O => \N__4932\,
            I => \RnW_c\
        );

    \I__734\ : IoInMux
    port map (
            O => \N__4927\,
            I => \N__4924\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4924\,
            I => \N__4921\
        );

    \I__732\ : Span4Mux_s2_h
    port map (
            O => \N__4921\,
            I => \N__4918\
        );

    \I__731\ : Sp12to4
    port map (
            O => \N__4918\,
            I => \N__4915\
        );

    \I__730\ : Span12Mux_s6_v
    port map (
            O => \N__4915\,
            I => \N__4912\
        );

    \I__729\ : Span12Mux_h
    port map (
            O => \N__4912\,
            I => \N__4909\
        );

    \I__728\ : Odrv12
    port map (
            O => \N__4909\,
            I => \DRDDIR_i_m4_i_m2\
        );

    \I__727\ : InMux
    port map (
            O => \N__4906\,
            I => \N__4902\
        );

    \I__726\ : InMux
    port map (
            O => \N__4905\,
            I => \N__4899\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4902\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__4899\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__723\ : InMux
    port map (
            O => \N__4894\,
            I => \N__4890\
        );

    \I__722\ : InMux
    port map (
            O => \N__4893\,
            I => \N__4887\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4890\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4887\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__4882\,
            I => \N__4878\
        );

    \I__718\ : InMux
    port map (
            O => \N__4881\,
            I => \N__4875\
        );

    \I__717\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4872\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4875\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4872\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__4867\,
            I => \N__4864\
        );

    \I__713\ : InMux
    port map (
            O => \N__4864\,
            I => \N__4861\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4861\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_RNOZ0Z_0\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__4858\,
            I => \N__4850\
        );

    \I__710\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4847\
        );

    \I__709\ : InMux
    port map (
            O => \N__4856\,
            I => \N__4844\
        );

    \I__708\ : CascadeMux
    port map (
            O => \N__4855\,
            I => \N__4841\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__4854\,
            I => \N__4838\
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__4853\,
            I => \N__4835\
        );

    \I__705\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4832\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__4847\,
            I => \N__4825\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4844\,
            I => \N__4825\
        );

    \I__702\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4820\
        );

    \I__701\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4820\
        );

    \I__700\ : InMux
    port map (
            O => \N__4835\,
            I => \N__4817\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__4832\,
            I => \N__4814\
        );

    \I__698\ : InMux
    port map (
            O => \N__4831\,
            I => \N__4809\
        );

    \I__697\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4809\
        );

    \I__696\ : Odrv4
    port map (
            O => \N__4825\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4820\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4817\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__693\ : Odrv4
    port map (
            O => \N__4814\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4809\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__691\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4795\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4795\,
            I => \U712_REG_SM.N_265\
        );

    \I__689\ : InMux
    port map (
            O => \N__4792\,
            I => \N__4788\
        );

    \I__688\ : InMux
    port map (
            O => \N__4791\,
            I => \N__4785\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__4788\,
            I => \U712_REG_SM.N_183\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4785\,
            I => \U712_REG_SM.N_183\
        );

    \I__685\ : InMux
    port map (
            O => \N__4780\,
            I => \N__4777\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__4777\,
            I => \N__4772\
        );

    \I__683\ : InMux
    port map (
            O => \N__4776\,
            I => \N__4769\
        );

    \I__682\ : InMux
    port map (
            O => \N__4775\,
            I => \N__4766\
        );

    \I__681\ : Odrv4
    port map (
            O => \N__4772\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__4769\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__4766\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__678\ : InMux
    port map (
            O => \N__4759\,
            I => \N__4753\
        );

    \I__677\ : InMux
    port map (
            O => \N__4758\,
            I => \N__4750\
        );

    \I__676\ : InMux
    port map (
            O => \N__4757\,
            I => \N__4747\
        );

    \I__675\ : InMux
    port map (
            O => \N__4756\,
            I => \N__4744\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__4753\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4750\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4747\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4744\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__670\ : InMux
    port map (
            O => \N__4735\,
            I => \N__4731\
        );

    \I__669\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4728\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4731\,
            I => \N__4725\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__4728\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__666\ : Odrv12
    port map (
            O => \N__4725\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__665\ : CascadeMux
    port map (
            O => \N__4720\,
            I => \N__4717\
        );

    \I__664\ : InMux
    port map (
            O => \N__4717\,
            I => \N__4713\
        );

    \I__663\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4710\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__4713\,
            I => \N__4707\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4710\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__4707\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__659\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4699\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4699\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__657\ : InMux
    port map (
            O => \N__4696\,
            I => \N__4693\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__4693\,
            I => \N__4689\
        );

    \I__655\ : InMux
    port map (
            O => \N__4692\,
            I => \N__4685\
        );

    \I__654\ : Span4Mux_h
    port map (
            O => \N__4689\,
            I => \N__4682\
        );

    \I__653\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4679\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__4685\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__651\ : Odrv4
    port map (
            O => \N__4682\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4679\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__649\ : InMux
    port map (
            O => \N__4672\,
            I => \N__4669\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4669\,
            I => \U712_CHIP_RAM.DBR_SYNCZ0Z_2\
        );

    \I__647\ : InMux
    port map (
            O => \N__4666\,
            I => \N__4662\
        );

    \I__646\ : InMux
    port map (
            O => \N__4665\,
            I => \N__4659\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4662\,
            I => \N__4656\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4659\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__643\ : Odrv4
    port map (
            O => \N__4656\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__4651\,
            I => \U712_CHIP_RAM.N_177_cascade_\
        );

    \I__641\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4645\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4645\,
            I => \N__4641\
        );

    \I__639\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4638\
        );

    \I__638\ : Odrv4
    port map (
            O => \N__4641\,
            I => \U712_CHIP_RAM.N_197\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4638\,
            I => \U712_CHIP_RAM.N_197\
        );

    \I__636\ : InMux
    port map (
            O => \N__4633\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__635\ : InMux
    port map (
            O => \N__4630\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__634\ : InMux
    port map (
            O => \N__4627\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__633\ : InMux
    port map (
            O => \N__4624\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__632\ : InMux
    port map (
            O => \N__4621\,
            I => \N__4617\
        );

    \I__631\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4614\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4617\,
            I => \N__4611\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__4614\,
            I => \N__4608\
        );

    \I__628\ : Span4Mux_v
    port map (
            O => \N__4611\,
            I => \N__4605\
        );

    \I__627\ : Span4Mux_v
    port map (
            O => \N__4608\,
            I => \N__4602\
        );

    \I__626\ : Sp12to4
    port map (
            O => \N__4605\,
            I => \N__4599\
        );

    \I__625\ : Span4Mux_h
    port map (
            O => \N__4602\,
            I => \N__4596\
        );

    \I__624\ : Span12Mux_h
    port map (
            O => \N__4599\,
            I => \N__4591\
        );

    \I__623\ : Sp12to4
    port map (
            O => \N__4596\,
            I => \N__4591\
        );

    \I__622\ : Span12Mux_v
    port map (
            O => \N__4591\,
            I => \N__4588\
        );

    \I__621\ : Odrv12
    port map (
            O => \N__4588\,
            I => \TSn_c\
        );

    \I__620\ : CascadeMux
    port map (
            O => \N__4585\,
            I => \N__4582\
        );

    \I__619\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4579\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__4579\,
            I => \N__4576\
        );

    \I__617\ : Span4Mux_v
    port map (
            O => \N__4576\,
            I => \N__4573\
        );

    \I__616\ : Sp12to4
    port map (
            O => \N__4573\,
            I => \N__4570\
        );

    \I__615\ : Span12Mux_h
    port map (
            O => \N__4570\,
            I => \N__4567\
        );

    \I__614\ : Span12Mux_v
    port map (
            O => \N__4567\,
            I => \N__4564\
        );

    \I__613\ : Odrv12
    port map (
            O => \N__4564\,
            I => \RAMSPACEn_c\
        );

    \I__612\ : InMux
    port map (
            O => \N__4561\,
            I => \N__4557\
        );

    \I__611\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4552\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4557\,
            I => \N__4549\
        );

    \I__609\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4546\
        );

    \I__608\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4543\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__4552\,
            I => \N__4540\
        );

    \I__606\ : Odrv4
    port map (
            O => \N__4549\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4546\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4543\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__603\ : Odrv12
    port map (
            O => \N__4540\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__602\ : InMux
    port map (
            O => \N__4531\,
            I => \N__4527\
        );

    \I__601\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4524\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__4527\,
            I => \N__4519\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4524\,
            I => \N__4519\
        );

    \I__598\ : Odrv4
    port map (
            O => \N__4519\,
            I => \U712_REG_SM.N_325\
        );

    \I__597\ : InMux
    port map (
            O => \N__4516\,
            I => \N__4512\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__4515\,
            I => \N__4509\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4512\,
            I => \N__4505\
        );

    \I__594\ : InMux
    port map (
            O => \N__4509\,
            I => \N__4502\
        );

    \I__593\ : InMux
    port map (
            O => \N__4508\,
            I => \N__4496\
        );

    \I__592\ : Span4Mux_h
    port map (
            O => \N__4505\,
            I => \N__4493\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4502\,
            I => \N__4490\
        );

    \I__590\ : InMux
    port map (
            O => \N__4501\,
            I => \N__4487\
        );

    \I__589\ : InMux
    port map (
            O => \N__4500\,
            I => \N__4482\
        );

    \I__588\ : InMux
    port map (
            O => \N__4499\,
            I => \N__4482\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4496\,
            I => \U712_REG_SM.N_201\
        );

    \I__586\ : Odrv4
    port map (
            O => \N__4493\,
            I => \U712_REG_SM.N_201\
        );

    \I__585\ : Odrv4
    port map (
            O => \N__4490\,
            I => \U712_REG_SM.N_201\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4487\,
            I => \U712_REG_SM.N_201\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__4482\,
            I => \U712_REG_SM.N_201\
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__4471\,
            I => \N__4468\
        );

    \I__581\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4463\
        );

    \I__580\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4460\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__4466\,
            I => \N__4457\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__4463\,
            I => \N__4452\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__4460\,
            I => \N__4452\
        );

    \I__576\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4449\
        );

    \I__575\ : Span4Mux_v
    port map (
            O => \N__4452\,
            I => \N__4446\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4449\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__573\ : Odrv4
    port map (
            O => \N__4446\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__572\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4437\
        );

    \I__571\ : IoInMux
    port map (
            O => \N__4440\,
            I => \N__4434\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4437\,
            I => \N__4431\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__4434\,
            I => \N__4428\
        );

    \I__568\ : Span4Mux_v
    port map (
            O => \N__4431\,
            I => \N__4425\
        );

    \I__567\ : IoSpan4Mux
    port map (
            O => \N__4428\,
            I => \N__4422\
        );

    \I__566\ : Sp12to4
    port map (
            O => \N__4425\,
            I => \N__4419\
        );

    \I__565\ : IoSpan4Mux
    port map (
            O => \N__4422\,
            I => \N__4416\
        );

    \I__564\ : Span12Mux_h
    port map (
            O => \N__4419\,
            I => \N__4413\
        );

    \I__563\ : IoSpan4Mux
    port map (
            O => \N__4416\,
            I => \N__4410\
        );

    \I__562\ : Odrv12
    port map (
            O => \N__4413\,
            I => \C3_c\
        );

    \I__561\ : Odrv4
    port map (
            O => \N__4410\,
            I => \C3_c\
        );

    \I__560\ : InMux
    port map (
            O => \N__4405\,
            I => \N__4400\
        );

    \I__559\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4394\
        );

    \I__558\ : InMux
    port map (
            O => \N__4403\,
            I => \N__4394\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__4400\,
            I => \N__4391\
        );

    \I__556\ : InMux
    port map (
            O => \N__4399\,
            I => \N__4388\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4394\,
            I => \N__4385\
        );

    \I__554\ : Odrv12
    port map (
            O => \N__4391\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__4388\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__552\ : Odrv4
    port map (
            O => \N__4385\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__4378\,
            I => \N__4374\
        );

    \I__550\ : InMux
    port map (
            O => \N__4377\,
            I => \N__4371\
        );

    \I__549\ : InMux
    port map (
            O => \N__4374\,
            I => \N__4368\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4371\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4368\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__546\ : IoInMux
    port map (
            O => \N__4363\,
            I => \N__4360\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__4360\,
            I => \N__4357\
        );

    \I__544\ : IoSpan4Mux
    port map (
            O => \N__4357\,
            I => \N__4354\
        );

    \I__543\ : IoSpan4Mux
    port map (
            O => \N__4354\,
            I => \N__4351\
        );

    \I__542\ : Span4Mux_s0_v
    port map (
            O => \N__4351\,
            I => \N__4348\
        );

    \I__541\ : Sp12to4
    port map (
            O => \N__4348\,
            I => \N__4345\
        );

    \I__540\ : Span12Mux_v
    port map (
            O => \N__4345\,
            I => \N__4342\
        );

    \I__539\ : Odrv12
    port map (
            O => \N__4342\,
            I => \U712_REG_SM_un1_LDSn_i\
        );

    \I__538\ : InMux
    port map (
            O => \N__4339\,
            I => \N__4333\
        );

    \I__537\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4333\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4333\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0\
        );

    \I__535\ : InMux
    port map (
            O => \N__4330\,
            I => \bfn_9_9_0_\
        );

    \I__534\ : InMux
    port map (
            O => \N__4327\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__533\ : InMux
    port map (
            O => \N__4324\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__532\ : InMux
    port map (
            O => \N__4321\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__4318\,
            I => \U712_REG_SM.N_215_cascade_\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__4315\,
            I => \U712_REG_SM.N_200_cascade_\
        );

    \I__529\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4308\
        );

    \I__528\ : InMux
    port map (
            O => \N__4311\,
            I => \N__4305\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4308\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4305\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__525\ : InMux
    port map (
            O => \N__4300\,
            I => \N__4296\
        );

    \I__524\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4293\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4296\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4293\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__521\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4281\
        );

    \I__520\ : InMux
    port map (
            O => \N__4287\,
            I => \N__4281\
        );

    \I__519\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4278\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4281\,
            I => \U712_REG_SM.N_200\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4278\,
            I => \U712_REG_SM.N_200\
        );

    \I__516\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4269\
        );

    \I__515\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4266\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__4269\,
            I => \U712_REG_SM.N_219\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4266\,
            I => \U712_REG_SM.N_219\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__4261\,
            I => \U712_REG_SM.N_325_cascade_\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__4258\,
            I => \N__4249\
        );

    \I__510\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4246\
        );

    \I__509\ : InMux
    port map (
            O => \N__4256\,
            I => \N__4241\
        );

    \I__508\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4241\
        );

    \I__507\ : InMux
    port map (
            O => \N__4254\,
            I => \N__4238\
        );

    \I__506\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4231\
        );

    \I__505\ : InMux
    port map (
            O => \N__4252\,
            I => \N__4231\
        );

    \I__504\ : InMux
    port map (
            O => \N__4249\,
            I => \N__4231\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4246\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4241\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__4238\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4231\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__499\ : InMux
    port map (
            O => \N__4222\,
            I => \N__4219\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4219\,
            I => \N__4216\
        );

    \I__497\ : Odrv4
    port map (
            O => \N__4216\,
            I => \U712_REG_SM.N_198\
        );

    \I__496\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4210\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4210\,
            I => \N__4205\
        );

    \I__494\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4202\
        );

    \I__493\ : InMux
    port map (
            O => \N__4208\,
            I => \N__4199\
        );

    \I__492\ : Odrv4
    port map (
            O => \N__4205\,
            I => \U712_REG_SM.N_212\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4202\,
            I => \U712_REG_SM.N_212\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4199\,
            I => \U712_REG_SM.N_212\
        );

    \I__489\ : InMux
    port map (
            O => \N__4192\,
            I => \N__4187\
        );

    \I__488\ : InMux
    port map (
            O => \N__4191\,
            I => \N__4184\
        );

    \I__487\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4181\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__4187\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__4184\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4181\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__4174\,
            I => \U712_REG_SM.N_198_cascade_\
        );

    \I__482\ : CascadeMux
    port map (
            O => \N__4171\,
            I => \U712_REG_SM.DS_EN_RNOZ0Z_0_cascade_\
        );

    \I__481\ : CascadeMux
    port map (
            O => \N__4168\,
            I => \U712_BYTE_ENABLE.N_271_cascade_\
        );

    \I__480\ : IoInMux
    port map (
            O => \N__4165\,
            I => \N__4162\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4162\,
            I => \N__4159\
        );

    \I__478\ : Span4Mux_s3_h
    port map (
            O => \N__4159\,
            I => \N__4156\
        );

    \I__477\ : Span4Mux_v
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__476\ : Sp12to4
    port map (
            O => \N__4153\,
            I => \N__4150\
        );

    \I__475\ : Span12Mux_s11_h
    port map (
            O => \N__4150\,
            I => \N__4147\
        );

    \I__474\ : Odrv12
    port map (
            O => \N__4147\,
            I => \N_44_i\
        );

    \I__473\ : InMux
    port map (
            O => \N__4144\,
            I => \N__4135\
        );

    \I__472\ : InMux
    port map (
            O => \N__4143\,
            I => \N__4135\
        );

    \I__471\ : InMux
    port map (
            O => \N__4142\,
            I => \N__4135\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4135\,
            I => \N__4131\
        );

    \I__469\ : InMux
    port map (
            O => \N__4134\,
            I => \N__4128\
        );

    \I__468\ : Span4Mux_h
    port map (
            O => \N__4131\,
            I => \N__4121\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4128\,
            I => \N__4121\
        );

    \I__466\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4118\
        );

    \I__465\ : InMux
    port map (
            O => \N__4126\,
            I => \N__4115\
        );

    \I__464\ : Span4Mux_v
    port map (
            O => \N__4121\,
            I => \N__4110\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4118\,
            I => \N__4110\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4115\,
            I => \N__4107\
        );

    \I__461\ : Span4Mux_v
    port map (
            O => \N__4110\,
            I => \N__4104\
        );

    \I__460\ : Span12Mux_v
    port map (
            O => \N__4107\,
            I => \N__4099\
        );

    \I__459\ : Sp12to4
    port map (
            O => \N__4104\,
            I => \N__4099\
        );

    \I__458\ : Odrv12
    port map (
            O => \N__4099\,
            I => \A_c_0\
        );

    \I__457\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4086\
        );

    \I__456\ : InMux
    port map (
            O => \N__4095\,
            I => \N__4086\
        );

    \I__455\ : InMux
    port map (
            O => \N__4094\,
            I => \N__4086\
        );

    \I__454\ : InMux
    port map (
            O => \N__4093\,
            I => \N__4083\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__4086\,
            I => \N__4078\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4083\,
            I => \N__4078\
        );

    \I__451\ : Span12Mux_v
    port map (
            O => \N__4078\,
            I => \N__4075\
        );

    \I__450\ : Odrv12
    port map (
            O => \N__4075\,
            I => \A_c_1\
        );

    \I__449\ : InMux
    port map (
            O => \N__4072\,
            I => \N__4069\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4069\,
            I => \U712_BYTE_ENABLE.N_277\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__4066\,
            I => \N__4063\
        );

    \I__446\ : InMux
    port map (
            O => \N__4063\,
            I => \N__4059\
        );

    \I__445\ : CascadeMux
    port map (
            O => \N__4062\,
            I => \N__4056\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__4059\,
            I => \N__4052\
        );

    \I__443\ : InMux
    port map (
            O => \N__4056\,
            I => \N__4047\
        );

    \I__442\ : InMux
    port map (
            O => \N__4055\,
            I => \N__4047\
        );

    \I__441\ : Span4Mux_h
    port map (
            O => \N__4052\,
            I => \N__4042\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4047\,
            I => \N__4042\
        );

    \I__439\ : Span4Mux_v
    port map (
            O => \N__4042\,
            I => \N__4039\
        );

    \I__438\ : Sp12to4
    port map (
            O => \N__4039\,
            I => \N__4036\
        );

    \I__437\ : Span12Mux_h
    port map (
            O => \N__4036\,
            I => \N__4033\
        );

    \I__436\ : Span12Mux_v
    port map (
            O => \N__4033\,
            I => \N__4030\
        );

    \I__435\ : Odrv12
    port map (
            O => \N__4030\,
            I => \SIZ_c_1\
        );

    \I__434\ : InMux
    port map (
            O => \N__4027\,
            I => \N__4024\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__4024\,
            I => \N__4019\
        );

    \I__432\ : InMux
    port map (
            O => \N__4023\,
            I => \N__4016\
        );

    \I__431\ : InMux
    port map (
            O => \N__4022\,
            I => \N__4013\
        );

    \I__430\ : Span4Mux_v
    port map (
            O => \N__4019\,
            I => \N__4006\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4016\,
            I => \N__4006\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__4013\,
            I => \N__4006\
        );

    \I__427\ : Sp12to4
    port map (
            O => \N__4006\,
            I => \N__4003\
        );

    \I__426\ : Span12Mux_v
    port map (
            O => \N__4003\,
            I => \N__4000\
        );

    \I__425\ : Odrv12
    port map (
            O => \N__4000\,
            I => \SIZ_c_0\
        );

    \I__424\ : InMux
    port map (
            O => \N__3997\,
            I => \N__3985\
        );

    \I__423\ : InMux
    port map (
            O => \N__3996\,
            I => \N__3985\
        );

    \I__422\ : InMux
    port map (
            O => \N__3995\,
            I => \N__3985\
        );

    \I__421\ : InMux
    port map (
            O => \N__3994\,
            I => \N__3985\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3985\,
            I => \U712_BYTE_ENABLE.N_270\
        );

    \I__419\ : IoInMux
    port map (
            O => \N__3982\,
            I => \N__3979\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3979\,
            I => \N__3975\
        );

    \I__417\ : IoInMux
    port map (
            O => \N__3978\,
            I => \N__3972\
        );

    \I__416\ : Span4Mux_s0_v
    port map (
            O => \N__3975\,
            I => \N__3969\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3972\,
            I => \N__3966\
        );

    \I__414\ : Span4Mux_h
    port map (
            O => \N__3969\,
            I => \N__3963\
        );

    \I__413\ : Span4Mux_s0_v
    port map (
            O => \N__3966\,
            I => \N__3960\
        );

    \I__412\ : Sp12to4
    port map (
            O => \N__3963\,
            I => \N__3957\
        );

    \I__411\ : Sp12to4
    port map (
            O => \N__3960\,
            I => \N__3954\
        );

    \I__410\ : Span12Mux_h
    port map (
            O => \N__3957\,
            I => \N__3949\
        );

    \I__409\ : Span12Mux_s11_h
    port map (
            O => \N__3954\,
            I => \N__3949\
        );

    \I__408\ : Span12Mux_v
    port map (
            O => \N__3949\,
            I => \N__3945\
        );

    \I__407\ : InMux
    port map (
            O => \N__3948\,
            I => \N__3942\
        );

    \I__406\ : Odrv12
    port map (
            O => \N__3945\,
            I => \ASn_c\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__3942\,
            I => \ASn_c\
        );

    \I__404\ : CascadeMux
    port map (
            O => \N__3937\,
            I => \U712_REG_SM.N_266_cascade_\
        );

    \I__403\ : InMux
    port map (
            O => \N__3934\,
            I => \N__3931\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3931\,
            I => \U712_REG_SM.N_215\
        );

    \I__401\ : IoInMux
    port map (
            O => \N__3928\,
            I => \N__3925\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3925\,
            I => \N__3922\
        );

    \I__399\ : IoSpan4Mux
    port map (
            O => \N__3922\,
            I => \N__3919\
        );

    \I__398\ : Span4Mux_s2_h
    port map (
            O => \N__3919\,
            I => \N__3916\
        );

    \I__397\ : Span4Mux_h
    port map (
            O => \N__3916\,
            I => \N__3913\
        );

    \I__396\ : Span4Mux_h
    port map (
            O => \N__3913\,
            I => \N__3910\
        );

    \I__395\ : Odrv4
    port map (
            O => \N__3910\,
            I => \N_944_i\
        );

    \I__394\ : IoInMux
    port map (
            O => \N__3907\,
            I => \N__3904\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3904\,
            I => \N__3901\
        );

    \I__392\ : Span12Mux_s5_v
    port map (
            O => \N__3901\,
            I => \N__3898\
        );

    \I__391\ : Odrv12
    port map (
            O => \N__3898\,
            I => \VBENn_c\
        );

    \I__390\ : CascadeMux
    port map (
            O => \N__3895\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_cascade_\
        );

    \I__389\ : IoInMux
    port map (
            O => \N__3892\,
            I => \N__3889\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3889\,
            I => \N__3886\
        );

    \I__387\ : Span12Mux_s11_v
    port map (
            O => \N__3886\,
            I => \N__3883\
        );

    \I__386\ : Odrv12
    port map (
            O => \N__3883\,
            I => \N_41_i\
        );

    \I__385\ : InMux
    port map (
            O => \N__3880\,
            I => \N__3877\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3877\,
            I => \N__3874\
        );

    \I__383\ : Odrv4
    port map (
            O => \N__3874\,
            I => \U712_BYTE_ENABLE.N_273\
        );

    \I__382\ : IoInMux
    port map (
            O => \N__3871\,
            I => \N__3868\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__3868\,
            I => \N__3865\
        );

    \I__380\ : Span12Mux_s8_h
    port map (
            O => \N__3865\,
            I => \N__3862\
        );

    \I__379\ : Span12Mux_h
    port map (
            O => \N__3862\,
            I => \N__3859\
        );

    \I__378\ : Span12Mux_v
    port map (
            O => \N__3859\,
            I => \N__3856\
        );

    \I__377\ : Odrv12
    port map (
            O => \N__3856\,
            I => \N_43_i\
        );

    \I__376\ : InMux
    port map (
            O => \N__3853\,
            I => \N__3850\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__3850\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0\
        );

    \I__374\ : CascadeMux
    port map (
            O => \N__3847\,
            I => \U712_BYTE_ENABLE.N_275_cascade_\
        );

    \I__373\ : IoInMux
    port map (
            O => \N__3844\,
            I => \N__3841\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3841\,
            I => \N__3838\
        );

    \I__371\ : Span12Mux_s5_h
    port map (
            O => \N__3838\,
            I => \N__3835\
        );

    \I__370\ : Span12Mux_h
    port map (
            O => \N__3835\,
            I => \N__3832\
        );

    \I__369\ : Span12Mux_v
    port map (
            O => \N__3832\,
            I => \N__3829\
        );

    \I__368\ : Odrv12
    port map (
            O => \N__3829\,
            I => \N_42_i\
        );

    \I__367\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3822\
        );

    \I__366\ : InMux
    port map (
            O => \N__3825\,
            I => \N__3819\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__3822\,
            I => \U712_REG_SM.REG_CYCLE_GOZ0\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3819\,
            I => \U712_REG_SM.REG_CYCLE_GOZ0\
        );

    \I__363\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3811\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__3811\,
            I => \U712_REG_SM.UDS_OUT_2_0_a2_0_a3_0\
        );

    \I__361\ : InMux
    port map (
            O => \N__3808\,
            I => \N__3805\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3805\,
            I => \N__3801\
        );

    \I__359\ : IoInMux
    port map (
            O => \N__3804\,
            I => \N__3798\
        );

    \I__358\ : Span4Mux_h
    port map (
            O => \N__3801\,
            I => \N__3795\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__3798\,
            I => \N__3792\
        );

    \I__356\ : Span4Mux_h
    port map (
            O => \N__3795\,
            I => \N__3787\
        );

    \I__355\ : Span4Mux_s3_h
    port map (
            O => \N__3792\,
            I => \N__3787\
        );

    \I__354\ : Sp12to4
    port map (
            O => \N__3787\,
            I => \N__3784\
        );

    \I__353\ : Span12Mux_v
    port map (
            O => \N__3784\,
            I => \N__3781\
        );

    \I__352\ : Odrv12
    port map (
            O => \N__3781\,
            I => \C1_c\
        );

    \I__351\ : CascadeMux
    port map (
            O => \N__3778\,
            I => \U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1_cascade_\
        );

    \I__350\ : InMux
    port map (
            O => \N__3775\,
            I => \N__3769\
        );

    \I__349\ : InMux
    port map (
            O => \N__3774\,
            I => \N__3769\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3769\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__347\ : InMux
    port map (
            O => \N__3766\,
            I => \N__3763\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__3763\,
            I => \U712_REG_SM.LDS_OUT_2_0_a2_0_a3_0\
        );

    \I__345\ : InMux
    port map (
            O => \N__3760\,
            I => \N__3750\
        );

    \I__344\ : InMux
    port map (
            O => \N__3759\,
            I => \N__3750\
        );

    \I__343\ : InMux
    port map (
            O => \N__3758\,
            I => \N__3750\
        );

    \I__342\ : InMux
    port map (
            O => \N__3757\,
            I => \N__3747\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__3750\,
            I => \N__3744\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__3747\,
            I => \U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1\
        );

    \I__339\ : Odrv4
    port map (
            O => \N__3744\,
            I => \U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1\
        );

    \I__338\ : IoInMux
    port map (
            O => \N__3739\,
            I => \N__3736\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__3736\,
            I => \N__3733\
        );

    \I__336\ : Span4Mux_s2_v
    port map (
            O => \N__3733\,
            I => \N__3730\
        );

    \I__335\ : Span4Mux_v
    port map (
            O => \N__3730\,
            I => \N__3727\
        );

    \I__334\ : Odrv4
    port map (
            O => \N__3727\,
            I => \CLK80_OUT_i_i\
        );

    \I__333\ : IoInMux
    port map (
            O => \N__3724\,
            I => \N__3721\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__3721\,
            I => \N__3718\
        );

    \I__331\ : Odrv12
    port map (
            O => \N__3718\,
            I => \CLK40_OUT_i_i\
        );

    \I__330\ : CascadeMux
    port map (
            O => \N__3715\,
            I => \N__3712\
        );

    \I__329\ : InMux
    port map (
            O => \N__3712\,
            I => \N__3709\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__3709\,
            I => \N__3706\
        );

    \I__327\ : Span4Mux_v
    port map (
            O => \N__3706\,
            I => \N__3703\
        );

    \I__326\ : Span4Mux_h
    port map (
            O => \N__3703\,
            I => \N__3700\
        );

    \I__325\ : Sp12to4
    port map (
            O => \N__3700\,
            I => \N__3697\
        );

    \I__324\ : Span12Mux_v
    port map (
            O => \N__3697\,
            I => \N__3694\
        );

    \I__323\ : Odrv12
    port map (
            O => \N__3694\,
            I => \REGSPACEn_c\
        );

    \I__322\ : IoInMux
    port map (
            O => \N__3691\,
            I => \N__3688\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__3688\,
            I => \N__3685\
        );

    \I__320\ : IoSpan4Mux
    port map (
            O => \N__3685\,
            I => \N__3682\
        );

    \I__319\ : Span4Mux_s2_v
    port map (
            O => \N__3682\,
            I => \N__3679\
        );

    \I__318\ : Sp12to4
    port map (
            O => \N__3679\,
            I => \N__3676\
        );

    \I__317\ : Span12Mux_v
    port map (
            O => \N__3676\,
            I => \N__3673\
        );

    \I__316\ : Odrv12
    port map (
            O => \N__3673\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__9309\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_8C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_8C_net\,
            I => \N__9307\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__9308\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__9304\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__9305\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__9306\
        );

    \IN_MUX_bfv_10_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_14_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7771\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3804\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4440\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_3_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8788\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK40C_obuf_RNO_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8074\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_RNO_0_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__4985\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4134\,
            lcout => \U712_REG_SM.UDS_OUT_2_0_a2_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDS_OUT_RNO_0_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4969\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4127\,
            lcout => \U712_REG_SM.LDS_OUT_2_0_a2_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001101"
        )
    port map (
            in0 => \N__4620\,
            in1 => \N__4555\,
            in2 => \N__3715\,
            in3 => \N__3826\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8772\,
            ce => 'H',
            sr => \N__9496\
        );

    \U712_REG_SM.C3_SYNC_2_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4759\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => 'H',
            sr => \N__9490\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__3759\,
            in1 => \N__4191\,
            in2 => \_gnd_net_\,
            in3 => \N__4213\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => 'H',
            sr => \N__9490\
        );

    \U712_REG_SM.C1_SYNC_2_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4257\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => 'H',
            sr => \N__9490\
        );

    \U712_REG_SM.REG_CYCLE_GO_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__3758\,
            in1 => \N__4556\,
            in2 => \N__4471\,
            in3 => \N__3825\,
            lcout => \U712_REG_SM.REG_CYCLE_GOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => 'H',
            sr => \N__9490\
        );

    \U712_REG_SM.UDS_OUT_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001110111"
        )
    port map (
            in0 => \N__4023\,
            in1 => \N__3814\,
            in2 => \N__5019\,
            in3 => \N__3760\,
            lcout => \U712_REG_SM.UDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => 'H',
            sr => \N__9490\
        );

    \U712_REG_SM.C1_SYNC_1_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4857\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => 'H',
            sr => \N__9490\
        );

    \U712_REG_SM.C1_SYNC_0_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3808\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8777\,
            ce => 'H',
            sr => \N__9490\
        );

    \U712_REG_SM.C1_SYNC_RNITQLC2_1_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4273\,
            in1 => \N__4254\,
            in2 => \N__4853\,
            in3 => \N__4501\,
            lcout => \U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1\,
            ltout => \U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__4467\,
            in1 => \N__4561\,
            in2 => \N__3778\,
            in3 => \N__3775\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8780\,
            ce => 'H',
            sr => \N__9483\
        );

    \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__3774\,
            in1 => \N__4776\,
            in2 => \_gnd_net_\,
            in3 => \N__4757\,
            lcout => \U712_REG_SM.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4399\,
            in2 => \_gnd_net_\,
            in3 => \N__4312\,
            lcout => \U712_REG_SM.N_201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDS_OUT_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001110111"
        )
    port map (
            in0 => \N__3766\,
            in1 => \N__4022\,
            in2 => \N__4378\,
            in3 => \N__3757\,
            lcout => \U712_REG_SM.LDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8784\,
            ce => 'H',
            sr => \N__9472\
        );

    \TACKn_obuft_RNO_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5728\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_944_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_0_a3_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8420\,
            in2 => \_gnd_net_\,
            in3 => \N__7683\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__4095\,
            in1 => \N__4143\,
            in2 => \N__4066\,
            in3 => \N__8389\,
            lcout => \U712_BYTE_ENABLE.N_273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5874\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7733\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0\,
            ltout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_41_i_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__4072\,
            in1 => \N__3994\,
            in2 => \N__3895\,
            in3 => \N__5115\,
            lcout => \N_41_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_43_i_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__3996\,
            in1 => \N__3880\,
            in2 => \N__5119\,
            in3 => \N__4338\,
            lcout => \N_43_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4094\,
            in1 => \N__4142\,
            in2 => \_gnd_net_\,
            in3 => \N__8388\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_275_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_42_i_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__3995\,
            in1 => \N__3853\,
            in2 => \N__3847\,
            in3 => \N__5154\,
            lcout => \N_42_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_0_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4096\,
            in1 => \N__4144\,
            in2 => \_gnd_net_\,
            in3 => \N__8390\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_271_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_44_i_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__3997\,
            in1 => \N__4339\,
            in2 => \N__4168\,
            in3 => \N__5155\,
            lcout => \N_44_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__4126\,
            in1 => \N__4093\,
            in2 => \N__8419\,
            in3 => \N__4055\,
            lcout => \U712_BYTE_ENABLE.N_277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8387\,
            in2 => \N__4062\,
            in3 => \N__4027\,
            lcout => \U712_BYTE_ENABLE.N_270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000000010"
        )
    port map (
            in0 => \N__5310\,
            in1 => \N__5293\,
            in2 => \N__7407\,
            in3 => \N__7374\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8768\,
            ce => 'H',
            sr => \N__9491\
        );

    \U712_REG_SM.REGENn_1_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__4531\,
            in1 => \N__3948\,
            in2 => \N__4515\,
            in3 => \N__4222\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8768\,
            ce => 'H',
            sr => \N__9491\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001000000000"
        )
    port map (
            in0 => \N__4192\,
            in1 => \N__4209\,
            in2 => \N__5314\,
            in3 => \N__5292\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8768\,
            ce => 'H',
            sr => \N__9491\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4256\,
            in1 => \N__4500\,
            in2 => \N__4855\,
            in3 => \N__4288\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_266_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100000010"
        )
    port map (
            in0 => \N__7336\,
            in1 => \N__3934\,
            in2 => \N__3937\,
            in3 => \N__4300\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8773\,
            ce => 'H',
            sr => \N__9484\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4255\,
            in1 => \N__4499\,
            in2 => \N__4854\,
            in3 => \N__4287\,
            lcout => \U712_REG_SM.N_215\,
            ltout => \U712_REG_SM.N_215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100000"
        )
    port map (
            in0 => \N__7337\,
            in1 => \N__7403\,
            in2 => \N__4318\,
            in3 => \N__7373\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8773\,
            ce => 'H',
            sr => \N__9484\
        );

    \U712_REG_SM.C3_SYNC_1_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4405\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8773\,
            ce => 'H',
            sr => \N__9484\
        );

    \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4775\,
            in2 => \_gnd_net_\,
            in3 => \N__4756\,
            lcout => \U712_REG_SM.N_200\,
            ltout => \U712_REG_SM.N_200_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4792\,
            in2 => \N__4315\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.N_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4311\,
            in1 => \N__4830\,
            in2 => \N__4258\,
            in3 => \N__4403\,
            lcout => \U712_REG_SM.N_183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4252\,
            in1 => \N__4299\,
            in2 => \N__4858\,
            in3 => \N__4286\,
            lcout => \U712_REG_SM.N_325\,
            ltout => \U712_REG_SM.N_325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIJS6A3_1_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__4831\,
            in1 => \N__4272\,
            in2 => \N__4261\,
            in3 => \N__4253\,
            lcout => \U712_REG_SM.N_198\,
            ltout => \U712_REG_SM.N_198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__4208\,
            in1 => \N__4190\,
            in2 => \N__4174\,
            in3 => \N__4508\,
            lcout => OPEN,
            ltout => \U712_REG_SM.DS_EN_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__4404\,
            in1 => \N__5039\,
            in2 => \N__4171\,
            in3 => \N__4798\,
            lcout => \U712_REG_SM.DS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8778\,
            ce => 'H',
            sr => \N__9473\
        );

    \U712_CHIP_RAM.DBR_SYNC_2_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4692\,
            lcout => \U712_CHIP_RAM.DBR_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8781\,
            ce => 'H',
            sr => \N__9468\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5061\,
            lcout => \U712_REG_SM_DBR_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8781\,
            ce => 'H',
            sr => \N__9468\
        );

    \U712_REG_SM.C3_SYNC_0_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4441\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8781\,
            ce => 'H',
            sr => \N__9468\
        );

    \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5046\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4377\,
            lcout => \U712_REG_SM_un1_LDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7732\,
            in2 => \_gnd_net_\,
            in3 => \N__5873\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4906\,
            in2 => \_gnd_net_\,
            in3 => \N__4330\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__9303\,
            ce => 'H',
            sr => \N__5323\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5383\,
            in2 => \_gnd_net_\,
            in3 => \N__4327\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__9303\,
            ce => 'H',
            sr => \N__5323\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4894\,
            in2 => \_gnd_net_\,
            in3 => \N__4324\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__9303\,
            ce => 'H',
            sr => \N__5323\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4734\,
            in2 => \_gnd_net_\,
            in3 => \N__4321\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__9303\,
            ce => 'H',
            sr => \N__5323\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4881\,
            in2 => \_gnd_net_\,
            in3 => \N__4633\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__9303\,
            ce => 'H',
            sr => \N__5323\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5181\,
            in2 => \_gnd_net_\,
            in3 => \N__4630\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__9303\,
            ce => 'H',
            sr => \N__5323\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5196\,
            in2 => \_gnd_net_\,
            in3 => \N__4627\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__9303\,
            ce => 'H',
            sr => \N__5323\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4716\,
            in2 => \_gnd_net_\,
            in3 => \N__4624\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9303\,
            ce => 'H',
            sr => \N__5323\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100000011"
        )
    port map (
            in0 => \N__8330\,
            in1 => \N__4621\,
            in2 => \N__4585\,
            in3 => \N__4665\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8764\,
            ce => 'H',
            sr => \N__9485\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__4560\,
            in1 => \N__4530\,
            in2 => \N__4466\,
            in3 => \N__4516\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8764\,
            ce => 'H',
            sr => \N__9485\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__5506\,
            in1 => \N__6066\,
            in2 => \N__4867\,
            in3 => \N__4648\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8764\,
            ce => 'H',
            sr => \N__9485\
        );

    \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__4696\,
            in1 => \N__7369\,
            in2 => \_gnd_net_\,
            in3 => \N__5062\,
            lcout => \U712_REG_SM.N_209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7537\,
            in1 => \N__7047\,
            in2 => \N__6016\,
            in3 => \N__6634\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8769\,
            ce => \N__5458\,
            sr => \N__9474\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4986\,
            in1 => \N__5267\,
            in2 => \_gnd_net_\,
            in3 => \N__6678\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4987\,
            in2 => \_gnd_net_\,
            in3 => \N__4856\,
            lcout => \U712_REG_SM.N_265\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__4791\,
            in1 => \N__4780\,
            in2 => \_gnd_net_\,
            in3 => \N__4758\,
            lcout => \U712_REG_SM.N_187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111111011"
        )
    port map (
            in0 => \N__4735\,
            in1 => \N__5167\,
            in2 => \N__4720\,
            in3 => \N__5371\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8774\,
            ce => 'H',
            sr => \N__9469\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001010"
        )
    port map (
            in0 => \N__6677\,
            in1 => \N__5073\,
            in2 => \N__7739\,
            in3 => \N__4702\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8774\,
            ce => 'H',
            sr => \N__9469\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5074\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8774\,
            ce => 'H',
            sr => \N__9469\
        );

    \U712_CHIP_RAM.DBR_SYNC_RNIMGL61_2_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__4688\,
            in1 => \N__4672\,
            in2 => \_gnd_net_\,
            in3 => \N__4666\,
            lcout => \U712_CHIP_RAM.N_177\,
            ltout => \U712_CHIP_RAM.N_177_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIH3B52_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5427\,
            in2 => \N__4651\,
            in3 => \N__6676\,
            lcout => \U712_CHIP_RAM.N_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5444\,
            in2 => \_gnd_net_\,
            in3 => \N__4644\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a3_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5197\,
            in2 => \_gnd_net_\,
            in3 => \N__5182\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIRILU_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5426\,
            in2 => \_gnd_net_\,
            in3 => \N__6673\,
            lcout => \U712_CHIP_RAM.N_307\,
            ltout => \U712_CHIP_RAM.N_307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNI6A2O6_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5443\,
            in1 => \N__5488\,
            in2 => \N__5161\,
            in3 => \N__7218\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNI6A2O6_0_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5158\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5145\,
            in2 => \_gnd_net_\,
            in3 => \N__5109\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8782\,
            ce => 'H',
            sr => \N__9451\
        );

    \U712_CHIP_RAM.DBR_SYNC_0_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9275\,
            lcout => \U712_REG_SM_DBR_SYNC_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8782\,
            ce => 'H',
            sr => \N__9451\
        );

    \U712_REG_SM.UDS_OUT_RNIUP9B_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5047\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5023\,
            lcout => \U712_REG_SM_un1_UDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_i_m4_i_m2_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__4976\,
            in1 => \N__5268\,
            in2 => \_gnd_net_\,
            in3 => \N__7746\,
            lcout => \DRDDIR_i_m4_i_m2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100111111"
        )
    port map (
            in0 => \N__4905\,
            in1 => \N__4893\,
            in2 => \N__4882\,
            in3 => \N__5382\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5359\,
            in1 => \N__5344\,
            in2 => \_gnd_net_\,
            in3 => \N__8546\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8547\,
            in1 => \N__8400\,
            in2 => \N__5326\,
            in3 => \N__8200\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6235\,
            in1 => \N__9025\,
            in2 => \N__6203\,
            in3 => \N__8545\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101110"
        )
    port map (
            in0 => \N__5309\,
            in1 => \N__7670\,
            in2 => \N__7348\,
            in3 => \N__5291\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8761\,
            ce => 'H',
            sr => \N__9475\
        );

    \U712_CHIP_RAM.DBDIR_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__5278\,
            in1 => \N__5217\,
            in2 => \_gnd_net_\,
            in3 => \N__5910\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8761\,
            ce => 'H',
            sr => \N__9475\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI7MG83_3_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6885\,
            in1 => \N__7524\,
            in2 => \N__7977\,
            in3 => \N__6001\,
            lcout => \U712_CHIP_RAM.N_323\,
            ltout => \U712_CHIP_RAM.N_323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISS7R7_3_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__6002\,
            in1 => \N__5203\,
            in2 => \N__5206\,
            in3 => \N__5446\,
            lcout => \U712_CHIP_RAM.N_238\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000001000"
        )
    port map (
            in0 => \N__7041\,
            in1 => \N__7523\,
            in2 => \N__6898\,
            in3 => \N__7960\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_4_0_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7961\,
            in1 => \N__7042\,
            in2 => \N__6900\,
            in3 => \N__6062\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a3_3_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5445\,
            in1 => \N__6003\,
            in2 => \N__5467\,
            in3 => \N__7525\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__6004\,
            in1 => \N__6595\,
            in2 => \N__5464\,
            in3 => \N__5518\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_188_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000001"
        )
    port map (
            in0 => \N__5404\,
            in1 => \N__5398\,
            in2 => \N__5461\,
            in3 => \N__6192\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8765\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9524\,
            in2 => \_gnd_net_\,
            in3 => \N__5473\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7842\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7137\,
            lcout => \U712_CHIP_RAM.N_306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIM32A1_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__7138\,
            in1 => \N__5428\,
            in2 => \_gnd_net_\,
            in3 => \N__6675\,
            lcout => \U712_CHIP_RAM.N_221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIRGPAB_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__7843\,
            in1 => \N__7139\,
            in2 => \N__6582\,
            in3 => \N__5410\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIND16J_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5397\,
            in2 => \N__5386\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5524\,
            in2 => \_gnd_net_\,
            in3 => \N__7140\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7051\,
            in1 => \N__7841\,
            in2 => \N__7897\,
            in3 => \N__6889\,
            lcout => \U712_CHIP_RAM.N_240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__7526\,
            in1 => \N__7050\,
            in2 => \N__6899\,
            in3 => \N__5991\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7845\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6129\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5541\,
            in1 => \N__5556\,
            in2 => \N__5578\,
            in3 => \N__5739\,
            lcout => \U712_CHIP_RAM.N_10\,
            ltout => \U712_CHIP_RAM.N_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_1_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7503\,
            in1 => \N__7028\,
            in2 => \N__5512\,
            in3 => \N__6621\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER16\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5509\,
            in3 => \N__7157\,
            lcout => \U712_CHIP_RAM.N_328\,
            ltout => \U712_CHIP_RAM.N_328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5497\,
            in2 => \N__5491\,
            in3 => \N__5487\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_251_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__7029\,
            in1 => \N__6092\,
            in2 => \N__5476\,
            in3 => \N__7883\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__6674\,
            in1 => \_gnd_net_\,
            in2 => \N__7162\,
            in3 => \N__7219\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_1_esr_RNO_0_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__7030\,
            in1 => \N__6091\,
            in2 => \N__5593\,
            in3 => \N__7884\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7049\,
            in2 => \_gnd_net_\,
            in3 => \N__5590\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \bfn_10_14_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7271\,
            in1 => \N__7516\,
            in2 => \_gnd_net_\,
            in3 => \N__5587\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__8779\,
            ce => \N__7183\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6893\,
            in2 => \_gnd_net_\,
            in3 => \N__5584\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7272\,
            in1 => \N__7959\,
            in2 => \_gnd_net_\,
            in3 => \N__5581\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__8779\,
            ce => \N__7183\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7266\,
            in1 => \N__5574\,
            in2 => \_gnd_net_\,
            in3 => \N__5560\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__8779\,
            ce => \N__7183\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7273\,
            in1 => \N__5557\,
            in2 => \_gnd_net_\,
            in3 => \N__5545\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__8779\,
            ce => \N__7183\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7267\,
            in1 => \N__5542\,
            in2 => \_gnd_net_\,
            in3 => \N__5530\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__8779\,
            ce => \N__7183\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__5740\,
            in1 => \N__7268\,
            in2 => \_gnd_net_\,
            in3 => \N__5527\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8779\,
            ce => \N__7183\,
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101011111"
        )
    port map (
            in0 => \N__8110\,
            in1 => \_gnd_net_\,
            in2 => \N__7849\,
            in3 => \N__8140\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8783\,
            ce => \N__6451\,
            sr => \N__9445\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5716\,
            in1 => \N__5695\,
            in2 => \_gnd_net_\,
            in3 => \N__8528\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8423\,
            in1 => \N__8548\,
            in2 => \N__5674\,
            in3 => \N__9151\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__8909\,
            in1 => \N__7600\,
            in2 => \N__8849\,
            in3 => \N__5665\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8754\,
            ce => \N__8664\,
            sr => \N__9486\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__8910\,
            in1 => \N__8840\,
            in2 => \N__7612\,
            in3 => \N__5830\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8754\,
            ce => \N__8664\,
            sr => \N__9486\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000111"
        )
    port map (
            in0 => \N__8523\,
            in1 => \N__9026\,
            in2 => \N__6245\,
            in3 => \N__6196\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA30_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5632\,
            in3 => \N__9526\,
            lcout => \U712_CHIP_RAM.un1_CMA30_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5629\,
            in1 => \N__5611\,
            in2 => \_gnd_net_\,
            in3 => \N__8526\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8527\,
            in1 => \N__8417\,
            in2 => \N__5833\,
            in3 => \N__9598\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5824\,
            in1 => \N__5803\,
            in2 => \_gnd_net_\,
            in3 => \N__8525\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5785\,
            in1 => \N__5767\,
            in2 => \_gnd_net_\,
            in3 => \N__8524\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_2_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__9020\,
            in1 => \N__8499\,
            in2 => \_gnd_net_\,
            in3 => \N__6185\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_2_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9021\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6186\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9MVM2_1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__7135\,
            in1 => \N__7535\,
            in2 => \N__6897\,
            in3 => \N__7441\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9MVM2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101010"
        )
    port map (
            in0 => \N__5752\,
            in1 => \N__7044\,
            in2 => \N__7161\,
            in3 => \N__6630\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110010"
        )
    port map (
            in0 => \N__7045\,
            in1 => \N__7978\,
            in2 => \N__5746\,
            in3 => \N__6880\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5743\,
            in3 => \N__5925\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8762\,
            ce => \N__6118\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110110"
        )
    port map (
            in0 => \N__7046\,
            in1 => \N__7979\,
            in2 => \N__6012\,
            in3 => \N__6879\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_66_0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__6881\,
            in1 => \N__5917\,
            in2 => \N__5929\,
            in3 => \N__5926\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8762\,
            ce => \N__6118\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111011101"
        )
    port map (
            in0 => \N__7043\,
            in1 => \N__7151\,
            in2 => \_gnd_net_\,
            in3 => \N__7534\,
            lcout => \U712_CHIP_RAM.N_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__7896\,
            in1 => \N__6992\,
            in2 => \N__5911\,
            in3 => \N__6093\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010110011111100"
        )
    port map (
            in0 => \N__6993\,
            in1 => \N__5856\,
            in2 => \N__5893\,
            in3 => \N__7549\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8766\,
            ce => 'H',
            sr => \N__9452\
        );

    \U712_CHIP_RAM.DMA_CYCLE_1_esr_RNO_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9523\,
            in2 => \_gnd_net_\,
            in3 => \N__5845\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_3_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7965\,
            in2 => \_gnd_net_\,
            in3 => \N__6844\,
            lcout => \U712_CHIP_RAM.N_305\,
            ltout => \U712_CHIP_RAM.N_305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6991\,
            in1 => \N__5989\,
            in2 => \N__5839\,
            in3 => \N__7527\,
            lcout => \U712_CHIP_RAM.N_254_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__7440\,
            in1 => \N__7001\,
            in2 => \_gnd_net_\,
            in3 => \N__6622\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__7002\,
            in1 => \N__7131\,
            in2 => \N__5836\,
            in3 => \N__7522\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__7007\,
            in1 => \N__6433\,
            in2 => \N__6133\,
            in3 => \N__6130\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8770\,
            ce => \N__6117\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7937\,
            in2 => \_gnd_net_\,
            in3 => \N__6828\,
            lcout => \U712_CHIP_RAM.N_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__7130\,
            in1 => \N__5990\,
            in2 => \_gnd_net_\,
            in3 => \N__7509\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__6097\,
            in1 => \N__7000\,
            in2 => \N__5938\,
            in3 => \N__7892\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__6030\,
            in1 => \N__7003\,
            in2 => \N__6073\,
            in3 => \N__6070\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8775\,
            ce => 'H',
            sr => \N__9446\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7156\,
            in2 => \_gnd_net_\,
            in3 => \N__6583\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOF0DC_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__7844\,
            in1 => \N__7858\,
            in2 => \N__6019\,
            in3 => \N__7220\,
            lcout => \U712_CHIP_RAM.N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7155\,
            in1 => \N__5979\,
            in2 => \_gnd_net_\,
            in3 => \N__7504\,
            lcout => \U712_CHIP_RAM.N_312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__6999\,
            in1 => \N__7505\,
            in2 => \N__6005\,
            in3 => \N__7063\,
            lcout => \U712_CHIP_RAM.N_260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7057\,
            in2 => \_gnd_net_\,
            in3 => \N__9521\,
            lcout => \U712_CYCLE_TERM.N_214_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000010"
        )
    port map (
            in0 => \N__7048\,
            in1 => \N__7958\,
            in2 => \N__6901\,
            in3 => \N__6442\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CRCSn_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6246\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8747\,
            ce => 'H',
            sr => \N__9495\
        );

    \U712_CHIP_RAM.WEn_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6211\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8747\,
            ce => 'H',
            sr => \N__9495\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__8430\,
            in1 => \N__6364\,
            in2 => \N__6349\,
            in3 => \N__6742\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8749\,
            ce => \N__8668\,
            sr => \N__9489\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__6741\,
            in1 => \N__6310\,
            in2 => \N__9337\,
            in3 => \N__8431\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8749\,
            ce => \N__8668\,
            sr => \N__9489\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__8911\,
            in1 => \N__8844\,
            in2 => \N__8932\,
            in3 => \N__6496\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8750\,
            ce => \N__8654\,
            sr => \N__9482\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__9033\,
            in1 => \N__6247\,
            in2 => \N__8572\,
            in3 => \N__6210\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8750\,
            ce => \N__8654\,
            sr => \N__9482\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__8912\,
            in1 => \N__9226\,
            in2 => \N__8850\,
            in3 => \N__6559\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8750\,
            ce => \N__8654\,
            sr => \N__9482\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6532\,
            in1 => \N__6517\,
            in2 => \_gnd_net_\,
            in3 => \N__8562\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8395\,
            in1 => \N__8564\,
            in2 => \N__6499\,
            in3 => \N__9187\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8394\,
            in2 => \_gnd_net_\,
            in3 => \N__8561\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__6490\,
            in1 => \N__8563\,
            in2 => \N__7561\,
            in3 => \N__8396\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000001010"
        )
    port map (
            in0 => \N__8889\,
            in1 => \N__8415\,
            in2 => \N__8570\,
            in3 => \N__8154\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111011"
        )
    port map (
            in0 => \N__8155\,
            in1 => \N__8554\,
            in2 => \N__8429\,
            in3 => \N__8890\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__6484\,
            in1 => \N__8416\,
            in2 => \N__8571\,
            in3 => \N__7567\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6478\,
            in2 => \N__6472\,
            in3 => \N__6469\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8753\,
            ce => \N__8671\,
            sr => \N__9467\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6691\,
            in1 => \N__6748\,
            in2 => \_gnd_net_\,
            in3 => \N__6754\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8753\,
            ce => \N__8671\,
            sr => \N__9467\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6775\,
            in1 => \N__8401\,
            in2 => \_gnd_net_\,
            in3 => \N__8188\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_316_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8888\,
            in2 => \N__6757\,
            in3 => \N__8565\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__6714\,
            in1 => \N__6731\,
            in2 => \N__8422\,
            in3 => \N__9114\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110110011"
        )
    port map (
            in0 => \N__8402\,
            in1 => \N__6732\,
            in2 => \N__6718\,
            in3 => \N__9115\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_1_esr_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7136\,
            in1 => \N__6685\,
            in2 => \_gnd_net_\,
            in3 => \N__7238\,
            lcout => \RAMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8759\,
            ce => \N__6640\,
            sr => \N__9450\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__7821\,
            in1 => \N__7133\,
            in2 => \N__7039\,
            in3 => \N__6626\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a3_2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6581\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8760\,
            ce => 'H',
            sr => \N__9448\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1_1_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__7822\,
            in1 => \N__6998\,
            in2 => \_gnd_net_\,
            in3 => \N__7536\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__8418\,
            in1 => \N__7420\,
            in2 => \N__7040\,
            in3 => \N__7429\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8760\,
            ce => 'H',
            sr => \N__9448\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7311\,
            in2 => \_gnd_net_\,
            in3 => \N__7419\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101110"
        )
    port map (
            in0 => \N__7312\,
            in1 => \N__7408\,
            in2 => \N__7381\,
            in3 => \N__7344\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8760\,
            ce => 'H',
            sr => \N__9448\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7303\,
            in1 => \N__7269\,
            in2 => \N__7239\,
            in3 => \N__7294\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8763\,
            ce => \N__7182\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7282\,
            in1 => \N__7270\,
            in2 => \N__7240\,
            in3 => \N__7195\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8763\,
            ce => \N__7182\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_2_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__7132\,
            in1 => \N__7980\,
            in2 => \_gnd_net_\,
            in3 => \N__6869\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__7823\,
            in1 => \N__8099\,
            in2 => \N__9049\,
            in3 => \N__8136\,
            lcout => \U712_CYCLE_TERM.N_214_i_0_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000000000"
        )
    port map (
            in0 => \N__6994\,
            in1 => \N__6845\,
            in2 => \N__7981\,
            in3 => \N__7885\,
            lcout => \U712_CHIP_RAM.N_243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7824\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7728\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7687\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__8919\,
            in1 => \N__8845\,
            in2 => \N__8242\,
            in3 => \N__7633\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8752\,
            ce => \N__8669\,
            sr => \N__9492\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8227\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9093\,
            ce => \N__9692\,
            sr => \N__9487\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7591\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9093\,
            ce => \N__9692\,
            sr => \N__9487\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7590\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__9588\,
            sr => \N__9476\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8182\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__9588\,
            sr => \N__9476\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8275\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9585\,
            sr => \N__9470\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8226\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9585\,
            sr => \N__9470\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8949\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9585\,
            sr => \N__9470\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8178\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9090\,
            ce => \N__9667\,
            sr => \N__9460\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011101100"
        )
    port map (
            in0 => \N__8062\,
            in1 => \N__8103\,
            in2 => \N__8035\,
            in3 => \N__8135\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8767\,
            ce => 'H',
            sr => \N__9453\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8030\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8064\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8771\,
            ce => 'H',
            sr => \N__9449\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9062\,
            in2 => \_gnd_net_\,
            in3 => \N__8082\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010001000100"
        )
    port map (
            in0 => \N__8029\,
            in1 => \N__9048\,
            in2 => \N__8143\,
            in3 => \N__8134\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8771\,
            ce => 'H',
            sr => \N__9449\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8083\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8771\,
            ce => 'H',
            sr => \N__9449\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110110000"
        )
    port map (
            in0 => \N__8063\,
            in1 => \N__8031\,
            in2 => \N__7998\,
            in3 => \N__9063\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8771\,
            ce => 'H',
            sr => \N__9449\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9064\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8776\,
            ce => 'H',
            sr => \N__9447\
        );

    \U712_CHIP_RAM.RASn_LC_14_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9034\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8748\,
            ce => 'H',
            sr => \N__9502\
        );

    \U712_CHIP_RAM.CASn_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8569\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8751\,
            ce => 'H',
            sr => \N__9501\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8956\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9094\,
            ce => \N__9691\,
            sr => \N__9497\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__8920\,
            in1 => \N__9217\,
            in2 => \N__8851\,
            in3 => \N__8281\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8758\,
            ce => \N__8670\,
            sr => \N__9493\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8608\,
            in1 => \N__8590\,
            in2 => \_gnd_net_\,
            in3 => \N__8552\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8553\,
            in1 => \N__8421\,
            in2 => \N__8284\,
            in3 => \N__9322\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8268\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9091\,
            ce => \N__9678\,
            sr => \N__9477\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9175\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9091\,
            ce => \N__9678\,
            sr => \N__9477\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9139\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__9578\,
            sr => \N__9471\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_8_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__9525\,
            in1 => \N__9277\,
            in2 => \_gnd_net_\,
            in3 => \N__9313\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_ctle_8_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__9522\,
            in1 => \N__9276\,
            in2 => \_gnd_net_\,
            in3 => \N__9100\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9211\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9096\,
            ce => \N__9694\,
            sr => \N__9500\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9631\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9095\,
            ce => \N__9693\,
            sr => \N__9498\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9204\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__9587\,
            sr => \N__9494\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_8_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9174\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_8C_net\,
            ce => \N__9586\,
            sr => \N__9488\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9138\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9092\,
            ce => \N__9668\,
            sr => \N__9478\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9630\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__9589\,
            sr => \N__9499\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 17 2025 18:30:33

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__12064\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK40_PLL_iso_i\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \N_929_i\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \LATCH_CLK_0_i\ : std_logic;
signal \C3_c\ : std_logic;
signal \INVU712_REG_SM.C3_SYNC_0C_net\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_390_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_346\ : std_logic;
signal \U712_CHIP_RAM.N_319\ : std_logic;
signal \U712_CHIP_RAM.N_229_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_345_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_\ : std_logic;
signal \LATCH_RAM\ : std_logic;
signal \U712_CHIP_RAM.N_379\ : std_logic;
signal \U712_CHIP_RAM.N_316_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0\ : std_logic;
signal \U712_CHIP_RAM.DBENn_8_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_316\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \LATCH_REG\ : std_logic;
signal \INVU712_REG_SM.C1_SYNC_1C_net\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_1\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \ASn_c\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.CYCLE_RUNZ0\ : std_logic;
signal \INVU712_REG_SM.C3_SYNC_1C_net\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \INVU712_REG_SM.C1_SYNC_0C_net\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_360\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.N_239_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto7_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_0_0_1_cascade_\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.N_323_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_367_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.N_374_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_418\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_418_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_0_a2_1_a2_0\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_229\ : std_logic;
signal \U712_CHIP_RAM.N_389_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_276\ : std_logic;
signal \U712_CHIP_RAM.N_389\ : std_logic;
signal \U712_CHIP_RAM.N_300\ : std_logic;
signal \U712_REG_SM.N_277_cascade_\ : std_logic;
signal \U712_REG_SM.N_236\ : std_logic;
signal \U712_REG_SM.N_277\ : std_logic;
signal \U712_REG_SM.N_236_cascade_\ : std_logic;
signal \U712_REG_SM.DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_437_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.N_244\ : std_logic;
signal \U712_REG_SM.N_244_cascade_\ : std_logic;
signal \U712_REG_SM.N_434\ : std_logic;
signal \N_275\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_9_4_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.N_57_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_436\ : std_logic;
signal \U712_CHIP_RAM.N_436_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_83\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_58\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_378\ : std_logic;
signal \U712_CHIP_RAM.N_367\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_237_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_3\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_5\ : std_logic;
signal \INVU712_REG_SM.STATE_COUNTER_5C_net\ : std_logic;
signal \U712_REG_SM.N_339\ : std_logic;
signal \U712_REG_SM.LDSn_7_iv_i_0\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \U712_REG_SM.UDSn_7_iv_i_0\ : std_logic;
signal \U712_REG_SM.N_337\ : std_logic;
signal \U712_REG_SM.N_169\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \REG_CPU_CYCLE\ : std_logic;
signal \U712_REG_SM.un15_0_i_0_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_7\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_255\ : std_logic;
signal \INVU712_REG_SM.LDSnC_net\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_6\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_274\ : std_logic;
signal \REG_WRITE_CYCLE\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERc_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_4\ : std_logic;
signal \U712_REG_SM.LATCH_REG_0_sqmuxa\ : std_logic;
signal \U712_REG_SM.REG_CPU_CYCLE_e_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_0_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_239\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_3\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_5_0_i_i_a2_0_a3_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_374\ : std_logic;
signal \WRITE_CYCLE\ : std_logic;
signal \U712_CHIP_RAM.N_130_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_60_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_57\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDs_0_6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \CLK40_PLL_g\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_r_sx_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_281\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_283\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_0\ : std_logic;
signal \U712_CHIP_RAM.N_130\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_292_cascade_\ : std_logic;
signal \N_207_i\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \N_205_i\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_248\ : std_logic;
signal \U712_CHIP_RAM.N_278\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_0_0_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_0_0_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_228\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_0_2\ : std_logic;
signal \U712_CHIP_RAM.N_50_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_50\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_263\ : std_logic;
signal \U712_CHIP_RAM.N_280_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDsr_0_3\ : std_logic;
signal \CLK40_PLL\ : std_logic;
signal \U712_CHIP_RAM.N_311\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDs_1_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDs_0_6\ : std_logic;
signal \U712_CHIP_RAM.N_377\ : std_logic;
signal \U712_CHIP_RAM.N_50_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.N_252_i_0_0_cascade_\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \CPU_TACK\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.un3_DMA_CYCLE_START\ : std_logic;
signal \U712_CYCLE_TERM.N_252_i_0_en\ : std_logic;
signal \U712_CYCLE_TERM.N_252_i_0_en_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_257\ : std_logic;
signal \U712_BYTE_ENABLE.N_258\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_BYTE_ENABLE.N_259\ : std_logic;
signal \N_222_i\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_11\ : std_logic;
signal \DMA_CYCLE\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_0Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_0Z0Z_0_cascade_\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \N_203_i\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_260\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \N_260_i\ : std_logic;
signal \N_259_i\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \N_257_i\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \N_258_i\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \RASn_c\ : std_logic;
signal \CASn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CPU_CYCLE\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \REG_CYCLE\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL\,
            REFERENCECLK => \N__4119\,
            RESETB => \N__6747\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12064\,
            DIN => \N__12063\,
            DOUT => \N__12062\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12064\,
            PADOUT => \N__12063\,
            PADIN => \N__12062\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8403\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12055\,
            DIN => \N__12054\,
            DOUT => \N__12053\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12055\,
            PADOUT => \N__12054\,
            PADIN => \N__12053\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12046\,
            DIN => \N__12045\,
            DOUT => \N__12044\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12046\,
            PADOUT => \N__12045\,
            PADIN => \N__12044\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9516\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12037\,
            DIN => \N__12036\,
            DOUT => \N__12035\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12037\,
            PADOUT => \N__12036\,
            PADIN => \N__12035\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4998\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12028\,
            DIN => \N__12027\,
            DOUT => \N__12026\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12028\,
            PADOUT => \N__12027\,
            PADIN => \N__12026\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12019\,
            DIN => \N__12018\,
            DOUT => \N__12017\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12019\,
            PADOUT => \N__12018\,
            PADIN => \N__12017\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12010\,
            DIN => \N__12009\,
            DOUT => \N__12008\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12010\,
            PADOUT => \N__12009\,
            PADIN => \N__12008\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12001\,
            DIN => \N__12000\,
            DOUT => \N__11999\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12001\,
            PADOUT => \N__12000\,
            PADIN => \N__11999\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11992\,
            DIN => \N__11991\,
            DOUT => \N__11990\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11992\,
            PADOUT => \N__11991\,
            PADIN => \N__11990\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11983\,
            DIN => \N__11982\,
            DOUT => \N__11981\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11983\,
            PADOUT => \N__11982\,
            PADIN => \N__11981\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11974\,
            DIN => \N__11973\,
            DOUT => \N__11972\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11974\,
            PADOUT => \N__11973\,
            PADIN => \N__11972\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8613\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11965\,
            DIN => \N__11964\,
            DOUT => \N__11963\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11965\,
            PADOUT => \N__11964\,
            PADIN => \N__11963\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8850\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11956\,
            DIN => \N__11955\,
            DOUT => \N__11954\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11956\,
            PADOUT => \N__11955\,
            PADIN => \N__11954\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11947\,
            DIN => \N__11946\,
            DOUT => \N__11945\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11947\,
            PADOUT => \N__11946\,
            PADIN => \N__11945\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11938\,
            DIN => \N__11937\,
            DOUT => \N__11936\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11938\,
            PADOUT => \N__11937\,
            PADIN => \N__11936\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11929\,
            DIN => \N__11928\,
            DOUT => \N__11927\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11929\,
            PADOUT => \N__11928\,
            PADIN => \N__11927\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4569\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11920\,
            DIN => \N__11919\,
            DOUT => \N__11918\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11920\,
            PADOUT => \N__11919\,
            PADIN => \N__11918\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11911\,
            DIN => \N__11910\,
            DOUT => \N__11909\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11911\,
            PADOUT => \N__11910\,
            PADIN => \N__11909\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11902\,
            DIN => \N__11901\,
            DOUT => \N__11900\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11902\,
            PADOUT => \N__11901\,
            PADIN => \N__11900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8724\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11893\,
            DIN => \N__11892\,
            DOUT => \N__11891\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11893\,
            PADOUT => \N__11892\,
            PADIN => \N__11891\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11884\,
            DIN => \N__11883\,
            DOUT => \N__11882\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11884\,
            PADOUT => \N__11883\,
            PADIN => \N__11882\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9543\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11875\,
            DIN => \N__11874\,
            DOUT => \N__11873\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11875\,
            PADOUT => \N__11874\,
            PADIN => \N__11873\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11866\,
            DIN => \N__11865\,
            DOUT => \N__11864\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11866\,
            PADOUT => \N__11865\,
            PADIN => \N__11864\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9894\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11857\,
            DIN => \N__11856\,
            DOUT => \N__11855\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11857\,
            PADOUT => \N__11856\,
            PADIN => \N__11855\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11848\,
            DIN => \N__11847\,
            DOUT => \N__11846\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11848\,
            PADOUT => \N__11847\,
            PADIN => \N__11846\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11839\,
            DIN => \N__11838\,
            DOUT => \N__11837\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11839\,
            PADOUT => \N__11838\,
            PADIN => \N__11837\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11830\,
            DIN => \N__11829\,
            DOUT => \N__11828\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11830\,
            PADOUT => \N__11829\,
            PADIN => \N__11828\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11821\,
            DIN => \N__11820\,
            DOUT => \N__11819\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11821\,
            PADOUT => \N__11820\,
            PADIN => \N__11819\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11812\,
            DIN => \N__11811\,
            DOUT => \N__11810\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11812\,
            PADOUT => \N__11811\,
            PADIN => \N__11810\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4994\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11803\,
            DIN => \N__11802\,
            DOUT => \N__11801\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11803\,
            PADOUT => \N__11802\,
            PADIN => \N__11801\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11794\,
            DIN => \N__11793\,
            DOUT => \N__11792\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11794\,
            PADOUT => \N__11793\,
            PADIN => \N__11792\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11785\,
            DIN => \N__11784\,
            DOUT => \N__11783\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11785\,
            PADOUT => \N__11784\,
            PADIN => \N__11783\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11776\,
            DIN => \N__11775\,
            DOUT => \N__11774\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11776\,
            PADOUT => \N__11775\,
            PADIN => \N__11774\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11767\,
            DIN => \N__11766\,
            DOUT => \N__11765\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11767\,
            PADOUT => \N__11766\,
            PADIN => \N__11765\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11758\,
            DIN => \N__11757\,
            DOUT => \N__11756\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11758\,
            PADOUT => \N__11757\,
            PADIN => \N__11756\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9528\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11749\,
            DIN => \N__11748\,
            DOUT => \N__11747\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11749\,
            PADOUT => \N__11748\,
            PADIN => \N__11747\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4710\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11740\,
            DIN => \N__11739\,
            DOUT => \N__11738\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11740\,
            PADOUT => \N__11739\,
            PADIN => \N__11738\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11731\,
            DIN => \N__11730\,
            DOUT => \N__11729\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11731\,
            PADOUT => \N__11730\,
            PADIN => \N__11729\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4491\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11722\,
            DIN => \N__11721\,
            DOUT => \N__11720\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11722\,
            PADOUT => \N__11721\,
            PADIN => \N__11720\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7857\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11713\,
            DIN => \N__11712\,
            DOUT => \N__11711\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11713\,
            PADOUT => \N__11712\,
            PADIN => \N__11711\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11704\,
            DIN => \N__11703\,
            DOUT => \N__11702\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11704\,
            PADOUT => \N__11703\,
            PADIN => \N__11702\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11695\,
            DIN => \N__11694\,
            DOUT => \N__11693\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11695\,
            PADOUT => \N__11694\,
            PADIN => \N__11693\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11686\,
            DIN => \N__11685\,
            DOUT => \N__11684\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11686\,
            PADOUT => \N__11685\,
            PADIN => \N__11684\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11677\,
            DIN => \N__11676\,
            DOUT => \N__11675\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11677\,
            PADOUT => \N__11676\,
            PADIN => \N__11675\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9144\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11668\,
            DIN => \N__11667\,
            DOUT => \N__11666\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11668\,
            PADOUT => \N__11667\,
            PADIN => \N__11666\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11659\,
            DIN => \N__11658\,
            DOUT => \N__11657\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11659\,
            PADOUT => \N__11658\,
            PADIN => \N__11657\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4228\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11650\,
            DIN => \N__11649\,
            DOUT => \N__11648\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11650\,
            PADOUT => \N__11649\,
            PADIN => \N__11648\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8649\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11641\,
            DIN => \N__11640\,
            DOUT => \N__11639\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11641\,
            PADOUT => \N__11640\,
            PADIN => \N__11639\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10971\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11632\,
            DIN => \N__11631\,
            DOUT => \N__11630\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11632\,
            PADOUT => \N__11631\,
            PADIN => \N__11630\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6693\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11623\,
            DIN => \N__11622\,
            DOUT => \N__11621\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11623\,
            PADOUT => \N__11622\,
            PADIN => \N__11621\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10704\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11614\,
            DIN => \N__11613\,
            DOUT => \N__11612\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11614\,
            PADOUT => \N__11613\,
            PADIN => \N__11612\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4518\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11605\,
            DIN => \N__11604\,
            DOUT => \N__11603\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11605\,
            PADOUT => \N__11604\,
            PADIN => \N__11603\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11596\,
            DIN => \N__11595\,
            DOUT => \N__11594\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11596\,
            PADOUT => \N__11595\,
            PADIN => \N__11594\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11587\,
            DIN => \N__11586\,
            DOUT => \N__11585\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11587\,
            PADOUT => \N__11586\,
            PADIN => \N__11585\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8079\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11578\,
            DIN => \N__11577\,
            DOUT => \N__11576\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11578\,
            PADOUT => \N__11577\,
            PADIN => \N__11576\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9495\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11569\,
            DIN => \N__11568\,
            DOUT => \N__11567\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11569\,
            PADOUT => \N__11568\,
            PADIN => \N__11567\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4425\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11560\,
            DIN => \N__11559\,
            DOUT => \N__11558\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11560\,
            PADOUT => \N__11559\,
            PADIN => \N__11558\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7497\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11551\,
            DIN => \N__11550\,
            DOUT => \N__11549\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11551\,
            PADOUT => \N__11550\,
            PADIN => \N__11549\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11542\,
            DIN => \N__11541\,
            DOUT => \N__11540\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11542\,
            PADOUT => \N__11541\,
            PADIN => \N__11540\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11533\,
            DIN => \N__11532\,
            DOUT => \N__11531\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11533\,
            PADOUT => \N__11532\,
            PADIN => \N__11531\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11524\,
            DIN => \N__11523\,
            DOUT => \N__11522\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11524\,
            PADOUT => \N__11523\,
            PADIN => \N__11522\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11515\,
            DIN => \N__11514\,
            DOUT => \N__11513\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11515\,
            PADOUT => \N__11514\,
            PADIN => \N__11513\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7869\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11506\,
            DIN => \N__11505\,
            DOUT => \N__11504\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11506\,
            PADOUT => \N__11505\,
            PADIN => \N__11504\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8835\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11497\,
            DIN => \N__11496\,
            DOUT => \N__11495\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11497\,
            PADOUT => \N__11496\,
            PADIN => \N__11495\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11488\,
            DIN => \N__11487\,
            DOUT => \N__11486\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11488\,
            PADOUT => \N__11487\,
            PADIN => \N__11486\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8337\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11479\,
            DIN => \N__11478\,
            DOUT => \N__11477\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11479\,
            PADOUT => \N__11478\,
            PADIN => \N__11477\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4170\,
            DIN0 => OPEN,
            DOUT0 => \N__4953\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11470\,
            DIN => \N__11469\,
            DOUT => \N__11468\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11470\,
            PADOUT => \N__11469\,
            PADIN => \N__11468\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8685\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11461\,
            DIN => \N__11460\,
            DOUT => \N__11459\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11461\,
            PADOUT => \N__11460\,
            PADIN => \N__11459\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11452\,
            DIN => \N__11451\,
            DOUT => \N__11450\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11452\,
            PADOUT => \N__11451\,
            PADIN => \N__11450\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11443\,
            DIN => \N__11442\,
            DOUT => \N__11441\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11443\,
            PADOUT => \N__11442\,
            PADIN => \N__11441\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10938\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11434\,
            DIN => \N__11433\,
            DOUT => \N__11432\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11434\,
            PADOUT => \N__11433\,
            PADIN => \N__11432\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11425\,
            DIN => \N__11424\,
            DOUT => \N__11423\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11425\,
            PADOUT => \N__11424\,
            PADIN => \N__11423\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11416\,
            DIN => \N__11415\,
            DOUT => \N__11414\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11416\,
            PADOUT => \N__11415\,
            PADIN => \N__11414\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11407\,
            DIN => \N__11406\,
            DOUT => \N__11405\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11407\,
            PADOUT => \N__11406\,
            PADIN => \N__11405\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11398\,
            DIN => \N__11397\,
            DOUT => \N__11396\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11398\,
            PADOUT => \N__11397\,
            PADIN => \N__11396\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8118\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11389\,
            DIN => \N__11388\,
            DOUT => \N__11387\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11389\,
            PADOUT => \N__11388\,
            PADIN => \N__11387\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5727\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11380\,
            DIN => \N__11379\,
            DOUT => \N__11378\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11380\,
            PADOUT => \N__11379\,
            PADIN => \N__11378\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9561\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11371\,
            DIN => \N__11370\,
            DOUT => \N__11369\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11371\,
            PADOUT => \N__11370\,
            PADIN => \N__11369\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6795\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11362\,
            DIN => \N__11361\,
            DOUT => \N__11360\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11362\,
            PADOUT => \N__11361\,
            PADIN => \N__11360\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11353\,
            DIN => \N__11352\,
            DOUT => \N__11351\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11353\,
            PADOUT => \N__11352\,
            PADIN => \N__11351\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11344\,
            DIN => \N__11343\,
            DOUT => \N__11342\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11344\,
            PADOUT => \N__11343\,
            PADIN => \N__11342\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8592\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11335\,
            DIN => \N__11334\,
            DOUT => \N__11333\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11335\,
            PADOUT => \N__11334\,
            PADIN => \N__11333\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11326\,
            DIN => \N__11325\,
            DOUT => \N__11324\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11326\,
            PADOUT => \N__11325\,
            PADIN => \N__11324\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11317\,
            DIN => \N__11316\,
            DOUT => \N__11315\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11317\,
            PADOUT => \N__11316\,
            PADIN => \N__11315\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4137\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11308\,
            DIN => \N__11307\,
            DOUT => \N__11306\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11308\,
            PADOUT => \N__11307\,
            PADIN => \N__11306\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5793\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11299\,
            DIN => \N__11298\,
            DOUT => \N__11297\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11299\,
            PADOUT => \N__11298\,
            PADIN => \N__11297\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4239\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11290\,
            DIN => \N__11289\,
            DOUT => \N__11288\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11290\,
            PADOUT => \N__11289\,
            PADIN => \N__11288\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11281\,
            DIN => \N__11280\,
            DOUT => \N__11279\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11281\,
            PADOUT => \N__11280\,
            PADIN => \N__11279\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4235\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11272\,
            DIN => \N__11271\,
            DOUT => \N__11270\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11272\,
            PADOUT => \N__11271\,
            PADIN => \N__11270\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4155\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2743\ : InMux
    port map (
            O => \N__11253\,
            I => \N__11246\
        );

    \I__2742\ : InMux
    port map (
            O => \N__11252\,
            I => \N__11243\
        );

    \I__2741\ : InMux
    port map (
            O => \N__11251\,
            I => \N__11240\
        );

    \I__2740\ : InMux
    port map (
            O => \N__11250\,
            I => \N__11237\
        );

    \I__2739\ : InMux
    port map (
            O => \N__11249\,
            I => \N__11234\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__11246\,
            I => \N__11229\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__11243\,
            I => \N__11226\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__11240\,
            I => \N__11219\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__11237\,
            I => \N__11189\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__11234\,
            I => \N__11182\
        );

    \I__2733\ : SRMux
    port map (
            O => \N__11233\,
            I => \N__11085\
        );

    \I__2732\ : SRMux
    port map (
            O => \N__11232\,
            I => \N__11085\
        );

    \I__2731\ : Glb2LocalMux
    port map (
            O => \N__11229\,
            I => \N__11085\
        );

    \I__2730\ : Glb2LocalMux
    port map (
            O => \N__11226\,
            I => \N__11085\
        );

    \I__2729\ : SRMux
    port map (
            O => \N__11225\,
            I => \N__11085\
        );

    \I__2728\ : SRMux
    port map (
            O => \N__11224\,
            I => \N__11085\
        );

    \I__2727\ : SRMux
    port map (
            O => \N__11223\,
            I => \N__11085\
        );

    \I__2726\ : SRMux
    port map (
            O => \N__11222\,
            I => \N__11085\
        );

    \I__2725\ : Glb2LocalMux
    port map (
            O => \N__11219\,
            I => \N__11085\
        );

    \I__2724\ : SRMux
    port map (
            O => \N__11218\,
            I => \N__11085\
        );

    \I__2723\ : SRMux
    port map (
            O => \N__11217\,
            I => \N__11085\
        );

    \I__2722\ : SRMux
    port map (
            O => \N__11216\,
            I => \N__11085\
        );

    \I__2721\ : SRMux
    port map (
            O => \N__11215\,
            I => \N__11085\
        );

    \I__2720\ : SRMux
    port map (
            O => \N__11214\,
            I => \N__11085\
        );

    \I__2719\ : SRMux
    port map (
            O => \N__11213\,
            I => \N__11085\
        );

    \I__2718\ : SRMux
    port map (
            O => \N__11212\,
            I => \N__11085\
        );

    \I__2717\ : SRMux
    port map (
            O => \N__11211\,
            I => \N__11085\
        );

    \I__2716\ : SRMux
    port map (
            O => \N__11210\,
            I => \N__11085\
        );

    \I__2715\ : SRMux
    port map (
            O => \N__11209\,
            I => \N__11085\
        );

    \I__2714\ : SRMux
    port map (
            O => \N__11208\,
            I => \N__11085\
        );

    \I__2713\ : SRMux
    port map (
            O => \N__11207\,
            I => \N__11085\
        );

    \I__2712\ : SRMux
    port map (
            O => \N__11206\,
            I => \N__11085\
        );

    \I__2711\ : SRMux
    port map (
            O => \N__11205\,
            I => \N__11085\
        );

    \I__2710\ : SRMux
    port map (
            O => \N__11204\,
            I => \N__11085\
        );

    \I__2709\ : SRMux
    port map (
            O => \N__11203\,
            I => \N__11085\
        );

    \I__2708\ : SRMux
    port map (
            O => \N__11202\,
            I => \N__11085\
        );

    \I__2707\ : SRMux
    port map (
            O => \N__11201\,
            I => \N__11085\
        );

    \I__2706\ : SRMux
    port map (
            O => \N__11200\,
            I => \N__11085\
        );

    \I__2705\ : SRMux
    port map (
            O => \N__11199\,
            I => \N__11085\
        );

    \I__2704\ : SRMux
    port map (
            O => \N__11198\,
            I => \N__11085\
        );

    \I__2703\ : SRMux
    port map (
            O => \N__11197\,
            I => \N__11085\
        );

    \I__2702\ : SRMux
    port map (
            O => \N__11196\,
            I => \N__11085\
        );

    \I__2701\ : SRMux
    port map (
            O => \N__11195\,
            I => \N__11085\
        );

    \I__2700\ : SRMux
    port map (
            O => \N__11194\,
            I => \N__11085\
        );

    \I__2699\ : SRMux
    port map (
            O => \N__11193\,
            I => \N__11085\
        );

    \I__2698\ : SRMux
    port map (
            O => \N__11192\,
            I => \N__11085\
        );

    \I__2697\ : Glb2LocalMux
    port map (
            O => \N__11189\,
            I => \N__11085\
        );

    \I__2696\ : SRMux
    port map (
            O => \N__11188\,
            I => \N__11085\
        );

    \I__2695\ : SRMux
    port map (
            O => \N__11187\,
            I => \N__11085\
        );

    \I__2694\ : SRMux
    port map (
            O => \N__11186\,
            I => \N__11085\
        );

    \I__2693\ : SRMux
    port map (
            O => \N__11185\,
            I => \N__11085\
        );

    \I__2692\ : Glb2LocalMux
    port map (
            O => \N__11182\,
            I => \N__11085\
        );

    \I__2691\ : SRMux
    port map (
            O => \N__11181\,
            I => \N__11085\
        );

    \I__2690\ : SRMux
    port map (
            O => \N__11180\,
            I => \N__11085\
        );

    \I__2689\ : SRMux
    port map (
            O => \N__11179\,
            I => \N__11085\
        );

    \I__2688\ : SRMux
    port map (
            O => \N__11178\,
            I => \N__11085\
        );

    \I__2687\ : GlobalMux
    port map (
            O => \N__11085\,
            I => \N__11082\
        );

    \I__2686\ : gio2CtrlBuf
    port map (
            O => \N__11082\,
            I => \RESETn_c_i_g\
        );

    \I__2685\ : InMux
    port map (
            O => \N__11079\,
            I => \N__11076\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__11076\,
            I => \N__11072\
        );

    \I__2683\ : InMux
    port map (
            O => \N__11075\,
            I => \N__11069\
        );

    \I__2682\ : Span4Mux_v
    port map (
            O => \N__11072\,
            I => \N__11064\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__11069\,
            I => \N__11064\
        );

    \I__2680\ : Span4Mux_v
    port map (
            O => \N__11064\,
            I => \N__11061\
        );

    \I__2679\ : Sp12to4
    port map (
            O => \N__11061\,
            I => \N__11057\
        );

    \I__2678\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11054\
        );

    \I__2677\ : Span12Mux_h
    port map (
            O => \N__11057\,
            I => \N__11049\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__11054\,
            I => \N__11049\
        );

    \I__2675\ : Span12Mux_v
    port map (
            O => \N__11049\,
            I => \N__11046\
        );

    \I__2674\ : Odrv12
    port map (
            O => \N__11046\,
            I => \CASLn_c\
        );

    \I__2673\ : InMux
    port map (
            O => \N__11043\,
            I => \N__11039\
        );

    \I__2672\ : InMux
    port map (
            O => \N__11042\,
            I => \N__11036\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__11039\,
            I => \N__11031\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__11036\,
            I => \N__11031\
        );

    \I__2669\ : Span4Mux_v
    port map (
            O => \N__11031\,
            I => \N__11027\
        );

    \I__2668\ : InMux
    port map (
            O => \N__11030\,
            I => \N__11024\
        );

    \I__2667\ : Sp12to4
    port map (
            O => \N__11027\,
            I => \N__11021\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__11024\,
            I => \N__11018\
        );

    \I__2665\ : Span12Mux_h
    port map (
            O => \N__11021\,
            I => \N__11015\
        );

    \I__2664\ : Span4Mux_h
    port map (
            O => \N__11018\,
            I => \N__11012\
        );

    \I__2663\ : Span12Mux_v
    port map (
            O => \N__11015\,
            I => \N__11009\
        );

    \I__2662\ : Span4Mux_v
    port map (
            O => \N__11012\,
            I => \N__11006\
        );

    \I__2661\ : Odrv12
    port map (
            O => \N__11009\,
            I => \CASUn_c\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__11006\,
            I => \CASUn_c\
        );

    \I__2659\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10998\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__10998\,
            I => \N__10995\
        );

    \I__2657\ : Span12Mux_v
    port map (
            O => \N__10995\,
            I => \N__10991\
        );

    \I__2656\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10988\
        );

    \I__2655\ : Span12Mux_h
    port map (
            O => \N__10991\,
            I => \N__10984\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__10988\,
            I => \N__10981\
        );

    \I__2653\ : InMux
    port map (
            O => \N__10987\,
            I => \N__10978\
        );

    \I__2652\ : Odrv12
    port map (
            O => \N__10984\,
            I => \REG_CYCLE\
        );

    \I__2651\ : Odrv4
    port map (
            O => \N__10981\,
            I => \REG_CYCLE\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__10978\,
            I => \REG_CYCLE\
        );

    \I__2649\ : IoInMux
    port map (
            O => \N__10971\,
            I => \N__10968\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__10968\,
            I => \N__10965\
        );

    \I__2647\ : Span4Mux_s3_v
    port map (
            O => \N__10965\,
            I => \N__10962\
        );

    \I__2646\ : Span4Mux_v
    port map (
            O => \N__10962\,
            I => \N__10959\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__10959\,
            I => \DRDENn_c\
        );

    \I__2644\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10953\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__10953\,
            I => \N__10950\
        );

    \I__2642\ : Sp12to4
    port map (
            O => \N__10950\,
            I => \N__10947\
        );

    \I__2641\ : Span12Mux_v
    port map (
            O => \N__10947\,
            I => \N__10944\
        );

    \I__2640\ : Span12Mux_h
    port map (
            O => \N__10944\,
            I => \N__10941\
        );

    \I__2639\ : Odrv12
    port map (
            O => \N__10941\,
            I => \A_c_17\
        );

    \I__2638\ : IoInMux
    port map (
            O => \N__10938\,
            I => \N__10935\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__10935\,
            I => \N__10932\
        );

    \I__2636\ : IoSpan4Mux
    port map (
            O => \N__10932\,
            I => \N__10929\
        );

    \I__2635\ : Span4Mux_s0_h
    port map (
            O => \N__10929\,
            I => \N__10926\
        );

    \I__2634\ : Sp12to4
    port map (
            O => \N__10926\,
            I => \N__10923\
        );

    \I__2633\ : Span12Mux_h
    port map (
            O => \N__10923\,
            I => \N__10920\
        );

    \I__2632\ : Odrv12
    port map (
            O => \N__10920\,
            I => \CMA_c_8\
        );

    \I__2631\ : InMux
    port map (
            O => \N__10917\,
            I => \N__10913\
        );

    \I__2630\ : InMux
    port map (
            O => \N__10916\,
            I => \N__10910\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__10913\,
            I => \N__10903\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__10910\,
            I => \N__10903\
        );

    \I__2627\ : InMux
    port map (
            O => \N__10909\,
            I => \N__10898\
        );

    \I__2626\ : InMux
    port map (
            O => \N__10908\,
            I => \N__10898\
        );

    \I__2625\ : Odrv12
    port map (
            O => \N__10903\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__10898\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__2623\ : CascadeMux
    port map (
            O => \N__10893\,
            I => \N__10890\
        );

    \I__2622\ : InMux
    port map (
            O => \N__10890\,
            I => \N__10887\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__10887\,
            I => \N__10884\
        );

    \I__2620\ : Sp12to4
    port map (
            O => \N__10884\,
            I => \N__10881\
        );

    \I__2619\ : Span12Mux_v
    port map (
            O => \N__10881\,
            I => \N__10878\
        );

    \I__2618\ : Span12Mux_h
    port map (
            O => \N__10878\,
            I => \N__10875\
        );

    \I__2617\ : Odrv12
    port map (
            O => \N__10875\,
            I => \A_c_19\
        );

    \I__2616\ : CascadeMux
    port map (
            O => \N__10872\,
            I => \N__10868\
        );

    \I__2615\ : InMux
    port map (
            O => \N__10871\,
            I => \N__10859\
        );

    \I__2614\ : InMux
    port map (
            O => \N__10868\,
            I => \N__10856\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__10867\,
            I => \N__10850\
        );

    \I__2612\ : InMux
    port map (
            O => \N__10866\,
            I => \N__10845\
        );

    \I__2611\ : InMux
    port map (
            O => \N__10865\,
            I => \N__10839\
        );

    \I__2610\ : InMux
    port map (
            O => \N__10864\,
            I => \N__10834\
        );

    \I__2609\ : InMux
    port map (
            O => \N__10863\,
            I => \N__10834\
        );

    \I__2608\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10830\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__10859\,
            I => \N__10825\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__10856\,
            I => \N__10825\
        );

    \I__2605\ : InMux
    port map (
            O => \N__10855\,
            I => \N__10822\
        );

    \I__2604\ : InMux
    port map (
            O => \N__10854\,
            I => \N__10817\
        );

    \I__2603\ : InMux
    port map (
            O => \N__10853\,
            I => \N__10817\
        );

    \I__2602\ : InMux
    port map (
            O => \N__10850\,
            I => \N__10812\
        );

    \I__2601\ : InMux
    port map (
            O => \N__10849\,
            I => \N__10812\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__10848\,
            I => \N__10808\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__10845\,
            I => \N__10805\
        );

    \I__2598\ : InMux
    port map (
            O => \N__10844\,
            I => \N__10797\
        );

    \I__2597\ : InMux
    port map (
            O => \N__10843\,
            I => \N__10797\
        );

    \I__2596\ : InMux
    port map (
            O => \N__10842\,
            I => \N__10797\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__10839\,
            I => \N__10789\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__10834\,
            I => \N__10789\
        );

    \I__2593\ : InMux
    port map (
            O => \N__10833\,
            I => \N__10786\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__10830\,
            I => \N__10775\
        );

    \I__2591\ : Span4Mux_h
    port map (
            O => \N__10825\,
            I => \N__10775\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__10822\,
            I => \N__10775\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__10817\,
            I => \N__10775\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__10812\,
            I => \N__10775\
        );

    \I__2587\ : InMux
    port map (
            O => \N__10811\,
            I => \N__10772\
        );

    \I__2586\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10768\
        );

    \I__2585\ : Span4Mux_v
    port map (
            O => \N__10805\,
            I => \N__10764\
        );

    \I__2584\ : InMux
    port map (
            O => \N__10804\,
            I => \N__10761\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__10797\,
            I => \N__10758\
        );

    \I__2582\ : InMux
    port map (
            O => \N__10796\,
            I => \N__10751\
        );

    \I__2581\ : InMux
    port map (
            O => \N__10795\,
            I => \N__10751\
        );

    \I__2580\ : InMux
    port map (
            O => \N__10794\,
            I => \N__10751\
        );

    \I__2579\ : Span4Mux_h
    port map (
            O => \N__10789\,
            I => \N__10748\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__10786\,
            I => \N__10741\
        );

    \I__2577\ : Span4Mux_h
    port map (
            O => \N__10775\,
            I => \N__10741\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__10772\,
            I => \N__10741\
        );

    \I__2575\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10738\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__10768\,
            I => \N__10735\
        );

    \I__2573\ : InMux
    port map (
            O => \N__10767\,
            I => \N__10732\
        );

    \I__2572\ : Sp12to4
    port map (
            O => \N__10764\,
            I => \N__10723\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__10761\,
            I => \N__10723\
        );

    \I__2570\ : Sp12to4
    port map (
            O => \N__10758\,
            I => \N__10723\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__10751\,
            I => \N__10723\
        );

    \I__2568\ : Span4Mux_h
    port map (
            O => \N__10748\,
            I => \N__10720\
        );

    \I__2567\ : Span4Mux_h
    port map (
            O => \N__10741\,
            I => \N__10717\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__10738\,
            I => \CPU_CYCLE\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__10735\,
            I => \CPU_CYCLE\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__10732\,
            I => \CPU_CYCLE\
        );

    \I__2563\ : Odrv12
    port map (
            O => \N__10723\,
            I => \CPU_CYCLE\
        );

    \I__2562\ : Odrv4
    port map (
            O => \N__10720\,
            I => \CPU_CYCLE\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__10717\,
            I => \CPU_CYCLE\
        );

    \I__2560\ : IoInMux
    port map (
            O => \N__10704\,
            I => \N__10701\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__10701\,
            I => \N__10698\
        );

    \I__2558\ : Span4Mux_s2_h
    port map (
            O => \N__10698\,
            I => \N__10695\
        );

    \I__2557\ : Span4Mux_v
    port map (
            O => \N__10695\,
            I => \N__10692\
        );

    \I__2556\ : Sp12to4
    port map (
            O => \N__10692\,
            I => \N__10689\
        );

    \I__2555\ : Span12Mux_h
    port map (
            O => \N__10689\,
            I => \N__10686\
        );

    \I__2554\ : Odrv12
    port map (
            O => \N__10686\,
            I => \CMA_c_9\
        );

    \I__2553\ : InMux
    port map (
            O => \N__10683\,
            I => \N__10680\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10680\,
            I => \N__10653\
        );

    \I__2551\ : ClkMux
    port map (
            O => \N__10679\,
            I => \N__10575\
        );

    \I__2550\ : ClkMux
    port map (
            O => \N__10678\,
            I => \N__10575\
        );

    \I__2549\ : ClkMux
    port map (
            O => \N__10677\,
            I => \N__10575\
        );

    \I__2548\ : ClkMux
    port map (
            O => \N__10676\,
            I => \N__10575\
        );

    \I__2547\ : ClkMux
    port map (
            O => \N__10675\,
            I => \N__10575\
        );

    \I__2546\ : ClkMux
    port map (
            O => \N__10674\,
            I => \N__10575\
        );

    \I__2545\ : ClkMux
    port map (
            O => \N__10673\,
            I => \N__10575\
        );

    \I__2544\ : ClkMux
    port map (
            O => \N__10672\,
            I => \N__10575\
        );

    \I__2543\ : ClkMux
    port map (
            O => \N__10671\,
            I => \N__10575\
        );

    \I__2542\ : ClkMux
    port map (
            O => \N__10670\,
            I => \N__10575\
        );

    \I__2541\ : ClkMux
    port map (
            O => \N__10669\,
            I => \N__10575\
        );

    \I__2540\ : ClkMux
    port map (
            O => \N__10668\,
            I => \N__10575\
        );

    \I__2539\ : ClkMux
    port map (
            O => \N__10667\,
            I => \N__10575\
        );

    \I__2538\ : ClkMux
    port map (
            O => \N__10666\,
            I => \N__10575\
        );

    \I__2537\ : ClkMux
    port map (
            O => \N__10665\,
            I => \N__10575\
        );

    \I__2536\ : ClkMux
    port map (
            O => \N__10664\,
            I => \N__10575\
        );

    \I__2535\ : ClkMux
    port map (
            O => \N__10663\,
            I => \N__10575\
        );

    \I__2534\ : ClkMux
    port map (
            O => \N__10662\,
            I => \N__10575\
        );

    \I__2533\ : ClkMux
    port map (
            O => \N__10661\,
            I => \N__10575\
        );

    \I__2532\ : ClkMux
    port map (
            O => \N__10660\,
            I => \N__10575\
        );

    \I__2531\ : ClkMux
    port map (
            O => \N__10659\,
            I => \N__10575\
        );

    \I__2530\ : ClkMux
    port map (
            O => \N__10658\,
            I => \N__10575\
        );

    \I__2529\ : ClkMux
    port map (
            O => \N__10657\,
            I => \N__10575\
        );

    \I__2528\ : ClkMux
    port map (
            O => \N__10656\,
            I => \N__10575\
        );

    \I__2527\ : Glb2LocalMux
    port map (
            O => \N__10653\,
            I => \N__10575\
        );

    \I__2526\ : ClkMux
    port map (
            O => \N__10652\,
            I => \N__10575\
        );

    \I__2525\ : ClkMux
    port map (
            O => \N__10651\,
            I => \N__10575\
        );

    \I__2524\ : ClkMux
    port map (
            O => \N__10650\,
            I => \N__10575\
        );

    \I__2523\ : ClkMux
    port map (
            O => \N__10649\,
            I => \N__10575\
        );

    \I__2522\ : ClkMux
    port map (
            O => \N__10648\,
            I => \N__10575\
        );

    \I__2521\ : ClkMux
    port map (
            O => \N__10647\,
            I => \N__10575\
        );

    \I__2520\ : ClkMux
    port map (
            O => \N__10646\,
            I => \N__10575\
        );

    \I__2519\ : ClkMux
    port map (
            O => \N__10645\,
            I => \N__10575\
        );

    \I__2518\ : ClkMux
    port map (
            O => \N__10644\,
            I => \N__10575\
        );

    \I__2517\ : GlobalMux
    port map (
            O => \N__10575\,
            I => \CLK80_PLL\
        );

    \I__2516\ : CEMux
    port map (
            O => \N__10572\,
            I => \N__10567\
        );

    \I__2515\ : CEMux
    port map (
            O => \N__10571\,
            I => \N__10561\
        );

    \I__2514\ : CEMux
    port map (
            O => \N__10570\,
            I => \N__10558\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__10567\,
            I => \N__10554\
        );

    \I__2512\ : CEMux
    port map (
            O => \N__10566\,
            I => \N__10551\
        );

    \I__2511\ : CEMux
    port map (
            O => \N__10565\,
            I => \N__10548\
        );

    \I__2510\ : CEMux
    port map (
            O => \N__10564\,
            I => \N__10545\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__10561\,
            I => \N__10542\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10558\,
            I => \N__10539\
        );

    \I__2507\ : CEMux
    port map (
            O => \N__10557\,
            I => \N__10536\
        );

    \I__2506\ : Span4Mux_h
    port map (
            O => \N__10554\,
            I => \N__10533\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__10551\,
            I => \N__10528\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__10548\,
            I => \N__10528\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10545\,
            I => \N__10525\
        );

    \I__2502\ : Span4Mux_h
    port map (
            O => \N__10542\,
            I => \N__10522\
        );

    \I__2501\ : Span4Mux_v
    port map (
            O => \N__10539\,
            I => \N__10519\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__10536\,
            I => \N__10516\
        );

    \I__2499\ : Span4Mux_h
    port map (
            O => \N__10533\,
            I => \N__10511\
        );

    \I__2498\ : Span4Mux_v
    port map (
            O => \N__10528\,
            I => \N__10511\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__10525\,
            I => \N__10508\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__10522\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2495\ : Odrv4
    port map (
            O => \N__10519\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2494\ : Odrv12
    port map (
            O => \N__10516\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2493\ : Odrv4
    port map (
            O => \N__10511\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__10508\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2491\ : InMux
    port map (
            O => \N__10497\,
            I => \N__10494\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10494\,
            I => \N__10491\
        );

    \I__2489\ : Span4Mux_v
    port map (
            O => \N__10491\,
            I => \N__10488\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__10488\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2487\ : InMux
    port map (
            O => \N__10485\,
            I => \N__10479\
        );

    \I__2486\ : InMux
    port map (
            O => \N__10484\,
            I => \N__10476\
        );

    \I__2485\ : InMux
    port map (
            O => \N__10483\,
            I => \N__10473\
        );

    \I__2484\ : InMux
    port map (
            O => \N__10482\,
            I => \N__10470\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__10479\,
            I => \N__10467\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__10476\,
            I => \N__10460\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__10473\,
            I => \N__10460\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__10470\,
            I => \N__10460\
        );

    \I__2479\ : Sp12to4
    port map (
            O => \N__10467\,
            I => \N__10457\
        );

    \I__2478\ : Span4Mux_v
    port map (
            O => \N__10460\,
            I => \N__10454\
        );

    \I__2477\ : Span12Mux_v
    port map (
            O => \N__10457\,
            I => \N__10449\
        );

    \I__2476\ : Sp12to4
    port map (
            O => \N__10454\,
            I => \N__10449\
        );

    \I__2475\ : Span12Mux_h
    port map (
            O => \N__10449\,
            I => \N__10446\
        );

    \I__2474\ : Odrv12
    port map (
            O => \N__10446\,
            I => \DRA_c_8\
        );

    \I__2473\ : InMux
    port map (
            O => \N__10443\,
            I => \N__10440\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__10440\,
            I => \N__10437\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__10437\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2470\ : InMux
    port map (
            O => \N__10434\,
            I => \N__10430\
        );

    \I__2469\ : InMux
    port map (
            O => \N__10433\,
            I => \N__10426\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__10430\,
            I => \N__10423\
        );

    \I__2467\ : InMux
    port map (
            O => \N__10429\,
            I => \N__10420\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10426\,
            I => \N__10416\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__10423\,
            I => \N__10411\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__10420\,
            I => \N__10411\
        );

    \I__2463\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10408\
        );

    \I__2462\ : Span4Mux_v
    port map (
            O => \N__10416\,
            I => \N__10403\
        );

    \I__2461\ : Span4Mux_v
    port map (
            O => \N__10411\,
            I => \N__10403\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__10408\,
            I => \N__10398\
        );

    \I__2459\ : Sp12to4
    port map (
            O => \N__10403\,
            I => \N__10398\
        );

    \I__2458\ : Span12Mux_h
    port map (
            O => \N__10398\,
            I => \N__10395\
        );

    \I__2457\ : Span12Mux_v
    port map (
            O => \N__10395\,
            I => \N__10392\
        );

    \I__2456\ : Odrv12
    port map (
            O => \N__10392\,
            I => \DRA_c_1\
        );

    \I__2455\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10386\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__10386\,
            I => \N__10383\
        );

    \I__2453\ : Span4Mux_v
    port map (
            O => \N__10383\,
            I => \N__10379\
        );

    \I__2452\ : InMux
    port map (
            O => \N__10382\,
            I => \N__10376\
        );

    \I__2451\ : Sp12to4
    port map (
            O => \N__10379\,
            I => \N__10371\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10376\,
            I => \N__10371\
        );

    \I__2449\ : Span12Mux_h
    port map (
            O => \N__10371\,
            I => \N__10368\
        );

    \I__2448\ : Span12Mux_v
    port map (
            O => \N__10368\,
            I => \N__10365\
        );

    \I__2447\ : Odrv12
    port map (
            O => \N__10365\,
            I => \DRA_c_0\
        );

    \I__2446\ : InMux
    port map (
            O => \N__10362\,
            I => \N__10359\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__10359\,
            I => \N__10356\
        );

    \I__2444\ : Span4Mux_v
    port map (
            O => \N__10356\,
            I => \N__10353\
        );

    \I__2443\ : Odrv4
    port map (
            O => \N__10353\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10350\,
            I => \N__10347\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__10347\,
            I => \N__10342\
        );

    \I__2440\ : InMux
    port map (
            O => \N__10346\,
            I => \N__10339\
        );

    \I__2439\ : InMux
    port map (
            O => \N__10345\,
            I => \N__10335\
        );

    \I__2438\ : Span4Mux_h
    port map (
            O => \N__10342\,
            I => \N__10330\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__10339\,
            I => \N__10330\
        );

    \I__2436\ : InMux
    port map (
            O => \N__10338\,
            I => \N__10327\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__10335\,
            I => \N__10320\
        );

    \I__2434\ : Span4Mux_h
    port map (
            O => \N__10330\,
            I => \N__10320\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__10327\,
            I => \N__10320\
        );

    \I__2432\ : Span4Mux_v
    port map (
            O => \N__10320\,
            I => \N__10317\
        );

    \I__2431\ : Sp12to4
    port map (
            O => \N__10317\,
            I => \N__10314\
        );

    \I__2430\ : Span12Mux_h
    port map (
            O => \N__10314\,
            I => \N__10311\
        );

    \I__2429\ : Odrv12
    port map (
            O => \N__10311\,
            I => \DRA_c_7\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__10308\,
            I => \N__10305\
        );

    \I__2427\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10302\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__10302\,
            I => \N__10299\
        );

    \I__2425\ : Odrv4
    port map (
            O => \N__10299\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2424\ : InMux
    port map (
            O => \N__10296\,
            I => \N__10293\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__10293\,
            I => \N__10290\
        );

    \I__2422\ : Span12Mux_h
    port map (
            O => \N__10290\,
            I => \N__10287\
        );

    \I__2421\ : Odrv12
    port map (
            O => \N__10287\,
            I => \RAS0n_c\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__10284\,
            I => \N__10280\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10277\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10280\,
            I => \N__10274\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__10277\,
            I => \N__10269\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__10274\,
            I => \N__10266\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10273\,
            I => \N__10263\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10272\,
            I => \N__10260\
        );

    \I__2413\ : Span4Mux_h
    port map (
            O => \N__10269\,
            I => \N__10251\
        );

    \I__2412\ : Span4Mux_v
    port map (
            O => \N__10266\,
            I => \N__10251\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__10263\,
            I => \N__10251\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__10260\,
            I => \N__10251\
        );

    \I__2409\ : Span4Mux_h
    port map (
            O => \N__10251\,
            I => \N__10248\
        );

    \I__2408\ : Span4Mux_v
    port map (
            O => \N__10248\,
            I => \N__10245\
        );

    \I__2407\ : Sp12to4
    port map (
            O => \N__10245\,
            I => \N__10242\
        );

    \I__2406\ : Span12Mux_v
    port map (
            O => \N__10242\,
            I => \N__10239\
        );

    \I__2405\ : Odrv12
    port map (
            O => \N__10239\,
            I => \DRA_c_9\
        );

    \I__2404\ : InMux
    port map (
            O => \N__10236\,
            I => \N__10233\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__10233\,
            I => \N__10230\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__10230\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2401\ : InMux
    port map (
            O => \N__10227\,
            I => \N__10221\
        );

    \I__2400\ : InMux
    port map (
            O => \N__10226\,
            I => \N__10216\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10225\,
            I => \N__10216\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10224\,
            I => \N__10213\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__10221\,
            I => \N__10208\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__10216\,
            I => \N__10208\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__10213\,
            I => \N__10205\
        );

    \I__2394\ : Span12Mux_v
    port map (
            O => \N__10208\,
            I => \N__10202\
        );

    \I__2393\ : Sp12to4
    port map (
            O => \N__10205\,
            I => \N__10199\
        );

    \I__2392\ : Span12Mux_h
    port map (
            O => \N__10202\,
            I => \N__10196\
        );

    \I__2391\ : Span12Mux_v
    port map (
            O => \N__10199\,
            I => \N__10193\
        );

    \I__2390\ : Odrv12
    port map (
            O => \N__10196\,
            I => \DRA_c_5\
        );

    \I__2389\ : Odrv12
    port map (
            O => \N__10193\,
            I => \DRA_c_5\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10188\,
            I => \N__10183\
        );

    \I__2387\ : InMux
    port map (
            O => \N__10187\,
            I => \N__10180\
        );

    \I__2386\ : InMux
    port map (
            O => \N__10186\,
            I => \N__10177\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__10183\,
            I => \N__10173\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10180\,
            I => \N__10168\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__10177\,
            I => \N__10168\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10176\,
            I => \N__10165\
        );

    \I__2381\ : Span4Mux_v
    port map (
            O => \N__10173\,
            I => \N__10162\
        );

    \I__2380\ : Span4Mux_h
    port map (
            O => \N__10168\,
            I => \N__10159\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__10165\,
            I => \N__10156\
        );

    \I__2378\ : Span4Mux_v
    port map (
            O => \N__10162\,
            I => \N__10153\
        );

    \I__2377\ : Sp12to4
    port map (
            O => \N__10159\,
            I => \N__10148\
        );

    \I__2376\ : Sp12to4
    port map (
            O => \N__10156\,
            I => \N__10148\
        );

    \I__2375\ : Sp12to4
    port map (
            O => \N__10153\,
            I => \N__10143\
        );

    \I__2374\ : Span12Mux_v
    port map (
            O => \N__10148\,
            I => \N__10143\
        );

    \I__2373\ : Odrv12
    port map (
            O => \N__10143\,
            I => \DRA_c_6\
        );

    \I__2372\ : InMux
    port map (
            O => \N__10140\,
            I => \N__10137\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10137\,
            I => \N__10134\
        );

    \I__2370\ : Span4Mux_v
    port map (
            O => \N__10134\,
            I => \N__10126\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10123\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10132\,
            I => \N__10120\
        );

    \I__2367\ : InMux
    port map (
            O => \N__10131\,
            I => \N__10117\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10114\
        );

    \I__2365\ : CascadeMux
    port map (
            O => \N__10129\,
            I => \N__10105\
        );

    \I__2364\ : Span4Mux_v
    port map (
            O => \N__10126\,
            I => \N__10099\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__10123\,
            I => \N__10094\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10120\,
            I => \N__10094\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__10117\,
            I => \N__10089\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__10114\,
            I => \N__10089\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10113\,
            I => \N__10086\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10112\,
            I => \N__10083\
        );

    \I__2357\ : InMux
    port map (
            O => \N__10111\,
            I => \N__10080\
        );

    \I__2356\ : InMux
    port map (
            O => \N__10110\,
            I => \N__10077\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10109\,
            I => \N__10074\
        );

    \I__2354\ : InMux
    port map (
            O => \N__10108\,
            I => \N__10057\
        );

    \I__2353\ : InMux
    port map (
            O => \N__10105\,
            I => \N__10057\
        );

    \I__2352\ : InMux
    port map (
            O => \N__10104\,
            I => \N__10057\
        );

    \I__2351\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10057\
        );

    \I__2350\ : InMux
    port map (
            O => \N__10102\,
            I => \N__10057\
        );

    \I__2349\ : Span4Mux_h
    port map (
            O => \N__10099\,
            I => \N__10052\
        );

    \I__2348\ : Span4Mux_v
    port map (
            O => \N__10094\,
            I => \N__10052\
        );

    \I__2347\ : Span4Mux_v
    port map (
            O => \N__10089\,
            I => \N__10047\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10086\,
            I => \N__10047\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10083\,
            I => \N__10038\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__10080\,
            I => \N__10038\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__10077\,
            I => \N__10038\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__10074\,
            I => \N__10038\
        );

    \I__2341\ : InMux
    port map (
            O => \N__10073\,
            I => \N__10029\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10072\,
            I => \N__10029\
        );

    \I__2339\ : InMux
    port map (
            O => \N__10071\,
            I => \N__10029\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10070\,
            I => \N__10029\
        );

    \I__2337\ : InMux
    port map (
            O => \N__10069\,
            I => \N__10026\
        );

    \I__2336\ : InMux
    port map (
            O => \N__10068\,
            I => \N__10023\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__10057\,
            I => \N__10020\
        );

    \I__2334\ : Span4Mux_h
    port map (
            O => \N__10052\,
            I => \N__10015\
        );

    \I__2333\ : Span4Mux_v
    port map (
            O => \N__10047\,
            I => \N__10015\
        );

    \I__2332\ : Span4Mux_v
    port map (
            O => \N__10038\,
            I => \N__10012\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__10029\,
            I => \N__10005\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__10026\,
            I => \N__10005\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10023\,
            I => \N__10005\
        );

    \I__2328\ : Span12Mux_v
    port map (
            O => \N__10020\,
            I => \N__9998\
        );

    \I__2327\ : Sp12to4
    port map (
            O => \N__10015\,
            I => \N__9998\
        );

    \I__2326\ : Sp12to4
    port map (
            O => \N__10012\,
            I => \N__9998\
        );

    \I__2325\ : Span12Mux_h
    port map (
            O => \N__10005\,
            I => \N__9995\
        );

    \I__2324\ : Span12Mux_h
    port map (
            O => \N__9998\,
            I => \N__9992\
        );

    \I__2323\ : Span12Mux_v
    port map (
            O => \N__9995\,
            I => \N__9989\
        );

    \I__2322\ : Span12Mux_v
    port map (
            O => \N__9992\,
            I => \N__9986\
        );

    \I__2321\ : Odrv12
    port map (
            O => \N__9989\,
            I => \AGNUS_REV_c\
        );

    \I__2320\ : Odrv12
    port map (
            O => \N__9986\,
            I => \AGNUS_REV_c\
        );

    \I__2319\ : InMux
    port map (
            O => \N__9981\,
            I => \N__9975\
        );

    \I__2318\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9975\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__9975\,
            I => \N__9972\
        );

    \I__2316\ : Odrv12
    port map (
            O => \N__9972\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2315\ : ClkMux
    port map (
            O => \N__9969\,
            I => \N__9951\
        );

    \I__2314\ : ClkMux
    port map (
            O => \N__9968\,
            I => \N__9951\
        );

    \I__2313\ : ClkMux
    port map (
            O => \N__9967\,
            I => \N__9951\
        );

    \I__2312\ : ClkMux
    port map (
            O => \N__9966\,
            I => \N__9951\
        );

    \I__2311\ : ClkMux
    port map (
            O => \N__9965\,
            I => \N__9951\
        );

    \I__2310\ : ClkMux
    port map (
            O => \N__9964\,
            I => \N__9951\
        );

    \I__2309\ : GlobalMux
    port map (
            O => \N__9951\,
            I => \N__9948\
        );

    \I__2308\ : gio2CtrlBuf
    port map (
            O => \N__9948\,
            I => \C3_c_g\
        );

    \I__2307\ : CEMux
    port map (
            O => \N__9945\,
            I => \N__9912\
        );

    \I__2306\ : CEMux
    port map (
            O => \N__9944\,
            I => \N__9912\
        );

    \I__2305\ : CEMux
    port map (
            O => \N__9943\,
            I => \N__9912\
        );

    \I__2304\ : CEMux
    port map (
            O => \N__9942\,
            I => \N__9912\
        );

    \I__2303\ : CEMux
    port map (
            O => \N__9941\,
            I => \N__9912\
        );

    \I__2302\ : CEMux
    port map (
            O => \N__9940\,
            I => \N__9912\
        );

    \I__2301\ : CEMux
    port map (
            O => \N__9939\,
            I => \N__9912\
        );

    \I__2300\ : CEMux
    port map (
            O => \N__9938\,
            I => \N__9912\
        );

    \I__2299\ : CEMux
    port map (
            O => \N__9937\,
            I => \N__9912\
        );

    \I__2298\ : CEMux
    port map (
            O => \N__9936\,
            I => \N__9912\
        );

    \I__2297\ : CEMux
    port map (
            O => \N__9935\,
            I => \N__9912\
        );

    \I__2296\ : GlobalMux
    port map (
            O => \N__9912\,
            I => \N__9909\
        );

    \I__2295\ : gio2CtrlBuf
    port map (
            O => \N__9909\,
            I => \DBRn_c_i_0_g\
        );

    \I__2294\ : InMux
    port map (
            O => \N__9906\,
            I => \N__9903\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__9903\,
            I => \N__9900\
        );

    \I__2292\ : Span12Mux_h
    port map (
            O => \N__9900\,
            I => \N__9897\
        );

    \I__2291\ : Odrv12
    port map (
            O => \N__9897\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2290\ : IoInMux
    port map (
            O => \N__9894\,
            I => \N__9891\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__9891\,
            I => \N__9888\
        );

    \I__2288\ : Span4Mux_s2_v
    port map (
            O => \N__9888\,
            I => \N__9885\
        );

    \I__2287\ : Span4Mux_v
    port map (
            O => \N__9885\,
            I => \N__9882\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__9882\,
            I => \N_257_i\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__9879\,
            I => \N__9874\
        );

    \I__2284\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9866\
        );

    \I__2283\ : InMux
    port map (
            O => \N__9877\,
            I => \N__9859\
        );

    \I__2282\ : InMux
    port map (
            O => \N__9874\,
            I => \N__9859\
        );

    \I__2281\ : InMux
    port map (
            O => \N__9873\,
            I => \N__9859\
        );

    \I__2280\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9854\
        );

    \I__2279\ : InMux
    port map (
            O => \N__9871\,
            I => \N__9854\
        );

    \I__2278\ : InMux
    port map (
            O => \N__9870\,
            I => \N__9849\
        );

    \I__2277\ : InMux
    port map (
            O => \N__9869\,
            I => \N__9849\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__9866\,
            I => \N__9844\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__9859\,
            I => \N__9844\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__9854\,
            I => \N__9841\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__9849\,
            I => \N__9838\
        );

    \I__2272\ : Sp12to4
    port map (
            O => \N__9844\,
            I => \N__9835\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__9841\,
            I => \N__9832\
        );

    \I__2270\ : Span4Mux_v
    port map (
            O => \N__9838\,
            I => \N__9829\
        );

    \I__2269\ : Span12Mux_v
    port map (
            O => \N__9835\,
            I => \N__9826\
        );

    \I__2268\ : Sp12to4
    port map (
            O => \N__9832\,
            I => \N__9821\
        );

    \I__2267\ : Sp12to4
    port map (
            O => \N__9829\,
            I => \N__9821\
        );

    \I__2266\ : Span12Mux_h
    port map (
            O => \N__9826\,
            I => \N__9818\
        );

    \I__2265\ : Span12Mux_h
    port map (
            O => \N__9821\,
            I => \N__9815\
        );

    \I__2264\ : Odrv12
    port map (
            O => \N__9818\,
            I => \A_c_1\
        );

    \I__2263\ : Odrv12
    port map (
            O => \N__9815\,
            I => \A_c_1\
        );

    \I__2262\ : InMux
    port map (
            O => \N__9810\,
            I => \N__9802\
        );

    \I__2261\ : InMux
    port map (
            O => \N__9809\,
            I => \N__9799\
        );

    \I__2260\ : InMux
    port map (
            O => \N__9808\,
            I => \N__9792\
        );

    \I__2259\ : InMux
    port map (
            O => \N__9807\,
            I => \N__9792\
        );

    \I__2258\ : InMux
    port map (
            O => \N__9806\,
            I => \N__9787\
        );

    \I__2257\ : InMux
    port map (
            O => \N__9805\,
            I => \N__9787\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__9802\,
            I => \N__9782\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__9799\,
            I => \N__9782\
        );

    \I__2254\ : InMux
    port map (
            O => \N__9798\,
            I => \N__9777\
        );

    \I__2253\ : InMux
    port map (
            O => \N__9797\,
            I => \N__9777\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__9792\,
            I => \N__9770\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__9787\,
            I => \N__9770\
        );

    \I__2250\ : Span4Mux_v
    port map (
            O => \N__9782\,
            I => \N__9767\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__9777\,
            I => \N__9764\
        );

    \I__2248\ : InMux
    port map (
            O => \N__9776\,
            I => \N__9759\
        );

    \I__2247\ : InMux
    port map (
            O => \N__9775\,
            I => \N__9759\
        );

    \I__2246\ : Span4Mux_h
    port map (
            O => \N__9770\,
            I => \N__9756\
        );

    \I__2245\ : Sp12to4
    port map (
            O => \N__9767\,
            I => \N__9751\
        );

    \I__2244\ : Sp12to4
    port map (
            O => \N__9764\,
            I => \N__9751\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__9759\,
            I => \N__9748\
        );

    \I__2242\ : Span4Mux_v
    port map (
            O => \N__9756\,
            I => \N__9745\
        );

    \I__2241\ : Span12Mux_v
    port map (
            O => \N__9751\,
            I => \N__9742\
        );

    \I__2240\ : Span12Mux_v
    port map (
            O => \N__9748\,
            I => \N__9739\
        );

    \I__2239\ : Span4Mux_h
    port map (
            O => \N__9745\,
            I => \N__9736\
        );

    \I__2238\ : Span12Mux_h
    port map (
            O => \N__9742\,
            I => \N__9733\
        );

    \I__2237\ : Span12Mux_v
    port map (
            O => \N__9739\,
            I => \N__9728\
        );

    \I__2236\ : Sp12to4
    port map (
            O => \N__9736\,
            I => \N__9728\
        );

    \I__2235\ : Odrv12
    port map (
            O => \N__9733\,
            I => \SIZ_c_0\
        );

    \I__2234\ : Odrv12
    port map (
            O => \N__9728\,
            I => \SIZ_c_0\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__9723\,
            I => \N__9719\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__9722\,
            I => \N__9716\
        );

    \I__2231\ : InMux
    port map (
            O => \N__9719\,
            I => \N__9708\
        );

    \I__2230\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9708\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__9715\,
            I => \N__9704\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__9714\,
            I => \N__9700\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__9713\,
            I => \N__9696\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__9708\,
            I => \N__9693\
        );

    \I__2225\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9688\
        );

    \I__2224\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9688\
        );

    \I__2223\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9685\
        );

    \I__2222\ : InMux
    port map (
            O => \N__9700\,
            I => \N__9678\
        );

    \I__2221\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9678\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9678\
        );

    \I__2219\ : Span4Mux_h
    port map (
            O => \N__9693\,
            I => \N__9673\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__9688\,
            I => \N__9673\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__9685\,
            I => \N__9668\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__9678\,
            I => \N__9668\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__9673\,
            I => \N__9663\
        );

    \I__2214\ : Sp12to4
    port map (
            O => \N__9668\,
            I => \N__9660\
        );

    \I__2213\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9655\
        );

    \I__2212\ : InMux
    port map (
            O => \N__9666\,
            I => \N__9655\
        );

    \I__2211\ : Sp12to4
    port map (
            O => \N__9663\,
            I => \N__9650\
        );

    \I__2210\ : Span12Mux_v
    port map (
            O => \N__9660\,
            I => \N__9650\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__9655\,
            I => \N__9647\
        );

    \I__2208\ : Span12Mux_h
    port map (
            O => \N__9650\,
            I => \N__9644\
        );

    \I__2207\ : Span12Mux_v
    port map (
            O => \N__9647\,
            I => \N__9641\
        );

    \I__2206\ : Odrv12
    port map (
            O => \N__9644\,
            I => \A_c_0\
        );

    \I__2205\ : Odrv12
    port map (
            O => \N__9641\,
            I => \A_c_0\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__9636\,
            I => \N__9633\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9633\,
            I => \N__9626\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9632\,
            I => \N__9623\
        );

    \I__2201\ : InMux
    port map (
            O => \N__9631\,
            I => \N__9618\
        );

    \I__2200\ : InMux
    port map (
            O => \N__9630\,
            I => \N__9618\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__9629\,
            I => \N__9613\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__9626\,
            I => \N__9609\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__9623\,
            I => \N__9604\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__9618\,
            I => \N__9604\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9599\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9616\,
            I => \N__9599\
        );

    \I__2193\ : InMux
    port map (
            O => \N__9613\,
            I => \N__9594\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9612\,
            I => \N__9594\
        );

    \I__2191\ : Span4Mux_v
    port map (
            O => \N__9609\,
            I => \N__9591\
        );

    \I__2190\ : Span4Mux_v
    port map (
            O => \N__9604\,
            I => \N__9588\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__9599\,
            I => \N__9583\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__9594\,
            I => \N__9583\
        );

    \I__2187\ : Sp12to4
    port map (
            O => \N__9591\,
            I => \N__9578\
        );

    \I__2186\ : Sp12to4
    port map (
            O => \N__9588\,
            I => \N__9578\
        );

    \I__2185\ : Sp12to4
    port map (
            O => \N__9583\,
            I => \N__9575\
        );

    \I__2184\ : Span12Mux_h
    port map (
            O => \N__9578\,
            I => \N__9572\
        );

    \I__2183\ : Span12Mux_v
    port map (
            O => \N__9575\,
            I => \N__9569\
        );

    \I__2182\ : Span12Mux_v
    port map (
            O => \N__9572\,
            I => \N__9564\
        );

    \I__2181\ : Span12Mux_h
    port map (
            O => \N__9569\,
            I => \N__9564\
        );

    \I__2180\ : Odrv12
    port map (
            O => \N__9564\,
            I => \SIZ_c_1\
        );

    \I__2179\ : IoInMux
    port map (
            O => \N__9561\,
            I => \N__9558\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9558\,
            I => \N__9555\
        );

    \I__2177\ : Span4Mux_s2_v
    port map (
            O => \N__9555\,
            I => \N__9552\
        );

    \I__2176\ : Span4Mux_h
    port map (
            O => \N__9552\,
            I => \N__9549\
        );

    \I__2175\ : Span4Mux_v
    port map (
            O => \N__9549\,
            I => \N__9546\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__9546\,
            I => \N_258_i\
        );

    \I__2173\ : IoInMux
    port map (
            O => \N__9543\,
            I => \N__9540\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9540\,
            I => \N__9537\
        );

    \I__2171\ : Span4Mux_s2_v
    port map (
            O => \N__9537\,
            I => \N__9534\
        );

    \I__2170\ : Span4Mux_h
    port map (
            O => \N__9534\,
            I => \N__9531\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__9531\,
            I => \CRCSn_c\
        );

    \I__2168\ : IoInMux
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9525\,
            I => \N__9522\
        );

    \I__2166\ : Span12Mux_s7_v
    port map (
            O => \N__9522\,
            I => \N__9519\
        );

    \I__2165\ : Odrv12
    port map (
            O => \N__9519\,
            I => \RASn_c\
        );

    \I__2164\ : IoInMux
    port map (
            O => \N__9516\,
            I => \N__9513\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__9513\,
            I => \N__9510\
        );

    \I__2162\ : Span4Mux_s2_v
    port map (
            O => \N__9510\,
            I => \N__9507\
        );

    \I__2161\ : Span4Mux_v
    port map (
            O => \N__9507\,
            I => \N__9504\
        );

    \I__2160\ : Span4Mux_h
    port map (
            O => \N__9504\,
            I => \N__9501\
        );

    \I__2159\ : Span4Mux_h
    port map (
            O => \N__9501\,
            I => \N__9498\
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__9498\,
            I => \CASn_c\
        );

    \I__2157\ : IoInMux
    port map (
            O => \N__9495\,
            I => \N__9492\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__9492\,
            I => \N__9489\
        );

    \I__2155\ : Span4Mux_s1_h
    port map (
            O => \N__9489\,
            I => \N__9486\
        );

    \I__2154\ : Sp12to4
    port map (
            O => \N__9486\,
            I => \N__9483\
        );

    \I__2153\ : Span12Mux_s6_v
    port map (
            O => \N__9483\,
            I => \N__9480\
        );

    \I__2152\ : Span12Mux_h
    port map (
            O => \N__9480\,
            I => \N__9477\
        );

    \I__2151\ : Odrv12
    port map (
            O => \N__9477\,
            I => \WEn_c\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9474\,
            I => \N__9471\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__9471\,
            I => \N__9467\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9470\,
            I => \N__9464\
        );

    \I__2147\ : Span4Mux_v
    port map (
            O => \N__9467\,
            I => \N__9458\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__9464\,
            I => \N__9458\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9463\,
            I => \N__9455\
        );

    \I__2144\ : Span4Mux_v
    port map (
            O => \N__9458\,
            I => \N__9451\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9455\,
            I => \N__9445\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9454\,
            I => \N__9442\
        );

    \I__2141\ : Span4Mux_h
    port map (
            O => \N__9451\,
            I => \N__9439\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9450\,
            I => \N__9436\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9433\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9448\,
            I => \N__9430\
        );

    \I__2137\ : Span4Mux_h
    port map (
            O => \N__9445\,
            I => \N__9427\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9442\,
            I => \N__9424\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__9439\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9436\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__9433\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9430\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2131\ : Odrv4
    port map (
            O => \N__9427\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__9424\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__9411\,
            I => \N__9404\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9400\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9397\
        );

    \I__2126\ : CascadeMux
    port map (
            O => \N__9408\,
            I => \N__9393\
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__9407\,
            I => \N__9388\
        );

    \I__2124\ : InMux
    port map (
            O => \N__9404\,
            I => \N__9384\
        );

    \I__2123\ : CascadeMux
    port map (
            O => \N__9403\,
            I => \N__9380\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9400\,
            I => \N__9375\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__9397\,
            I => \N__9375\
        );

    \I__2120\ : InMux
    port map (
            O => \N__9396\,
            I => \N__9372\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9365\
        );

    \I__2118\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9365\
        );

    \I__2117\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9365\
        );

    \I__2116\ : InMux
    port map (
            O => \N__9388\,
            I => \N__9359\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__9387\,
            I => \N__9355\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__9384\,
            I => \N__9352\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9383\,
            I => \N__9349\
        );

    \I__2112\ : InMux
    port map (
            O => \N__9380\,
            I => \N__9346\
        );

    \I__2111\ : Span4Mux_v
    port map (
            O => \N__9375\,
            I => \N__9339\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9372\,
            I => \N__9339\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__9365\,
            I => \N__9339\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9364\,
            I => \N__9325\
        );

    \I__2107\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9325\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9322\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__9359\,
            I => \N__9319\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9316\
        );

    \I__2103\ : InMux
    port map (
            O => \N__9355\,
            I => \N__9313\
        );

    \I__2102\ : Span4Mux_h
    port map (
            O => \N__9352\,
            I => \N__9310\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9349\,
            I => \N__9305\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__9346\,
            I => \N__9305\
        );

    \I__2099\ : Span4Mux_h
    port map (
            O => \N__9339\,
            I => \N__9302\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9295\
        );

    \I__2097\ : InMux
    port map (
            O => \N__9337\,
            I => \N__9295\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9336\,
            I => \N__9295\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9284\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9284\
        );

    \I__2093\ : InMux
    port map (
            O => \N__9333\,
            I => \N__9284\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9284\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9331\,
            I => \N__9284\
        );

    \I__2090\ : InMux
    port map (
            O => \N__9330\,
            I => \N__9281\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__9325\,
            I => \N__9274\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__9322\,
            I => \N__9274\
        );

    \I__2087\ : Span4Mux_h
    port map (
            O => \N__9319\,
            I => \N__9274\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9316\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__9313\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__9310\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__9305\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2082\ : Odrv4
    port map (
            O => \N__9302\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__9295\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9284\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__9281\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__9274\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9255\,
            I => \N__9251\
        );

    \I__2076\ : CascadeMux
    port map (
            O => \N__9254\,
            I => \N__9248\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__9251\,
            I => \N__9245\
        );

    \I__2074\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9242\
        );

    \I__2073\ : Span4Mux_v
    port map (
            O => \N__9245\,
            I => \N__9235\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__9242\,
            I => \N__9235\
        );

    \I__2071\ : InMux
    port map (
            O => \N__9241\,
            I => \N__9232\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__9240\,
            I => \N__9229\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__9235\,
            I => \N__9226\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__9232\,
            I => \N__9223\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9229\,
            I => \N__9220\
        );

    \I__2066\ : Span4Mux_h
    port map (
            O => \N__9226\,
            I => \N__9215\
        );

    \I__2065\ : Span4Mux_v
    port map (
            O => \N__9223\,
            I => \N__9215\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__9220\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__9215\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2062\ : InMux
    port map (
            O => \N__9210\,
            I => \N__9206\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9209\,
            I => \N__9203\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__9206\,
            I => \N__9195\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__9203\,
            I => \N__9195\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9202\,
            I => \N__9191\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9201\,
            I => \N__9188\
        );

    \I__2056\ : CascadeMux
    port map (
            O => \N__9200\,
            I => \N__9185\
        );

    \I__2055\ : Span4Mux_v
    port map (
            O => \N__9195\,
            I => \N__9182\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9194\,
            I => \N__9179\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9191\,
            I => \N__9176\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__9188\,
            I => \N__9172\
        );

    \I__2051\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9169\
        );

    \I__2050\ : Span4Mux_h
    port map (
            O => \N__9182\,
            I => \N__9164\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9179\,
            I => \N__9164\
        );

    \I__2048\ : Span4Mux_h
    port map (
            O => \N__9176\,
            I => \N__9161\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9175\,
            I => \N__9158\
        );

    \I__2046\ : Span4Mux_v
    port map (
            O => \N__9172\,
            I => \N__9155\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__9169\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__9164\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__9161\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9158\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__9155\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2040\ : IoInMux
    port map (
            O => \N__9144\,
            I => \N__9141\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__9141\,
            I => \N__9138\
        );

    \I__2038\ : Span4Mux_s3_v
    port map (
            O => \N__9138\,
            I => \N__9135\
        );

    \I__2037\ : Span4Mux_v
    port map (
            O => \N__9135\,
            I => \N__9132\
        );

    \I__2036\ : Span4Mux_h
    port map (
            O => \N__9132\,
            I => \N__9129\
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__9129\,
            I => \CMA_c_10\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9126\,
            I => \N__9123\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9123\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9120\,
            I => \N__9116\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__9119\,
            I => \N__9113\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9116\,
            I => \N__9110\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9113\,
            I => \N__9107\
        );

    \I__2028\ : Span4Mux_h
    port map (
            O => \N__9110\,
            I => \N__9104\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__9107\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2026\ : Odrv4
    port map (
            O => \N__9104\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9096\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9096\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2023\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9090\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__9090\,
            I => \N__9087\
        );

    \I__2021\ : Odrv4
    port map (
            O => \N__9087\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9076\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9083\,
            I => \N__9076\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9082\,
            I => \N__9071\
        );

    \I__2017\ : InMux
    port map (
            O => \N__9081\,
            I => \N__9071\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9076\,
            I => \N__9066\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9071\,
            I => \N__9066\
        );

    \I__2014\ : Span12Mux_v
    port map (
            O => \N__9066\,
            I => \N__9063\
        );

    \I__2013\ : Span12Mux_h
    port map (
            O => \N__9063\,
            I => \N__9060\
        );

    \I__2012\ : Odrv12
    port map (
            O => \N__9060\,
            I => \DRA_c_2\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__9057\,
            I => \N__9054\
        );

    \I__2010\ : InMux
    port map (
            O => \N__9054\,
            I => \N__9051\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__9051\,
            I => \N__9048\
        );

    \I__2008\ : Span4Mux_v
    port map (
            O => \N__9048\,
            I => \N__9045\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__9045\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2006\ : InMux
    port map (
            O => \N__9042\,
            I => \N__9039\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__9039\,
            I => \N__9036\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__9036\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9033\,
            I => \N__9030\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9030\,
            I => \N__9027\
        );

    \I__2001\ : Span4Mux_h
    port map (
            O => \N__9027\,
            I => \N__9024\
        );

    \I__2000\ : Odrv4
    port map (
            O => \N__9024\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__9021\,
            I => \N__9018\
        );

    \I__1998\ : InMux
    port map (
            O => \N__9018\,
            I => \N__9015\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__9015\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1996\ : InMux
    port map (
            O => \N__9012\,
            I => \N__9006\
        );

    \I__1995\ : InMux
    port map (
            O => \N__9011\,
            I => \N__9006\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__9006\,
            I => \N__9002\
        );

    \I__1993\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8999\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__9002\,
            I => \N__8993\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__8999\,
            I => \N__8993\
        );

    \I__1990\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8990\
        );

    \I__1989\ : Span4Mux_h
    port map (
            O => \N__8993\,
            I => \N__8987\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__8990\,
            I => \N__8984\
        );

    \I__1987\ : Sp12to4
    port map (
            O => \N__8987\,
            I => \N__8981\
        );

    \I__1986\ : Span12Mux_v
    port map (
            O => \N__8984\,
            I => \N__8978\
        );

    \I__1985\ : Span12Mux_v
    port map (
            O => \N__8981\,
            I => \N__8975\
        );

    \I__1984\ : Span12Mux_h
    port map (
            O => \N__8978\,
            I => \N__8972\
        );

    \I__1983\ : Odrv12
    port map (
            O => \N__8975\,
            I => \DRA_c_3\
        );

    \I__1982\ : Odrv12
    port map (
            O => \N__8972\,
            I => \DRA_c_3\
        );

    \I__1981\ : InMux
    port map (
            O => \N__8967\,
            I => \N__8960\
        );

    \I__1980\ : InMux
    port map (
            O => \N__8966\,
            I => \N__8960\
        );

    \I__1979\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8957\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__8960\,
            I => \N__8953\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__8957\,
            I => \N__8950\
        );

    \I__1976\ : InMux
    port map (
            O => \N__8956\,
            I => \N__8947\
        );

    \I__1975\ : Span4Mux_v
    port map (
            O => \N__8953\,
            I => \N__8940\
        );

    \I__1974\ : Span4Mux_h
    port map (
            O => \N__8950\,
            I => \N__8940\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__8947\,
            I => \N__8940\
        );

    \I__1972\ : Span4Mux_v
    port map (
            O => \N__8940\,
            I => \N__8937\
        );

    \I__1971\ : Span4Mux_v
    port map (
            O => \N__8937\,
            I => \N__8934\
        );

    \I__1970\ : Sp12to4
    port map (
            O => \N__8934\,
            I => \N__8931\
        );

    \I__1969\ : Span12Mux_h
    port map (
            O => \N__8931\,
            I => \N__8928\
        );

    \I__1968\ : Odrv12
    port map (
            O => \N__8928\,
            I => \DRA_c_4\
        );

    \I__1967\ : InMux
    port map (
            O => \N__8925\,
            I => \N__8922\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__8922\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1965\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8916\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__8916\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8910\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__8910\,
            I => \N__8907\
        );

    \I__1961\ : Odrv12
    port map (
            O => \N__8907\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1960\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8901\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__8901\,
            I => \N__8898\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__8898\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1957\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8891\
        );

    \I__1956\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8888\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__8891\,
            I => \N__8885\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__8888\,
            I => \N__8882\
        );

    \I__1953\ : Span12Mux_h
    port map (
            O => \N__8885\,
            I => \N__8879\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__8882\,
            I => \N__8876\
        );

    \I__1951\ : Odrv12
    port map (
            O => \N__8879\,
            I => \DBRn_c_i\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__8876\,
            I => \DBRn_c_i\
        );

    \I__1949\ : InMux
    port map (
            O => \N__8871\,
            I => \N__8868\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__8868\,
            I => \N__8865\
        );

    \I__1947\ : Span4Mux_h
    port map (
            O => \N__8865\,
            I => \N__8861\
        );

    \I__1946\ : InMux
    port map (
            O => \N__8864\,
            I => \N__8858\
        );

    \I__1945\ : Span4Mux_h
    port map (
            O => \N__8861\,
            I => \N__8855\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__8858\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__8855\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__1942\ : IoInMux
    port map (
            O => \N__8850\,
            I => \N__8847\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__8847\,
            I => \N__8844\
        );

    \I__1940\ : Span4Mux_s2_v
    port map (
            O => \N__8844\,
            I => \N__8841\
        );

    \I__1939\ : Span4Mux_v
    port map (
            O => \N__8841\,
            I => \N__8838\
        );

    \I__1938\ : Odrv4
    port map (
            O => \N__8838\,
            I => \N_260_i\
        );

    \I__1937\ : IoInMux
    port map (
            O => \N__8835\,
            I => \N__8832\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8832\,
            I => \N__8829\
        );

    \I__1935\ : Span4Mux_s2_v
    port map (
            O => \N__8829\,
            I => \N__8826\
        );

    \I__1934\ : Span4Mux_v
    port map (
            O => \N__8826\,
            I => \N__8823\
        );

    \I__1933\ : Odrv4
    port map (
            O => \N__8823\,
            I => \N_259_i\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8820\,
            I => \N__8812\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8819\,
            I => \N__8805\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8818\,
            I => \N__8805\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8817\,
            I => \N__8805\
        );

    \I__1928\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8802\
        );

    \I__1927\ : InMux
    port map (
            O => \N__8815\,
            I => \N__8799\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__8812\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__8805\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8802\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__8799\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__8790\,
            I => \N__8784\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__8789\,
            I => \N__8779\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__8788\,
            I => \N__8776\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__8787\,
            I => \N__8773\
        );

    \I__1918\ : InMux
    port map (
            O => \N__8784\,
            I => \N__8770\
        );

    \I__1917\ : InMux
    port map (
            O => \N__8783\,
            I => \N__8763\
        );

    \I__1916\ : InMux
    port map (
            O => \N__8782\,
            I => \N__8763\
        );

    \I__1915\ : InMux
    port map (
            O => \N__8779\,
            I => \N__8760\
        );

    \I__1914\ : InMux
    port map (
            O => \N__8776\,
            I => \N__8757\
        );

    \I__1913\ : InMux
    port map (
            O => \N__8773\,
            I => \N__8754\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__8770\,
            I => \N__8751\
        );

    \I__1911\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8748\
        );

    \I__1910\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8745\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__8763\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8760\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8757\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__8754\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1905\ : Odrv4
    port map (
            O => \N__8751\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8748\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__8745\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8730\,
            I => \N__8727\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__8727\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1900\ : IoInMux
    port map (
            O => \N__8724\,
            I => \N__8721\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__8721\,
            I => \N__8718\
        );

    \I__1898\ : Span4Mux_s2_v
    port map (
            O => \N__8718\,
            I => \N__8715\
        );

    \I__1897\ : Span4Mux_v
    port map (
            O => \N__8715\,
            I => \N__8712\
        );

    \I__1896\ : Span4Mux_v
    port map (
            O => \N__8712\,
            I => \N__8709\
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__8709\,
            I => \CMA_c_0\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8703\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__8703\,
            I => \N__8700\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__8700\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1891\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8694\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__8694\,
            I => \N__8691\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__8691\,
            I => \N__8688\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__8688\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1887\ : IoInMux
    port map (
            O => \N__8685\,
            I => \N__8682\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__8682\,
            I => \N__8679\
        );

    \I__1885\ : IoSpan4Mux
    port map (
            O => \N__8679\,
            I => \N__8676\
        );

    \I__1884\ : Sp12to4
    port map (
            O => \N__8676\,
            I => \N__8673\
        );

    \I__1883\ : Odrv12
    port map (
            O => \N__8673\,
            I => \CMA_c_2\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8670\,
            I => \N__8667\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__8667\,
            I => \N__8664\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__8664\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8661\,
            I => \N__8658\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8658\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1877\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8652\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8652\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1875\ : IoInMux
    port map (
            O => \N__8649\,
            I => \N__8646\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__8646\,
            I => \N__8643\
        );

    \I__1873\ : IoSpan4Mux
    port map (
            O => \N__8643\,
            I => \N__8640\
        );

    \I__1872\ : Sp12to4
    port map (
            O => \N__8640\,
            I => \N__8637\
        );

    \I__1871\ : Span12Mux_s9_v
    port map (
            O => \N__8637\,
            I => \N__8634\
        );

    \I__1870\ : Span12Mux_h
    port map (
            O => \N__8634\,
            I => \N__8631\
        );

    \I__1869\ : Odrv12
    port map (
            O => \N__8631\,
            I => \CMA_c_4\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8628\,
            I => \N__8625\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8625\,
            I => \N__8622\
        );

    \I__1866\ : Span4Mux_v
    port map (
            O => \N__8622\,
            I => \N__8619\
        );

    \I__1865\ : Odrv4
    port map (
            O => \N__8619\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__8616\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_\
        );

    \I__1863\ : IoInMux
    port map (
            O => \N__8613\,
            I => \N__8610\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8610\,
            I => \N__8607\
        );

    \I__1861\ : IoSpan4Mux
    port map (
            O => \N__8607\,
            I => \N__8604\
        );

    \I__1860\ : Span4Mux_s3_h
    port map (
            O => \N__8604\,
            I => \N__8601\
        );

    \I__1859\ : Sp12to4
    port map (
            O => \N__8601\,
            I => \N__8598\
        );

    \I__1858\ : Span12Mux_s11_v
    port map (
            O => \N__8598\,
            I => \N__8595\
        );

    \I__1857\ : Odrv12
    port map (
            O => \N__8595\,
            I => \CMA_c_7\
        );

    \I__1856\ : IoInMux
    port map (
            O => \N__8592\,
            I => \N__8589\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__8589\,
            I => \N__8586\
        );

    \I__1854\ : IoSpan4Mux
    port map (
            O => \N__8586\,
            I => \N__8583\
        );

    \I__1853\ : Span4Mux_s1_h
    port map (
            O => \N__8583\,
            I => \N__8580\
        );

    \I__1852\ : Sp12to4
    port map (
            O => \N__8580\,
            I => \N__8577\
        );

    \I__1851\ : Span12Mux_h
    port map (
            O => \N__8577\,
            I => \N__8574\
        );

    \I__1850\ : Odrv12
    port map (
            O => \N__8574\,
            I => \CMA_c_6\
        );

    \I__1849\ : InMux
    port map (
            O => \N__8571\,
            I => \N__8568\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8568\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8565\,
            I => \N__8562\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__8562\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1845\ : InMux
    port map (
            O => \N__8559\,
            I => \N__8556\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__8556\,
            I => \N__8553\
        );

    \I__1843\ : Span4Mux_v
    port map (
            O => \N__8553\,
            I => \N__8550\
        );

    \I__1842\ : Sp12to4
    port map (
            O => \N__8550\,
            I => \N__8547\
        );

    \I__1841\ : Span12Mux_h
    port map (
            O => \N__8547\,
            I => \N__8544\
        );

    \I__1840\ : Odrv12
    port map (
            O => \N__8544\,
            I => \A_c_12\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8541\,
            I => \N__8538\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8538\,
            I => \N__8535\
        );

    \I__1837\ : Span12Mux_v
    port map (
            O => \N__8535\,
            I => \N__8532\
        );

    \I__1836\ : Span12Mux_h
    port map (
            O => \N__8532\,
            I => \N__8529\
        );

    \I__1835\ : Odrv12
    port map (
            O => \N__8529\,
            I => \A_c_5\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__8526\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8523\,
            I => \N__8520\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8520\,
            I => \N__8517\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__8517\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1830\ : InMux
    port map (
            O => \N__8514\,
            I => \N__8511\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__8511\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8508\,
            I => \N__8505\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8505\,
            I => \N__8502\
        );

    \I__1826\ : Span4Mux_v
    port map (
            O => \N__8502\,
            I => \N__8499\
        );

    \I__1825\ : Span4Mux_v
    port map (
            O => \N__8499\,
            I => \N__8496\
        );

    \I__1824\ : Sp12to4
    port map (
            O => \N__8496\,
            I => \N__8493\
        );

    \I__1823\ : Span12Mux_h
    port map (
            O => \N__8493\,
            I => \N__8490\
        );

    \I__1822\ : Odrv12
    port map (
            O => \N__8490\,
            I => \A_c_4\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8487\,
            I => \N__8484\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8484\,
            I => \N__8481\
        );

    \I__1819\ : Span12Mux_v
    port map (
            O => \N__8481\,
            I => \N__8478\
        );

    \I__1818\ : Span12Mux_h
    port map (
            O => \N__8478\,
            I => \N__8475\
        );

    \I__1817\ : Odrv12
    port map (
            O => \N__8475\,
            I => \A_c_11\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8472\,
            I => \N__8466\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8471\,
            I => \N__8463\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__8470\,
            I => \N__8460\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8469\,
            I => \N__8456\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8466\,
            I => \N__8452\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8463\,
            I => \N__8449\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8460\,
            I => \N__8443\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8443\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8456\,
            I => \N__8440\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8437\
        );

    \I__1806\ : Span4Mux_h
    port map (
            O => \N__8452\,
            I => \N__8432\
        );

    \I__1805\ : Span4Mux_h
    port map (
            O => \N__8449\,
            I => \N__8432\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8448\,
            I => \N__8429\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8443\,
            I => \N__8426\
        );

    \I__1802\ : Odrv12
    port map (
            O => \N__8440\,
            I => \DMA_CYCLE\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8437\,
            I => \DMA_CYCLE\
        );

    \I__1800\ : Odrv4
    port map (
            O => \N__8432\,
            I => \DMA_CYCLE\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8429\,
            I => \DMA_CYCLE\
        );

    \I__1798\ : Odrv4
    port map (
            O => \N__8426\,
            I => \DMA_CYCLE\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8415\,
            I => \N__8412\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8412\,
            I => \N__8409\
        );

    \I__1795\ : Odrv12
    port map (
            O => \N__8409\,
            I => \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_0Z0Z_0\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__8406\,
            I => \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_0Z0Z_0_cascade_\
        );

    \I__1793\ : IoInMux
    port map (
            O => \N__8403\,
            I => \N__8400\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__8400\,
            I => \N__8395\
        );

    \I__1791\ : CascadeMux
    port map (
            O => \N__8399\,
            I => \N__8391\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__8398\,
            I => \N__8388\
        );

    \I__1789\ : Span4Mux_s3_v
    port map (
            O => \N__8395\,
            I => \N__8385\
        );

    \I__1788\ : InMux
    port map (
            O => \N__8394\,
            I => \N__8382\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8391\,
            I => \N__8379\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8388\,
            I => \N__8376\
        );

    \I__1785\ : Span4Mux_v
    port map (
            O => \N__8385\,
            I => \N__8372\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8382\,
            I => \N__8369\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8379\,
            I => \N__8364\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8376\,
            I => \N__8364\
        );

    \I__1781\ : InMux
    port map (
            O => \N__8375\,
            I => \N__8361\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__8372\,
            I => \N__8358\
        );

    \I__1779\ : Span4Mux_v
    port map (
            O => \N__8369\,
            I => \N__8351\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__8364\,
            I => \N__8351\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__8361\,
            I => \N__8351\
        );

    \I__1776\ : Span4Mux_h
    port map (
            O => \N__8358\,
            I => \N__8345\
        );

    \I__1775\ : Span4Mux_h
    port map (
            O => \N__8351\,
            I => \N__8345\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8342\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__8345\,
            I => \DBENn_c\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8342\,
            I => \DBENn_c\
        );

    \I__1771\ : IoInMux
    port map (
            O => \N__8337\,
            I => \N__8334\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8334\,
            I => \N__8331\
        );

    \I__1769\ : Span12Mux_s4_h
    port map (
            O => \N__8331\,
            I => \N__8328\
        );

    \I__1768\ : Span12Mux_h
    port map (
            O => \N__8328\,
            I => \N__8325\
        );

    \I__1767\ : Odrv12
    port map (
            O => \N__8325\,
            I => \N_203_i\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8322\,
            I => \N__8316\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8316\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8316\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8313\,
            I => \N__8310\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__8310\,
            I => \N__8307\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__8307\,
            I => \U712_BYTE_ENABLE.N_260\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__8304\,
            I => \N__8299\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__8303\,
            I => \N__8296\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__8302\,
            I => \N__8290\
        );

    \I__1757\ : InMux
    port map (
            O => \N__8299\,
            I => \N__8284\
        );

    \I__1756\ : InMux
    port map (
            O => \N__8296\,
            I => \N__8279\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8295\,
            I => \N__8279\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8294\,
            I => \N__8276\
        );

    \I__1753\ : InMux
    port map (
            O => \N__8293\,
            I => \N__8269\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8290\,
            I => \N__8269\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8289\,
            I => \N__8269\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8288\,
            I => \N__8266\
        );

    \I__1749\ : InMux
    port map (
            O => \N__8287\,
            I => \N__8262\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8284\,
            I => \N__8251\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8279\,
            I => \N__8251\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__8276\,
            I => \N__8251\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8269\,
            I => \N__8246\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__8266\,
            I => \N__8246\
        );

    \I__1743\ : InMux
    port map (
            O => \N__8265\,
            I => \N__8243\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__8262\,
            I => \N__8237\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8234\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8260\,
            I => \N__8227\
        );

    \I__1739\ : InMux
    port map (
            O => \N__8259\,
            I => \N__8227\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8258\,
            I => \N__8227\
        );

    \I__1737\ : Span4Mux_h
    port map (
            O => \N__8251\,
            I => \N__8224\
        );

    \I__1736\ : Span4Mux_v
    port map (
            O => \N__8246\,
            I => \N__8219\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8243\,
            I => \N__8219\
        );

    \I__1734\ : InMux
    port map (
            O => \N__8242\,
            I => \N__8216\
        );

    \I__1733\ : InMux
    port map (
            O => \N__8241\,
            I => \N__8213\
        );

    \I__1732\ : InMux
    port map (
            O => \N__8240\,
            I => \N__8209\
        );

    \I__1731\ : Span4Mux_v
    port map (
            O => \N__8237\,
            I => \N__8201\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__8234\,
            I => \N__8201\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8227\,
            I => \N__8201\
        );

    \I__1728\ : Span4Mux_v
    port map (
            O => \N__8224\,
            I => \N__8192\
        );

    \I__1727\ : Span4Mux_h
    port map (
            O => \N__8219\,
            I => \N__8192\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__8216\,
            I => \N__8192\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8213\,
            I => \N__8192\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8189\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8209\,
            I => \N__8186\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8208\,
            I => \N__8183\
        );

    \I__1721\ : Span4Mux_v
    port map (
            O => \N__8201\,
            I => \N__8180\
        );

    \I__1720\ : Sp12to4
    port map (
            O => \N__8192\,
            I => \N__8175\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8189\,
            I => \N__8175\
        );

    \I__1718\ : Span12Mux_v
    port map (
            O => \N__8186\,
            I => \N__8170\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8183\,
            I => \N__8170\
        );

    \I__1716\ : Sp12to4
    port map (
            O => \N__8180\,
            I => \N__8165\
        );

    \I__1715\ : Span12Mux_v
    port map (
            O => \N__8175\,
            I => \N__8165\
        );

    \I__1714\ : Span12Mux_h
    port map (
            O => \N__8170\,
            I => \N__8162\
        );

    \I__1713\ : Span12Mux_h
    port map (
            O => \N__8165\,
            I => \N__8159\
        );

    \I__1712\ : Odrv12
    port map (
            O => \N__8162\,
            I => \RESETn_c\
        );

    \I__1711\ : Odrv12
    port map (
            O => \N__8159\,
            I => \RESETn_c\
        );

    \I__1710\ : IoInMux
    port map (
            O => \N__8154\,
            I => \N__8151\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__8151\,
            I => \N__8147\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8150\,
            I => \N__8144\
        );

    \I__1707\ : Span12Mux_s9_v
    port map (
            O => \N__8147\,
            I => \N__8141\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8144\,
            I => \N__8138\
        );

    \I__1705\ : Odrv12
    port map (
            O => \N__8141\,
            I => \RESETn_c_i\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__8138\,
            I => \RESETn_c_i\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__8133\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8130\,
            I => \N__8127\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8127\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1700\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8121\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__8121\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__1698\ : IoInMux
    port map (
            O => \N__8118\,
            I => \N__8115\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__8115\,
            I => \N__8112\
        );

    \I__1696\ : IoSpan4Mux
    port map (
            O => \N__8112\,
            I => \N__8109\
        );

    \I__1695\ : Span4Mux_s2_h
    port map (
            O => \N__8109\,
            I => \N__8106\
        );

    \I__1694\ : Sp12to4
    port map (
            O => \N__8106\,
            I => \N__8103\
        );

    \I__1693\ : Span12Mux_h
    port map (
            O => \N__8103\,
            I => \N__8100\
        );

    \I__1692\ : Odrv12
    port map (
            O => \N__8100\,
            I => \CMA_c_5\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8094\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__8094\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8088\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8088\,
            I => \N__8085\
        );

    \I__1687\ : Span4Mux_v
    port map (
            O => \N__8085\,
            I => \N__8082\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__8082\,
            I => \U712_BYTE_ENABLE.N_259\
        );

    \I__1685\ : IoInMux
    port map (
            O => \N__8079\,
            I => \N__8076\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__8076\,
            I => \N__8073\
        );

    \I__1683\ : IoSpan4Mux
    port map (
            O => \N__8073\,
            I => \N__8070\
        );

    \I__1682\ : Span4Mux_s2_h
    port map (
            O => \N__8070\,
            I => \N__8067\
        );

    \I__1681\ : Sp12to4
    port map (
            O => \N__8067\,
            I => \N__8064\
        );

    \I__1680\ : Span12Mux_h
    port map (
            O => \N__8064\,
            I => \N__8061\
        );

    \I__1679\ : Odrv12
    port map (
            O => \N__8061\,
            I => \N_222_i\
        );

    \I__1678\ : InMux
    port map (
            O => \N__8058\,
            I => \N__8055\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__8055\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__8052\,
            I => \N__8049\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8049\,
            I => \N__8043\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8048\,
            I => \N__8043\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__8043\,
            I => \N__8040\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__8040\,
            I => \N__8037\
        );

    \I__1671\ : Span4Mux_v
    port map (
            O => \N__8037\,
            I => \N__8034\
        );

    \I__1670\ : Sp12to4
    port map (
            O => \N__8034\,
            I => \N__8031\
        );

    \I__1669\ : Span12Mux_h
    port map (
            O => \N__8031\,
            I => \N__8028\
        );

    \I__1668\ : Odrv12
    port map (
            O => \N__8028\,
            I => \A_c_14\
        );

    \I__1667\ : InMux
    port map (
            O => \N__8025\,
            I => \N__8022\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__8022\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1665\ : InMux
    port map (
            O => \N__8019\,
            I => \N__8015\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__8018\,
            I => \N__8012\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__8015\,
            I => \N__8009\
        );

    \I__1662\ : InMux
    port map (
            O => \N__8012\,
            I => \N__8006\
        );

    \I__1661\ : Odrv4
    port map (
            O => \N__8009\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__8006\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8001\,
            I => \N__7998\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__7998\,
            I => \N__7995\
        );

    \I__1657\ : Span4Mux_h
    port map (
            O => \N__7995\,
            I => \N__7992\
        );

    \I__1656\ : Span4Mux_v
    port map (
            O => \N__7992\,
            I => \N__7989\
        );

    \I__1655\ : Sp12to4
    port map (
            O => \N__7989\,
            I => \N__7986\
        );

    \I__1654\ : Span12Mux_h
    port map (
            O => \N__7986\,
            I => \N__7983\
        );

    \I__1653\ : Odrv12
    port map (
            O => \N__7983\,
            I => \A_c_8\
        );

    \I__1652\ : InMux
    port map (
            O => \N__7980\,
            I => \N__7977\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__7977\,
            I => \N__7974\
        );

    \I__1650\ : Span12Mux_v
    port map (
            O => \N__7974\,
            I => \N__7971\
        );

    \I__1649\ : Span12Mux_h
    port map (
            O => \N__7971\,
            I => \N__7968\
        );

    \I__1648\ : Odrv12
    port map (
            O => \N__7968\,
            I => \A_c_15\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7962\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__7962\,
            I => \N__7959\
        );

    \I__1645\ : Span12Mux_v
    port map (
            O => \N__7959\,
            I => \N__7956\
        );

    \I__1644\ : Span12Mux_h
    port map (
            O => \N__7956\,
            I => \N__7953\
        );

    \I__1643\ : Span12Mux_v
    port map (
            O => \N__7953\,
            I => \N__7950\
        );

    \I__1642\ : Odrv12
    port map (
            O => \N__7950\,
            I => \A_c_2\
        );

    \I__1641\ : InMux
    port map (
            O => \N__7947\,
            I => \N__7944\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__7944\,
            I => \N__7941\
        );

    \I__1639\ : Span4Mux_v
    port map (
            O => \N__7941\,
            I => \N__7938\
        );

    \I__1638\ : Sp12to4
    port map (
            O => \N__7938\,
            I => \N__7935\
        );

    \I__1637\ : Span12Mux_h
    port map (
            O => \N__7935\,
            I => \N__7932\
        );

    \I__1636\ : Odrv12
    port map (
            O => \N__7932\,
            I => \A_c_9\
        );

    \I__1635\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7926\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__7926\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1633\ : InMux
    port map (
            O => \N__7923\,
            I => \N__7920\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__7920\,
            I => \N__7917\
        );

    \I__1631\ : Span4Mux_h
    port map (
            O => \N__7917\,
            I => \N__7914\
        );

    \I__1630\ : Span4Mux_v
    port map (
            O => \N__7914\,
            I => \N__7911\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__7911\,
            I => \U712_CHIP_RAM.un3_DMA_CYCLE_START\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7905\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__7905\,
            I => \U712_CYCLE_TERM.N_252_i_0_en\
        );

    \I__1626\ : CEMux
    port map (
            O => \N__7902\,
            I => \N__7899\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__7899\,
            I => \N__7896\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__7896\,
            I => \U712_CYCLE_TERM.N_252_i_0_en_0\
        );

    \I__1623\ : InMux
    port map (
            O => \N__7893\,
            I => \N__7890\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__7890\,
            I => \N__7887\
        );

    \I__1621\ : Odrv12
    port map (
            O => \N__7887\,
            I => \U712_BYTE_ENABLE.N_257\
        );

    \I__1620\ : InMux
    port map (
            O => \N__7884\,
            I => \N__7881\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7881\,
            I => \N__7878\
        );

    \I__1618\ : Odrv12
    port map (
            O => \N__7878\,
            I => \U712_BYTE_ENABLE.N_258\
        );

    \I__1617\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7872\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__7872\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__1615\ : IoInMux
    port map (
            O => \N__7869\,
            I => \N__7866\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__7866\,
            I => \N__7863\
        );

    \I__1613\ : Span12Mux_s2_v
    port map (
            O => \N__7863\,
            I => \N__7860\
        );

    \I__1612\ : Odrv12
    port map (
            O => \N__7860\,
            I => \CMA_c_1\
        );

    \I__1611\ : IoInMux
    port map (
            O => \N__7857\,
            I => \N__7854\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__7854\,
            I => \N__7851\
        );

    \I__1609\ : Span4Mux_s3_h
    port map (
            O => \N__7851\,
            I => \N__7848\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__7848\,
            I => \N__7845\
        );

    \I__1607\ : Span4Mux_v
    port map (
            O => \N__7845\,
            I => \N__7842\
        );

    \I__1606\ : Span4Mux_h
    port map (
            O => \N__7842\,
            I => \N__7839\
        );

    \I__1605\ : Sp12to4
    port map (
            O => \N__7839\,
            I => \N__7836\
        );

    \I__1604\ : Odrv12
    port map (
            O => \N__7836\,
            I => \CMA_c_3\
        );

    \I__1603\ : InMux
    port map (
            O => \N__7833\,
            I => \N__7830\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__7830\,
            I => \N__7825\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7829\,
            I => \N__7822\
        );

    \I__1600\ : IoInMux
    port map (
            O => \N__7828\,
            I => \N__7819\
        );

    \I__1599\ : Span4Mux_v
    port map (
            O => \N__7825\,
            I => \N__7816\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__7822\,
            I => \N__7813\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__7819\,
            I => \N__7810\
        );

    \I__1596\ : Span4Mux_h
    port map (
            O => \N__7816\,
            I => \N__7805\
        );

    \I__1595\ : Span4Mux_v
    port map (
            O => \N__7813\,
            I => \N__7805\
        );

    \I__1594\ : Span12Mux_s3_h
    port map (
            O => \N__7810\,
            I => \N__7802\
        );

    \I__1593\ : Span4Mux_v
    port map (
            O => \N__7805\,
            I => \N__7799\
        );

    \I__1592\ : Span12Mux_v
    port map (
            O => \N__7802\,
            I => \N__7796\
        );

    \I__1591\ : Span4Mux_v
    port map (
            O => \N__7799\,
            I => \N__7793\
        );

    \I__1590\ : Span12Mux_h
    port map (
            O => \N__7796\,
            I => \N__7790\
        );

    \I__1589\ : IoSpan4Mux
    port map (
            O => \N__7793\,
            I => \N__7787\
        );

    \I__1588\ : Odrv12
    port map (
            O => \N__7790\,
            I => \CLK40_PLL\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__7787\,
            I => \CLK40_PLL\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7782\,
            I => \N__7779\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7779\,
            I => \U712_CHIP_RAM.N_311\
        );

    \I__1584\ : InMux
    port map (
            O => \N__7776\,
            I => \N__7772\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7769\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7772\,
            I => \U712_CHIP_RAM.SDRAM_CMDs_1_3\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__7769\,
            I => \U712_CHIP_RAM.SDRAM_CMDs_1_3\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__7764\,
            I => \N__7761\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7758\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__7758\,
            I => \N__7754\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7751\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__7754\,
            I => \U712_CHIP_RAM.SDRAM_CMDs_0_6\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7751\,
            I => \U712_CHIP_RAM.SDRAM_CMDs_0_6\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7743\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7743\,
            I => \N__7738\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7742\,
            I => \N__7735\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7732\
        );

    \I__1570\ : Odrv4
    port map (
            O => \N__7738\,
            I => \U712_CHIP_RAM.N_377\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7735\,
            I => \U712_CHIP_RAM.N_377\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7732\,
            I => \U712_CHIP_RAM.N_377\
        );

    \I__1567\ : CEMux
    port map (
            O => \N__7725\,
            I => \N__7722\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7722\,
            I => \N__7719\
        );

    \I__1565\ : Span4Mux_v
    port map (
            O => \N__7719\,
            I => \N__7716\
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__7716\,
            I => \U712_CHIP_RAM.N_50_0\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7713\,
            I => \N__7709\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7712\,
            I => \N__7705\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7709\,
            I => \N__7702\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7708\,
            I => \N__7699\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7705\,
            I => \N__7696\
        );

    \I__1558\ : Span4Mux_v
    port map (
            O => \N__7702\,
            I => \N__7691\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7699\,
            I => \N__7691\
        );

    \I__1556\ : Span4Mux_h
    port map (
            O => \N__7696\,
            I => \N__7688\
        );

    \I__1555\ : Odrv4
    port map (
            O => \N__7691\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__7688\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1553\ : CascadeMux
    port map (
            O => \N__7683\,
            I => \N__7680\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7680\,
            I => \N__7677\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7677\,
            I => \N__7673\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7676\,
            I => \N__7670\
        );

    \I__1549\ : Odrv12
    port map (
            O => \N__7673\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7670\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__7665\,
            I => \U712_CYCLE_TERM.N_252_i_0_0_cascade_\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__7662\,
            I => \N__7658\
        );

    \I__1545\ : CascadeMux
    port map (
            O => \N__7661\,
            I => \N__7655\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7658\,
            I => \N__7651\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7655\,
            I => \N__7646\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7654\,
            I => \N__7643\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__7651\,
            I => \N__7640\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7650\,
            I => \N__7637\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7649\,
            I => \N__7634\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7646\,
            I => \N__7631\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__7643\,
            I => \N__7628\
        );

    \I__1536\ : Odrv4
    port map (
            O => \N__7640\,
            I => \REG_TACK\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__7637\,
            I => \REG_TACK\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7634\,
            I => \REG_TACK\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__7631\,
            I => \REG_TACK\
        );

    \I__1532\ : Odrv4
    port map (
            O => \N__7628\,
            I => \REG_TACK\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7617\,
            I => \N__7613\
        );

    \I__1530\ : InMux
    port map (
            O => \N__7616\,
            I => \N__7610\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__7613\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7610\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7605\,
            I => \N__7598\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7604\,
            I => \N__7595\
        );

    \I__1525\ : InMux
    port map (
            O => \N__7603\,
            I => \N__7590\
        );

    \I__1524\ : InMux
    port map (
            O => \N__7602\,
            I => \N__7590\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7601\,
            I => \N__7587\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7598\,
            I => \N__7584\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7595\,
            I => \N__7579\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7590\,
            I => \N__7579\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7587\,
            I => \CPU_TACK\
        );

    \I__1518\ : Odrv12
    port map (
            O => \N__7584\,
            I => \CPU_TACK\
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__7579\,
            I => \CPU_TACK\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__7572\,
            I => \N__7567\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__7571\,
            I => \N__7561\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7556\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7567\,
            I => \N__7556\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__7566\,
            I => \N__7553\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7550\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7564\,
            I => \N__7545\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7561\,
            I => \N__7545\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7556\,
            I => \N__7542\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7553\,
            I => \N__7539\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7550\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7545\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1504\ : Odrv4
    port map (
            O => \N__7542\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7539\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7530\,
            I => \N__7527\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7527\,
            I => \N__7522\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7526\,
            I => \N__7519\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7525\,
            I => \N__7516\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__7522\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7519\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__7516\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7509\,
            I => \N__7506\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7506\,
            I => \N__7503\
        );

    \I__1493\ : Span4Mux_h
    port map (
            O => \N__7503\,
            I => \N__7500\
        );

    \I__1492\ : Odrv4
    port map (
            O => \N__7500\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0\
        );

    \I__1491\ : IoInMux
    port map (
            O => \N__7497\,
            I => \N__7494\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__7494\,
            I => \N__7491\
        );

    \I__1489\ : IoSpan4Mux
    port map (
            O => \N__7491\,
            I => \N__7488\
        );

    \I__1488\ : Span4Mux_s3_h
    port map (
            O => \N__7488\,
            I => \N__7485\
        );

    \I__1487\ : Sp12to4
    port map (
            O => \N__7485\,
            I => \N__7482\
        );

    \I__1486\ : Span12Mux_h
    port map (
            O => \N__7482\,
            I => \N__7479\
        );

    \I__1485\ : Odrv12
    port map (
            O => \N__7479\,
            I => \N_205_i\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7476\,
            I => \N__7473\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7473\,
            I => \N__7470\
        );

    \I__1482\ : Span4Mux_v
    port map (
            O => \N__7470\,
            I => \N__7467\
        );

    \I__1481\ : Sp12to4
    port map (
            O => \N__7467\,
            I => \N__7464\
        );

    \I__1480\ : Span12Mux_h
    port map (
            O => \N__7464\,
            I => \N__7461\
        );

    \I__1479\ : Span12Mux_v
    port map (
            O => \N__7461\,
            I => \N__7458\
        );

    \I__1478\ : Odrv12
    port map (
            O => \N__7458\,
            I => \A_c_3\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7455\,
            I => \N__7452\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7452\,
            I => \N__7449\
        );

    \I__1475\ : Span12Mux_h
    port map (
            O => \N__7449\,
            I => \N__7446\
        );

    \I__1474\ : Odrv12
    port map (
            O => \N__7446\,
            I => \A_c_10\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7443\,
            I => \N__7440\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__7440\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7437\,
            I => \N__7432\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7436\,
            I => \N__7429\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7435\,
            I => \N__7426\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7432\,
            I => \U712_CHIP_RAM.N_248\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__7429\,
            I => \U712_CHIP_RAM.N_248\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7426\,
            I => \U712_CHIP_RAM.N_248\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7415\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7418\,
            I => \N__7412\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7415\,
            I => \N__7409\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7412\,
            I => \U712_CHIP_RAM.N_278\
        );

    \I__1461\ : Odrv4
    port map (
            O => \N__7409\,
            I => \U712_CHIP_RAM.N_278\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7404\,
            I => \N__7401\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7401\,
            I => \N__7398\
        );

    \I__1458\ : Span4Mux_h
    port map (
            O => \N__7398\,
            I => \N__7395\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__7395\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_0_0_3\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__7392\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_0_0_2_cascade_\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7389\,
            I => \N__7381\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7388\,
            I => \N__7375\
        );

    \I__1453\ : InMux
    port map (
            O => \N__7387\,
            I => \N__7375\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7370\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7370\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7384\,
            I => \N__7367\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7381\,
            I => \N__7360\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7380\,
            I => \N__7357\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7375\,
            I => \N__7354\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7370\,
            I => \N__7349\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7367\,
            I => \N__7349\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7366\,
            I => \N__7346\
        );

    \I__1443\ : InMux
    port map (
            O => \N__7365\,
            I => \N__7339\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7364\,
            I => \N__7339\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7363\,
            I => \N__7339\
        );

    \I__1440\ : Span4Mux_v
    port map (
            O => \N__7360\,
            I => \N__7336\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__7357\,
            I => \U712_CHIP_RAM.N_228\
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__7354\,
            I => \U712_CHIP_RAM.N_228\
        );

    \I__1437\ : Odrv4
    port map (
            O => \N__7349\,
            I => \U712_CHIP_RAM.N_228\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7346\,
            I => \U712_CHIP_RAM.N_228\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__7339\,
            I => \U712_CHIP_RAM.N_228\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__7336\,
            I => \U712_CHIP_RAM.N_228\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7323\,
            I => \N__7320\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7320\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_0_2\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__7317\,
            I => \U712_CHIP_RAM.N_50_cascade_\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7314\,
            I => \N__7311\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7311\,
            I => \N__7306\
        );

    \I__1428\ : InMux
    port map (
            O => \N__7310\,
            I => \N__7303\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7309\,
            I => \N__7300\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__7306\,
            I => \U712_CHIP_RAM.N_50\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7303\,
            I => \U712_CHIP_RAM.N_50\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__7300\,
            I => \U712_CHIP_RAM.N_50\
        );

    \I__1423\ : InMux
    port map (
            O => \N__7293\,
            I => \N__7286\
        );

    \I__1422\ : InMux
    port map (
            O => \N__7292\,
            I => \N__7283\
        );

    \I__1421\ : InMux
    port map (
            O => \N__7291\,
            I => \N__7278\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7290\,
            I => \N__7273\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7289\,
            I => \N__7273\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__7286\,
            I => \N__7264\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__7283\,
            I => \N__7261\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7282\,
            I => \N__7256\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7281\,
            I => \N__7256\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__7278\,
            I => \N__7250\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__7273\,
            I => \N__7242\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7272\,
            I => \N__7235\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7235\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7270\,
            I => \N__7235\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7269\,
            I => \N__7232\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7268\,
            I => \N__7227\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7267\,
            I => \N__7227\
        );

    \I__1406\ : Span4Mux_v
    port map (
            O => \N__7264\,
            I => \N__7224\
        );

    \I__1405\ : Span4Mux_v
    port map (
            O => \N__7261\,
            I => \N__7219\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7256\,
            I => \N__7219\
        );

    \I__1403\ : InMux
    port map (
            O => \N__7255\,
            I => \N__7212\
        );

    \I__1402\ : InMux
    port map (
            O => \N__7254\,
            I => \N__7212\
        );

    \I__1401\ : InMux
    port map (
            O => \N__7253\,
            I => \N__7212\
        );

    \I__1400\ : Span4Mux_h
    port map (
            O => \N__7250\,
            I => \N__7209\
        );

    \I__1399\ : InMux
    port map (
            O => \N__7249\,
            I => \N__7200\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7248\,
            I => \N__7200\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7247\,
            I => \N__7200\
        );

    \I__1396\ : InMux
    port map (
            O => \N__7246\,
            I => \N__7200\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7245\,
            I => \N__7197\
        );

    \I__1394\ : Span4Mux_h
    port map (
            O => \N__7242\,
            I => \N__7192\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7235\,
            I => \N__7192\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7232\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7227\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__7224\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1389\ : Odrv4
    port map (
            O => \N__7219\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__7212\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__7209\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7200\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7197\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1384\ : Odrv4
    port map (
            O => \N__7192\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__7173\,
            I => \N__7168\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__7172\,
            I => \N__7161\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__7171\,
            I => \N__7157\
        );

    \I__1380\ : InMux
    port map (
            O => \N__7168\,
            I => \N__7154\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7150\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__7166\,
            I => \N__7145\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__7165\,
            I => \N__7142\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7164\,
            I => \N__7135\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7161\,
            I => \N__7135\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7160\,
            I => \N__7132\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7157\,
            I => \N__7129\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7154\,
            I => \N__7126\
        );

    \I__1371\ : InMux
    port map (
            O => \N__7153\,
            I => \N__7123\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__7150\,
            I => \N__7120\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7149\,
            I => \N__7115\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7148\,
            I => \N__7115\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7110\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7142\,
            I => \N__7110\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7141\,
            I => \N__7103\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7103\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__7135\,
            I => \N__7100\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__7132\,
            I => \N__7097\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__7129\,
            I => \N__7092\
        );

    \I__1360\ : Span4Mux_h
    port map (
            O => \N__7126\,
            I => \N__7089\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7123\,
            I => \N__7086\
        );

    \I__1358\ : Span4Mux_h
    port map (
            O => \N__7120\,
            I => \N__7081\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7115\,
            I => \N__7081\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7110\,
            I => \N__7078\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7109\,
            I => \N__7073\
        );

    \I__1354\ : InMux
    port map (
            O => \N__7108\,
            I => \N__7073\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__7103\,
            I => \N__7066\
        );

    \I__1352\ : Span4Mux_h
    port map (
            O => \N__7100\,
            I => \N__7066\
        );

    \I__1351\ : Span4Mux_h
    port map (
            O => \N__7097\,
            I => \N__7066\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7096\,
            I => \N__7061\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7095\,
            I => \N__7061\
        );

    \I__1348\ : Odrv4
    port map (
            O => \N__7092\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__7089\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1346\ : Odrv4
    port map (
            O => \N__7086\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1345\ : Odrv4
    port map (
            O => \N__7081\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1344\ : Odrv12
    port map (
            O => \N__7078\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__7073\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1342\ : Odrv4
    port map (
            O => \N__7066\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__7061\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__7044\,
            I => \N__7039\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7043\,
            I => \N__7034\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7042\,
            I => \N__7034\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7039\,
            I => \N__7031\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7034\,
            I => \N__7023\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7031\,
            I => \N__7023\
        );

    \I__1334\ : InMux
    port map (
            O => \N__7030\,
            I => \N__7014\
        );

    \I__1333\ : InMux
    port map (
            O => \N__7029\,
            I => \N__7011\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7028\,
            I => \N__7008\
        );

    \I__1331\ : Span4Mux_h
    port map (
            O => \N__7023\,
            I => \N__7005\
        );

    \I__1330\ : InMux
    port map (
            O => \N__7022\,
            I => \N__7002\
        );

    \I__1329\ : InMux
    port map (
            O => \N__7021\,
            I => \N__6997\
        );

    \I__1328\ : InMux
    port map (
            O => \N__7020\,
            I => \N__6997\
        );

    \I__1327\ : InMux
    port map (
            O => \N__7019\,
            I => \N__6992\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7018\,
            I => \N__6992\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7017\,
            I => \N__6989\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__7014\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__7011\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__7008\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__7005\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__7002\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6997\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__6992\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6989\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6972\,
            I => \N__6969\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__6969\,
            I => \N__6965\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6968\,
            I => \N__6962\
        );

    \I__1313\ : Span4Mux_h
    port map (
            O => \N__6965\,
            I => \N__6959\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6962\,
            I => \U712_CHIP_RAM.N_263\
        );

    \I__1311\ : Odrv4
    port map (
            O => \N__6959\,
            I => \U712_CHIP_RAM.N_263\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__6954\,
            I => \U712_CHIP_RAM.N_280_cascade_\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6951\,
            I => \N__6948\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__6948\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_0_3\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__6945\,
            I => \N__6941\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__6944\,
            I => \N__6929\
        );

    \I__1305\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6925\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6921\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__6939\,
            I => \N__6916\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6938\,
            I => \N__6913\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6910\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6936\,
            I => \N__6907\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6935\,
            I => \N__6902\
        );

    \I__1298\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6902\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6933\,
            I => \N__6893\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6893\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6929\,
            I => \N__6893\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6928\,
            I => \N__6893\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6925\,
            I => \N__6888\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6924\,
            I => \N__6885\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__6921\,
            I => \N__6882\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6920\,
            I => \N__6875\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6919\,
            I => \N__6875\
        );

    \I__1288\ : InMux
    port map (
            O => \N__6916\,
            I => \N__6875\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__6913\,
            I => \N__6870\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__6910\,
            I => \N__6870\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__6907\,
            I => \N__6863\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__6902\,
            I => \N__6863\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6893\,
            I => \N__6863\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6892\,
            I => \N__6860\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6891\,
            I => \N__6857\
        );

    \I__1280\ : Span4Mux_v
    port map (
            O => \N__6888\,
            I => \N__6852\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6885\,
            I => \N__6852\
        );

    \I__1278\ : Span4Mux_h
    port map (
            O => \N__6882\,
            I => \N__6849\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6875\,
            I => \N__6846\
        );

    \I__1276\ : Span4Mux_h
    port map (
            O => \N__6870\,
            I => \N__6843\
        );

    \I__1275\ : Span4Mux_h
    port map (
            O => \N__6863\,
            I => \N__6840\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__6860\,
            I => \N__6837\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__6857\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__6852\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__6849\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__6846\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__6843\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1268\ : Odrv4
    port map (
            O => \N__6840\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1267\ : Odrv12
    port map (
            O => \N__6837\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6822\,
            I => \N__6819\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6819\,
            I => \N__6816\
        );

    \I__1264\ : Odrv4
    port map (
            O => \N__6816\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6813\,
            I => \N__6810\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__6810\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_0\
        );

    \I__1261\ : InMux
    port map (
            O => \N__6807\,
            I => \N__6804\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6804\,
            I => \N__6801\
        );

    \I__1259\ : Span4Mux_v
    port map (
            O => \N__6801\,
            I => \N__6798\
        );

    \I__1258\ : Odrv4
    port map (
            O => \N__6798\,
            I => \U712_CHIP_RAM.N_130\
        );

    \I__1257\ : IoInMux
    port map (
            O => \N__6795\,
            I => \N__6792\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__6792\,
            I => \N__6789\
        );

    \I__1255\ : Span4Mux_s2_h
    port map (
            O => \N__6789\,
            I => \N__6786\
        );

    \I__1254\ : Span4Mux_h
    port map (
            O => \N__6786\,
            I => \N__6783\
        );

    \I__1253\ : Sp12to4
    port map (
            O => \N__6783\,
            I => \N__6780\
        );

    \I__1252\ : Span12Mux_s11_v
    port map (
            O => \N__6780\,
            I => \N__6777\
        );

    \I__1251\ : Span12Mux_h
    port map (
            O => \N__6777\,
            I => \N__6773\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6770\
        );

    \I__1249\ : Odrv12
    port map (
            O => \N__6773\,
            I => \CLK_EN_c\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6770\,
            I => \CLK_EN_c\
        );

    \I__1247\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6762\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6762\,
            I => \N__6759\
        );

    \I__1245\ : Span4Mux_v
    port map (
            O => \N__6759\,
            I => \N__6756\
        );

    \I__1244\ : Span4Mux_h
    port map (
            O => \N__6756\,
            I => \N__6753\
        );

    \I__1243\ : Span4Mux_v
    port map (
            O => \N__6753\,
            I => \N__6750\
        );

    \I__1242\ : Odrv4
    port map (
            O => \N__6750\,
            I => \TACK_EN_i_ess\
        );

    \I__1241\ : IoInMux
    port map (
            O => \N__6747\,
            I => \N__6744\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__6744\,
            I => \N__6741\
        );

    \I__1239\ : Span4Mux_s1_v
    port map (
            O => \N__6741\,
            I => \N__6737\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6740\,
            I => \N__6734\
        );

    \I__1237\ : Span4Mux_v
    port map (
            O => \N__6737\,
            I => \N__6731\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6734\,
            I => \N__6728\
        );

    \I__1235\ : Span4Mux_h
    port map (
            O => \N__6731\,
            I => \N__6725\
        );

    \I__1234\ : Span4Mux_v
    port map (
            O => \N__6728\,
            I => \N__6722\
        );

    \I__1233\ : Odrv4
    port map (
            O => \N__6725\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1232\ : Odrv4
    port map (
            O => \N__6722\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6717\,
            I => \N__6714\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__6714\,
            I => \N__6711\
        );

    \I__1229\ : Span4Mux_v
    port map (
            O => \N__6711\,
            I => \N__6708\
        );

    \I__1228\ : Span4Mux_v
    port map (
            O => \N__6708\,
            I => \N__6705\
        );

    \I__1227\ : Sp12to4
    port map (
            O => \N__6705\,
            I => \N__6702\
        );

    \I__1226\ : Span12Mux_h
    port map (
            O => \N__6702\,
            I => \N__6699\
        );

    \I__1225\ : Odrv12
    port map (
            O => \N__6699\,
            I => \A_c_7\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__6696\,
            I => \U712_CHIP_RAM.N_292_cascade_\
        );

    \I__1223\ : IoInMux
    port map (
            O => \N__6693\,
            I => \N__6690\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__6690\,
            I => \N__6687\
        );

    \I__1221\ : Span12Mux_s10_v
    port map (
            O => \N__6687\,
            I => \N__6684\
        );

    \I__1220\ : Odrv12
    port map (
            O => \N__6684\,
            I => \N_207_i\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6681\,
            I => \N__6678\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6678\,
            I => \N__6675\
        );

    \I__1217\ : Span4Mux_v
    port map (
            O => \N__6675\,
            I => \N__6672\
        );

    \I__1216\ : Sp12to4
    port map (
            O => \N__6672\,
            I => \N__6669\
        );

    \I__1215\ : Span12Mux_h
    port map (
            O => \N__6669\,
            I => \N__6666\
        );

    \I__1214\ : Odrv12
    port map (
            O => \N__6666\,
            I => \A_c_13\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6663\,
            I => \N__6660\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6660\,
            I => \N__6657\
        );

    \I__1211\ : Span4Mux_v
    port map (
            O => \N__6657\,
            I => \N__6654\
        );

    \I__1210\ : Span4Mux_v
    port map (
            O => \N__6654\,
            I => \N__6651\
        );

    \I__1209\ : Span4Mux_h
    port map (
            O => \N__6651\,
            I => \N__6648\
        );

    \I__1208\ : Sp12to4
    port map (
            O => \N__6648\,
            I => \N__6645\
        );

    \I__1207\ : Odrv12
    port map (
            O => \N__6645\,
            I => \A_c_6\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__6642\,
            I => \U712_CHIP_RAM.SDRAM_CMDs_0_6_cascade_\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__6639\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6631\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6621\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__6634\,
            I => \N__6618\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6631\,
            I => \N__6614\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6630\,
            I => \N__6607\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6604\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6628\,
            I => \N__6601\
        );

    \I__1197\ : InMux
    port map (
            O => \N__6627\,
            I => \N__6598\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6626\,
            I => \N__6593\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6625\,
            I => \N__6593\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6624\,
            I => \N__6590\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6621\,
            I => \N__6587\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6618\,
            I => \N__6584\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6617\,
            I => \N__6581\
        );

    \I__1190\ : Span4Mux_h
    port map (
            O => \N__6614\,
            I => \N__6578\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6575\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6612\,
            I => \N__6568\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6611\,
            I => \N__6568\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6568\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6607\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6604\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6601\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6598\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6593\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6590\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__6587\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6584\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6581\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__6578\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6575\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6568\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6543\,
            I => \N__6539\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6542\,
            I => \N__6536\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6539\,
            I => \N__6533\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6536\,
            I => \N__6524\
        );

    \I__1169\ : Glb2LocalMux
    port map (
            O => \N__6533\,
            I => \N__6507\
        );

    \I__1168\ : ClkMux
    port map (
            O => \N__6532\,
            I => \N__6507\
        );

    \I__1167\ : ClkMux
    port map (
            O => \N__6531\,
            I => \N__6507\
        );

    \I__1166\ : ClkMux
    port map (
            O => \N__6530\,
            I => \N__6507\
        );

    \I__1165\ : ClkMux
    port map (
            O => \N__6529\,
            I => \N__6507\
        );

    \I__1164\ : ClkMux
    port map (
            O => \N__6528\,
            I => \N__6507\
        );

    \I__1163\ : ClkMux
    port map (
            O => \N__6527\,
            I => \N__6507\
        );

    \I__1162\ : Glb2LocalMux
    port map (
            O => \N__6524\,
            I => \N__6507\
        );

    \I__1161\ : GlobalMux
    port map (
            O => \N__6507\,
            I => \N__6504\
        );

    \I__1160\ : gio2CtrlBuf
    port map (
            O => \N__6504\,
            I => \CLK40_PLL_g\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__6501\,
            I => \U712_CYCLE_TERM.TACK_STATE_r_sx_1_cascade_\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6495\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6495\,
            I => \U712_CHIP_RAM.N_281\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__6492\,
            I => \N__6483\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__6491\,
            I => \N__6480\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6490\,
            I => \N__6473\
        );

    \I__1153\ : InMux
    port map (
            O => \N__6489\,
            I => \N__6473\
        );

    \I__1152\ : InMux
    port map (
            O => \N__6488\,
            I => \N__6473\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6463\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6460\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6483\,
            I => \N__6457\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6454\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6473\,
            I => \N__6451\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6472\,
            I => \N__6444\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6471\,
            I => \N__6444\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6470\,
            I => \N__6444\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6469\,
            I => \N__6439\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6439\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6467\,
            I => \N__6434\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6466\,
            I => \N__6434\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6463\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__6460\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6457\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6454\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1135\ : Odrv4
    port map (
            O => \N__6451\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6444\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6439\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6434\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6417\,
            I => \N__6414\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__6414\,
            I => \U712_CHIP_RAM.N_283\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6411\,
            I => \N__6408\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6408\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_4\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6405\,
            I => \N__6402\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6402\,
            I => \N__6399\
        );

    \I__1125\ : Odrv12
    port map (
            O => \N__6399\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_5\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6396\,
            I => \N__6393\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6393\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_0_0\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6387\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6387\,
            I => \N__6384\
        );

    \I__1120\ : Span4Mux_v
    port map (
            O => \N__6384\,
            I => \N__6381\
        );

    \I__1119\ : Odrv4
    port map (
            O => \N__6381\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_3\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__6378\,
            I => \U712_CHIP_RAM.CLK_EN_5_0_i_i_a2_0_a3_1_cascade_\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6375\,
            I => \N__6372\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6372\,
            I => \N__6368\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6365\
        );

    \I__1114\ : Span4Mux_v
    port map (
            O => \N__6368\,
            I => \N__6361\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__6365\,
            I => \N__6358\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6364\,
            I => \N__6355\
        );

    \I__1111\ : Odrv4
    port map (
            O => \N__6361\,
            I => \U712_CHIP_RAM.N_374\
        );

    \I__1110\ : Odrv4
    port map (
            O => \N__6358\,
            I => \U712_CHIP_RAM.N_374\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6355\,
            I => \U712_CHIP_RAM.N_374\
        );

    \I__1108\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6343\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__6347\,
            I => \N__6338\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__6346\,
            I => \N__6335\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6343\,
            I => \N__6331\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6342\,
            I => \N__6326\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6341\,
            I => \N__6323\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6338\,
            I => \N__6316\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6316\
        );

    \I__1100\ : InMux
    port map (
            O => \N__6334\,
            I => \N__6316\
        );

    \I__1099\ : Span4Mux_v
    port map (
            O => \N__6331\,
            I => \N__6311\
        );

    \I__1098\ : InMux
    port map (
            O => \N__6330\,
            I => \N__6306\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6329\,
            I => \N__6306\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__6326\,
            I => \N__6299\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__6323\,
            I => \N__6299\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6316\,
            I => \N__6299\
        );

    \I__1093\ : InMux
    port map (
            O => \N__6315\,
            I => \N__6294\
        );

    \I__1092\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6294\
        );

    \I__1091\ : Odrv4
    port map (
            O => \N__6311\,
            I => \WRITE_CYCLE\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__6306\,
            I => \WRITE_CYCLE\
        );

    \I__1089\ : Odrv4
    port map (
            O => \N__6299\,
            I => \WRITE_CYCLE\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__6294\,
            I => \WRITE_CYCLE\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__6285\,
            I => \U712_CHIP_RAM.N_130_cascade_\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6282\,
            I => \N__6279\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6279\,
            I => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__6276\,
            I => \U712_CHIP_RAM.N_60_cascade_\
        );

    \I__1083\ : InMux
    port map (
            O => \N__6273\,
            I => \N__6270\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__6270\,
            I => \U712_CHIP_RAM.SDRAM_CMDsr_0_1\
        );

    \I__1081\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6263\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6266\,
            I => \N__6257\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6263\,
            I => \N__6254\
        );

    \I__1078\ : InMux
    port map (
            O => \N__6262\,
            I => \N__6251\
        );

    \I__1077\ : InMux
    port map (
            O => \N__6261\,
            I => \N__6246\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6246\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6257\,
            I => \U712_CHIP_RAM.N_57\
        );

    \I__1074\ : Odrv4
    port map (
            O => \N__6254\,
            I => \U712_CHIP_RAM.N_57\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__6251\,
            I => \U712_CHIP_RAM.N_57\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__6246\,
            I => \U712_CHIP_RAM.N_57\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6237\,
            I => \N__6234\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__6234\,
            I => \N__6230\
        );

    \I__1069\ : InMux
    port map (
            O => \N__6233\,
            I => \N__6226\
        );

    \I__1068\ : Span4Mux_v
    port map (
            O => \N__6230\,
            I => \N__6223\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6229\,
            I => \N__6220\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6226\,
            I => \N__6213\
        );

    \I__1065\ : Sp12to4
    port map (
            O => \N__6223\,
            I => \N__6213\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__6220\,
            I => \N__6213\
        );

    \I__1063\ : Span12Mux_h
    port map (
            O => \N__6213\,
            I => \N__6210\
        );

    \I__1062\ : Span12Mux_v
    port map (
            O => \N__6210\,
            I => \N__6207\
        );

    \I__1061\ : Odrv12
    port map (
            O => \N__6207\,
            I => \RnW_c\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__6204\,
            I => \N__6200\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__6203\,
            I => \N__6194\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6200\,
            I => \N__6191\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6186\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6186\
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__6197\,
            I => \N__6181\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6178\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__6191\,
            I => \N__6174\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6186\,
            I => \N__6171\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6168\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6163\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6163\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__6178\,
            I => \N__6160\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6177\,
            I => \N__6157\
        );

    \I__1046\ : Span4Mux_h
    port map (
            O => \N__6174\,
            I => \N__6152\
        );

    \I__1045\ : Span4Mux_v
    port map (
            O => \N__6171\,
            I => \N__6152\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__6168\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6163\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1042\ : Odrv4
    port map (
            O => \N__6160\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__6157\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1040\ : Odrv4
    port map (
            O => \N__6152\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6141\,
            I => \N__6135\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6132\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6139\,
            I => \N__6127\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6138\,
            I => \N__6127\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6135\,
            I => \U712_REG_SM.N_255\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6132\,
            I => \U712_REG_SM.N_255\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6127\,
            I => \U712_REG_SM.N_255\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6120\,
            I => \N__6115\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6119\,
            I => \N__6112\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6118\,
            I => \N__6109\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6115\,
            I => \N__6106\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__6112\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_6\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__6109\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_6\
        );

    \I__1026\ : Odrv12
    port map (
            O => \N__6106\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_6\
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__6099\,
            I => \N__6094\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6098\,
            I => \N__6089\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6082\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6079\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6074\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6074\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6089\,
            I => \N__6071\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6062\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6087\,
            I => \N__6062\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6086\,
            I => \N__6062\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6062\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__6082\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__6079\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6074\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1011\ : Odrv4
    port map (
            O => \N__6071\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__6062\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6048\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6048\,
            I => \U712_REG_SM.N_274\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6045\,
            I => \N__6040\
        );

    \I__1006\ : InMux
    port map (
            O => \N__6044\,
            I => \N__6037\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6043\,
            I => \N__6034\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6040\,
            I => \N__6029\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6037\,
            I => \N__6026\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6034\,
            I => \N__6023\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6033\,
            I => \N__6018\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6032\,
            I => \N__6018\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__6029\,
            I => \REG_WRITE_CYCLE\
        );

    \I__998\ : Odrv4
    port map (
            O => \N__6026\,
            I => \REG_WRITE_CYCLE\
        );

    \I__997\ : Odrv12
    port map (
            O => \N__6023\,
            I => \REG_WRITE_CYCLE\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__6018\,
            I => \REG_WRITE_CYCLE\
        );

    \I__995\ : InMux
    port map (
            O => \N__6009\,
            I => \N__6004\
        );

    \I__994\ : InMux
    port map (
            O => \N__6008\,
            I => \N__6001\
        );

    \I__993\ : InMux
    port map (
            O => \N__6007\,
            I => \N__5998\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__6004\,
            I => \U712_REG_SM.STATE_COUNTERc_1\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__6001\,
            I => \U712_REG_SM.STATE_COUNTERc_1\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__5998\,
            I => \U712_REG_SM.STATE_COUNTERc_1\
        );

    \I__989\ : CascadeMux
    port map (
            O => \N__5991\,
            I => \N__5988\
        );

    \I__988\ : InMux
    port map (
            O => \N__5988\,
            I => \N__5983\
        );

    \I__987\ : InMux
    port map (
            O => \N__5987\,
            I => \N__5980\
        );

    \I__986\ : InMux
    port map (
            O => \N__5986\,
            I => \N__5977\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__5983\,
            I => \N__5974\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5980\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_4\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5977\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_4\
        );

    \I__982\ : Odrv4
    port map (
            O => \N__5974\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_4\
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__5967\,
            I => \N__5963\
        );

    \I__980\ : InMux
    port map (
            O => \N__5966\,
            I => \N__5958\
        );

    \I__979\ : InMux
    port map (
            O => \N__5963\,
            I => \N__5958\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5958\,
            I => \N__5951\
        );

    \I__977\ : InMux
    port map (
            O => \N__5957\,
            I => \N__5944\
        );

    \I__976\ : InMux
    port map (
            O => \N__5956\,
            I => \N__5944\
        );

    \I__975\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5944\
        );

    \I__974\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5941\
        );

    \I__973\ : Odrv4
    port map (
            O => \N__5951\,
            I => \U712_REG_SM.LATCH_REG_0_sqmuxa\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5944\,
            I => \U712_REG_SM.LATCH_REG_0_sqmuxa\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__5941\,
            I => \U712_REG_SM.LATCH_REG_0_sqmuxa\
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__5934\,
            I => \N__5931\
        );

    \I__969\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5928\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5928\,
            I => \N__5925\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__5925\,
            I => \U712_REG_SM.REG_CPU_CYCLE_e_1\
        );

    \I__966\ : SRMux
    port map (
            O => \N__5922\,
            I => \N__5919\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__5919\,
            I => \N__5916\
        );

    \I__964\ : Odrv4
    port map (
            O => \N__5916\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__963\ : CascadeMux
    port map (
            O => \N__5913\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_0_2_cascade_\
        );

    \I__962\ : InMux
    port map (
            O => \N__5910\,
            I => \N__5907\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__5907\,
            I => \N__5903\
        );

    \I__960\ : InMux
    port map (
            O => \N__5906\,
            I => \N__5900\
        );

    \I__959\ : Span4Mux_v
    port map (
            O => \N__5903\,
            I => \N__5894\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__5900\,
            I => \N__5891\
        );

    \I__957\ : InMux
    port map (
            O => \N__5899\,
            I => \N__5886\
        );

    \I__956\ : InMux
    port map (
            O => \N__5898\,
            I => \N__5886\
        );

    \I__955\ : InMux
    port map (
            O => \N__5897\,
            I => \N__5883\
        );

    \I__954\ : Odrv4
    port map (
            O => \N__5894\,
            I => \U712_CHIP_RAM.N_239\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__5891\,
            I => \U712_CHIP_RAM.N_239\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__5886\,
            I => \U712_CHIP_RAM.N_239\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__5883\,
            I => \U712_CHIP_RAM.N_239\
        );

    \I__950\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5871\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5871\,
            I => \N__5868\
        );

    \I__948\ : Span12Mux_v
    port map (
            O => \N__5868\,
            I => \N__5865\
        );

    \I__947\ : Span12Mux_h
    port map (
            O => \N__5865\,
            I => \N__5862\
        );

    \I__946\ : Odrv12
    port map (
            O => \N__5862\,
            I => \A_c_16\
        );

    \I__945\ : InMux
    port map (
            O => \N__5859\,
            I => \N__5856\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5856\,
            I => \N__5853\
        );

    \I__943\ : Span12Mux_v
    port map (
            O => \N__5853\,
            I => \N__5850\
        );

    \I__942\ : Span12Mux_h
    port map (
            O => \N__5850\,
            I => \N__5847\
        );

    \I__941\ : Odrv12
    port map (
            O => \N__5847\,
            I => \A_c_18\
        );

    \I__940\ : InMux
    port map (
            O => \N__5844\,
            I => \N__5840\
        );

    \I__939\ : CascadeMux
    port map (
            O => \N__5843\,
            I => \N__5837\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5840\,
            I => \N__5834\
        );

    \I__937\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5830\
        );

    \I__936\ : Span4Mux_h
    port map (
            O => \N__5834\,
            I => \N__5827\
        );

    \I__935\ : InMux
    port map (
            O => \N__5833\,
            I => \N__5824\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5830\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_3\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__5827\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_3\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__5824\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_3\
        );

    \I__931\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5814\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__5814\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_5\
        );

    \I__929\ : InMux
    port map (
            O => \N__5811\,
            I => \N__5808\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5808\,
            I => \U712_REG_SM.N_339\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__5805\,
            I => \N__5802\
        );

    \I__926\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5799\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__5799\,
            I => \N__5796\
        );

    \I__924\ : Odrv4
    port map (
            O => \N__5796\,
            I => \U712_REG_SM.LDSn_7_iv_i_0\
        );

    \I__923\ : IoInMux
    port map (
            O => \N__5793\,
            I => \N__5790\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__5790\,
            I => \N__5787\
        );

    \I__921\ : Span4Mux_s1_v
    port map (
            O => \N__5787\,
            I => \N__5784\
        );

    \I__920\ : Span4Mux_v
    port map (
            O => \N__5784\,
            I => \N__5781\
        );

    \I__919\ : Sp12to4
    port map (
            O => \N__5781\,
            I => \N__5778\
        );

    \I__918\ : Span12Mux_s11_h
    port map (
            O => \N__5778\,
            I => \N__5775\
        );

    \I__917\ : Span12Mux_v
    port map (
            O => \N__5775\,
            I => \N__5769\
        );

    \I__916\ : InMux
    port map (
            O => \N__5774\,
            I => \N__5766\
        );

    \I__915\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5763\
        );

    \I__914\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5760\
        );

    \I__913\ : Odrv12
    port map (
            O => \N__5769\,
            I => \LDSn_c\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__5766\,
            I => \LDSn_c\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__5763\,
            I => \LDSn_c\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__5760\,
            I => \LDSn_c\
        );

    \I__909\ : InMux
    port map (
            O => \N__5751\,
            I => \N__5748\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__5748\,
            I => \U712_REG_SM.UDSn_7_iv_i_0\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__5745\,
            I => \N__5742\
        );

    \I__906\ : InMux
    port map (
            O => \N__5742\,
            I => \N__5739\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__5739\,
            I => \U712_REG_SM.N_337\
        );

    \I__904\ : InMux
    port map (
            O => \N__5736\,
            I => \N__5730\
        );

    \I__903\ : InMux
    port map (
            O => \N__5735\,
            I => \N__5730\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5730\,
            I => \U712_REG_SM.N_169\
        );

    \I__901\ : IoInMux
    port map (
            O => \N__5727\,
            I => \N__5724\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__5724\,
            I => \N__5721\
        );

    \I__899\ : Span4Mux_s0_v
    port map (
            O => \N__5721\,
            I => \N__5718\
        );

    \I__898\ : Span4Mux_v
    port map (
            O => \N__5718\,
            I => \N__5715\
        );

    \I__897\ : Span4Mux_v
    port map (
            O => \N__5715\,
            I => \N__5712\
        );

    \I__896\ : Sp12to4
    port map (
            O => \N__5712\,
            I => \N__5709\
        );

    \I__895\ : Span12Mux_h
    port map (
            O => \N__5709\,
            I => \N__5703\
        );

    \I__894\ : InMux
    port map (
            O => \N__5708\,
            I => \N__5700\
        );

    \I__893\ : InMux
    port map (
            O => \N__5707\,
            I => \N__5697\
        );

    \I__892\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5694\
        );

    \I__891\ : Odrv12
    port map (
            O => \N__5703\,
            I => \UDSn_c\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5700\,
            I => \UDSn_c\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__5697\,
            I => \UDSn_c\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5694\,
            I => \UDSn_c\
        );

    \I__887\ : InMux
    port map (
            O => \N__5685\,
            I => \N__5682\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5682\,
            I => \N__5679\
        );

    \I__885\ : Span4Mux_v
    port map (
            O => \N__5679\,
            I => \N__5675\
        );

    \I__884\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5672\
        );

    \I__883\ : Odrv4
    port map (
            O => \N__5675\,
            I => \REG_CPU_CYCLE\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__5672\,
            I => \REG_CPU_CYCLE\
        );

    \I__881\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5664\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5664\,
            I => \U712_REG_SM.un15_0_i_0_0\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__5661\,
            I => \N__5656\
        );

    \I__878\ : InMux
    port map (
            O => \N__5660\,
            I => \N__5653\
        );

    \I__877\ : InMux
    port map (
            O => \N__5659\,
            I => \N__5645\
        );

    \I__876\ : InMux
    port map (
            O => \N__5656\,
            I => \N__5642\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5653\,
            I => \N__5639\
        );

    \I__874\ : InMux
    port map (
            O => \N__5652\,
            I => \N__5632\
        );

    \I__873\ : InMux
    port map (
            O => \N__5651\,
            I => \N__5632\
        );

    \I__872\ : InMux
    port map (
            O => \N__5650\,
            I => \N__5632\
        );

    \I__871\ : InMux
    port map (
            O => \N__5649\,
            I => \N__5627\
        );

    \I__870\ : InMux
    port map (
            O => \N__5648\,
            I => \N__5627\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5645\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5642\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__867\ : Odrv4
    port map (
            O => \N__5639\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5632\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5627\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__864\ : InMux
    port map (
            O => \N__5616\,
            I => \N__5613\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5613\,
            I => \N__5606\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__5612\,
            I => \N__5601\
        );

    \I__861\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5598\
        );

    \I__860\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5595\
        );

    \I__859\ : InMux
    port map (
            O => \N__5609\,
            I => \N__5592\
        );

    \I__858\ : Span4Mux_v
    port map (
            O => \N__5606\,
            I => \N__5589\
        );

    \I__857\ : InMux
    port map (
            O => \N__5605\,
            I => \N__5582\
        );

    \I__856\ : InMux
    port map (
            O => \N__5604\,
            I => \N__5582\
        );

    \I__855\ : InMux
    port map (
            O => \N__5601\,
            I => \N__5582\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__5598\,
            I => \N__5577\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5595\,
            I => \N__5577\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5592\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__851\ : Odrv4
    port map (
            O => \N__5589\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5582\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__849\ : Odrv4
    port map (
            O => \N__5577\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__5568\,
            I => \N__5563\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__5567\,
            I => \N__5559\
        );

    \I__846\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5552\
        );

    \I__845\ : InMux
    port map (
            O => \N__5563\,
            I => \N__5552\
        );

    \I__844\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5549\
        );

    \I__843\ : InMux
    port map (
            O => \N__5559\,
            I => \N__5546\
        );

    \I__842\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5541\
        );

    \I__841\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5541\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5552\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5549\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5546\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5541\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__836\ : InMux
    port map (
            O => \N__5532\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__835\ : InMux
    port map (
            O => \N__5529\,
            I => \N__5525\
        );

    \I__834\ : InMux
    port map (
            O => \N__5528\,
            I => \N__5522\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__5525\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5522\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__831\ : InMux
    port map (
            O => \N__5517\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__830\ : InMux
    port map (
            O => \N__5514\,
            I => \N__5510\
        );

    \I__829\ : InMux
    port map (
            O => \N__5513\,
            I => \N__5507\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5510\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5507\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__826\ : InMux
    port map (
            O => \N__5502\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__825\ : InMux
    port map (
            O => \N__5499\,
            I => \N__5494\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__5498\,
            I => \N__5489\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__5497\,
            I => \N__5483\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5494\,
            I => \N__5480\
        );

    \I__821\ : InMux
    port map (
            O => \N__5493\,
            I => \N__5473\
        );

    \I__820\ : InMux
    port map (
            O => \N__5492\,
            I => \N__5473\
        );

    \I__819\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5473\
        );

    \I__818\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5464\
        );

    \I__817\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5464\
        );

    \I__816\ : InMux
    port map (
            O => \N__5486\,
            I => \N__5464\
        );

    \I__815\ : InMux
    port map (
            O => \N__5483\,
            I => \N__5464\
        );

    \I__814\ : Odrv12
    port map (
            O => \N__5480\,
            I => \U712_CHIP_RAM.N_58\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5473\,
            I => \U712_CHIP_RAM.N_58\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5464\,
            I => \U712_CHIP_RAM.N_58\
        );

    \I__811\ : InMux
    port map (
            O => \N__5457\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__810\ : InMux
    port map (
            O => \N__5454\,
            I => \N__5450\
        );

    \I__809\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5447\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5450\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__5447\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__806\ : CEMux
    port map (
            O => \N__5442\,
            I => \N__5439\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5439\,
            I => \N__5435\
        );

    \I__804\ : CEMux
    port map (
            O => \N__5438\,
            I => \N__5432\
        );

    \I__803\ : Span4Mux_h
    port map (
            O => \N__5435\,
            I => \N__5429\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5432\,
            I => \N__5426\
        );

    \I__801\ : Span4Mux_h
    port map (
            O => \N__5429\,
            I => \N__5423\
        );

    \I__800\ : Span4Mux_v
    port map (
            O => \N__5426\,
            I => \N__5420\
        );

    \I__799\ : Odrv4
    port map (
            O => \N__5423\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__798\ : Odrv4
    port map (
            O => \N__5420\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__797\ : InMux
    port map (
            O => \N__5415\,
            I => \N__5412\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5412\,
            I => \N__5409\
        );

    \I__795\ : Odrv12
    port map (
            O => \N__5409\,
            I => \U712_CHIP_RAM.N_378\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__5406\,
            I => \N__5403\
        );

    \I__793\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5395\
        );

    \I__792\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5395\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__5401\,
            I => \N__5390\
        );

    \I__790\ : InMux
    port map (
            O => \N__5400\,
            I => \N__5383\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5395\,
            I => \N__5380\
        );

    \I__788\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5377\
        );

    \I__787\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5370\
        );

    \I__786\ : InMux
    port map (
            O => \N__5390\,
            I => \N__5370\
        );

    \I__785\ : InMux
    port map (
            O => \N__5389\,
            I => \N__5370\
        );

    \I__784\ : InMux
    port map (
            O => \N__5388\,
            I => \N__5365\
        );

    \I__783\ : InMux
    port map (
            O => \N__5387\,
            I => \N__5365\
        );

    \I__782\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5362\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5383\,
            I => \U712_CHIP_RAM.N_367\
        );

    \I__780\ : Odrv4
    port map (
            O => \N__5380\,
            I => \U712_CHIP_RAM.N_367\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5377\,
            I => \U712_CHIP_RAM.N_367\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5370\,
            I => \U712_CHIP_RAM.N_367\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5365\,
            I => \U712_CHIP_RAM.N_367\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__5362\,
            I => \U712_CHIP_RAM.N_367\
        );

    \I__775\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5345\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__5348\,
            I => \N__5338\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__5345\,
            I => \N__5332\
        );

    \I__772\ : InMux
    port map (
            O => \N__5344\,
            I => \N__5328\
        );

    \I__771\ : InMux
    port map (
            O => \N__5343\,
            I => \N__5323\
        );

    \I__770\ : InMux
    port map (
            O => \N__5342\,
            I => \N__5323\
        );

    \I__769\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5320\
        );

    \I__768\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5315\
        );

    \I__767\ : InMux
    port map (
            O => \N__5337\,
            I => \N__5315\
        );

    \I__766\ : InMux
    port map (
            O => \N__5336\,
            I => \N__5312\
        );

    \I__765\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5309\
        );

    \I__764\ : Span4Mux_h
    port map (
            O => \N__5332\,
            I => \N__5306\
        );

    \I__763\ : InMux
    port map (
            O => \N__5331\,
            I => \N__5303\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__5328\,
            I => \N__5298\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__5323\,
            I => \N__5298\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__5320\,
            I => \N__5293\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5315\,
            I => \N__5293\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5312\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__5309\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__5306\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__5303\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__754\ : Odrv4
    port map (
            O => \N__5298\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__753\ : Odrv4
    port map (
            O => \N__5293\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__752\ : CEMux
    port map (
            O => \N__5280\,
            I => \N__5277\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__5277\,
            I => \N__5274\
        );

    \I__750\ : Span4Mux_h
    port map (
            O => \N__5274\,
            I => \N__5271\
        );

    \I__749\ : Odrv4
    port map (
            O => \N__5271\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__5268\,
            I => \U712_CHIP_RAM.N_237_cascade_\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__5265\,
            I => \N__5260\
        );

    \I__746\ : CascadeMux
    port map (
            O => \N__5264\,
            I => \N__5256\
        );

    \I__745\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5251\
        );

    \I__744\ : InMux
    port map (
            O => \N__5260\,
            I => \N__5251\
        );

    \I__743\ : InMux
    port map (
            O => \N__5259\,
            I => \N__5248\
        );

    \I__742\ : InMux
    port map (
            O => \N__5256\,
            I => \N__5245\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__5251\,
            I => \N__5242\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5248\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5245\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__738\ : Odrv4
    port map (
            O => \N__5242\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__5235\,
            I => \U712_CHIP_RAM.N_57_cascade_\
        );

    \I__736\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5229\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__5229\,
            I => \U712_CHIP_RAM.N_436\
        );

    \I__734\ : CascadeMux
    port map (
            O => \N__5226\,
            I => \U712_CHIP_RAM.N_436_cascade_\
        );

    \I__733\ : InMux
    port map (
            O => \N__5223\,
            I => \N__5220\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__5220\,
            I => \N__5217\
        );

    \I__731\ : Odrv4
    port map (
            O => \N__5217\,
            I => \U712_CHIP_RAM.N_83\
        );

    \I__730\ : InMux
    port map (
            O => \N__5214\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__729\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5207\
        );

    \I__728\ : InMux
    port map (
            O => \N__5210\,
            I => \N__5204\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__5207\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5204\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\
        );

    \I__725\ : InMux
    port map (
            O => \N__5199\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__724\ : InMux
    port map (
            O => \N__5196\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__723\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__5190\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__721\ : InMux
    port map (
            O => \N__5187\,
            I => \bfn_9_4_0_\
        );

    \I__720\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5180\
        );

    \I__719\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5177\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5180\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5177\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__716\ : InMux
    port map (
            O => \N__5172\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__715\ : InMux
    port map (
            O => \N__5169\,
            I => \N__5165\
        );

    \I__714\ : InMux
    port map (
            O => \N__5168\,
            I => \N__5162\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__5165\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__5162\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__711\ : InMux
    port map (
            O => \N__5157\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__710\ : InMux
    port map (
            O => \N__5154\,
            I => \N__5150\
        );

    \I__709\ : InMux
    port map (
            O => \N__5153\,
            I => \N__5147\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__5150\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__5147\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__706\ : InMux
    port map (
            O => \N__5142\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__705\ : CascadeMux
    port map (
            O => \N__5139\,
            I => \N__5135\
        );

    \I__704\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5132\
        );

    \I__703\ : InMux
    port map (
            O => \N__5135\,
            I => \N__5129\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5132\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5129\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__700\ : InMux
    port map (
            O => \N__5124\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__699\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5117\
        );

    \I__698\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5114\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5117\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5114\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__695\ : InMux
    port map (
            O => \N__5109\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__694\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5102\
        );

    \I__693\ : InMux
    port map (
            O => \N__5105\,
            I => \N__5099\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5102\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__5099\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__690\ : InMux
    port map (
            O => \N__5094\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__689\ : InMux
    port map (
            O => \N__5091\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__688\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5084\
        );

    \I__687\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5081\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5084\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__5081\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__684\ : ClkMux
    port map (
            O => \N__5076\,
            I => \N__5055\
        );

    \I__683\ : ClkMux
    port map (
            O => \N__5075\,
            I => \N__5055\
        );

    \I__682\ : ClkMux
    port map (
            O => \N__5074\,
            I => \N__5055\
        );

    \I__681\ : ClkMux
    port map (
            O => \N__5073\,
            I => \N__5055\
        );

    \I__680\ : ClkMux
    port map (
            O => \N__5072\,
            I => \N__5055\
        );

    \I__679\ : ClkMux
    port map (
            O => \N__5071\,
            I => \N__5055\
        );

    \I__678\ : ClkMux
    port map (
            O => \N__5070\,
            I => \N__5055\
        );

    \I__677\ : GlobalMux
    port map (
            O => \N__5055\,
            I => \N__5052\
        );

    \I__676\ : gio2CtrlBuf
    port map (
            O => \N__5052\,
            I => \C1_c_g\
        );

    \I__675\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5044\
        );

    \I__674\ : InMux
    port map (
            O => \N__5048\,
            I => \N__5041\
        );

    \I__673\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5038\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__5044\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_1\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__5041\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_1\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__5038\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_1\
        );

    \I__669\ : CascadeMux
    port map (
            O => \N__5031\,
            I => \U712_REG_SM.N_437_cascade_\
        );

    \I__668\ : InMux
    port map (
            O => \N__5028\,
            I => \N__5023\
        );

    \I__667\ : InMux
    port map (
            O => \N__5027\,
            I => \N__5018\
        );

    \I__666\ : InMux
    port map (
            O => \N__5026\,
            I => \N__5018\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5023\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__5018\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__663\ : InMux
    port map (
            O => \N__5013\,
            I => \N__5010\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__5010\,
            I => \U712_REG_SM.N_244\
        );

    \I__661\ : CascadeMux
    port map (
            O => \N__5007\,
            I => \U712_REG_SM.N_244_cascade_\
        );

    \I__660\ : InMux
    port map (
            O => \N__5004\,
            I => \N__5001\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__5001\,
            I => \U712_REG_SM.N_434\
        );

    \I__658\ : IoInMux
    port map (
            O => \N__4998\,
            I => \N__4995\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__4995\,
            I => \N__4991\
        );

    \I__656\ : IoInMux
    port map (
            O => \N__4994\,
            I => \N__4988\
        );

    \I__655\ : IoSpan4Mux
    port map (
            O => \N__4991\,
            I => \N__4985\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4988\,
            I => \N__4982\
        );

    \I__653\ : Span4Mux_s3_h
    port map (
            O => \N__4985\,
            I => \N__4979\
        );

    \I__652\ : IoSpan4Mux
    port map (
            O => \N__4982\,
            I => \N__4976\
        );

    \I__651\ : Sp12to4
    port map (
            O => \N__4979\,
            I => \N__4973\
        );

    \I__650\ : Span4Mux_s3_v
    port map (
            O => \N__4976\,
            I => \N__4970\
        );

    \I__649\ : Span12Mux_s11_h
    port map (
            O => \N__4973\,
            I => \N__4967\
        );

    \I__648\ : Span4Mux_v
    port map (
            O => \N__4970\,
            I => \N__4964\
        );

    \I__647\ : Span12Mux_v
    port map (
            O => \N__4967\,
            I => \N__4961\
        );

    \I__646\ : Sp12to4
    port map (
            O => \N__4964\,
            I => \N__4958\
        );

    \I__645\ : Odrv12
    port map (
            O => \N__4961\,
            I => \N_275\
        );

    \I__644\ : Odrv12
    port map (
            O => \N__4958\,
            I => \N_275\
        );

    \I__643\ : IoInMux
    port map (
            O => \N__4953\,
            I => \N__4950\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__4950\,
            I => \N__4947\
        );

    \I__641\ : Span12Mux_s11_h
    port map (
            O => \N__4947\,
            I => \N__4944\
        );

    \I__640\ : Span12Mux_v
    port map (
            O => \N__4944\,
            I => \N__4940\
        );

    \I__639\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4937\
        );

    \I__638\ : Odrv12
    port map (
            O => \N__4940\,
            I => \TACK_OUTn\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4937\,
            I => \TACK_OUTn\
        );

    \I__636\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4929\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4929\,
            I => \N__4926\
        );

    \I__634\ : Span4Mux_v
    port map (
            O => \N__4926\,
            I => \N__4922\
        );

    \I__633\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4919\
        );

    \I__632\ : Sp12to4
    port map (
            O => \N__4922\,
            I => \N__4914\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4919\,
            I => \N__4914\
        );

    \I__630\ : Span12Mux_h
    port map (
            O => \N__4914\,
            I => \N__4911\
        );

    \I__629\ : Span12Mux_v
    port map (
            O => \N__4911\,
            I => \N__4908\
        );

    \I__628\ : Odrv12
    port map (
            O => \N__4908\,
            I => \AWEn_c\
        );

    \I__627\ : InMux
    port map (
            O => \N__4905\,
            I => \N__4902\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__4902\,
            I => \N__4899\
        );

    \I__625\ : Odrv4
    port map (
            O => \N__4899\,
            I => \U712_CHIP_RAM.N_276\
        );

    \I__624\ : InMux
    port map (
            O => \N__4896\,
            I => \N__4893\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__4893\,
            I => \N__4889\
        );

    \I__622\ : InMux
    port map (
            O => \N__4892\,
            I => \N__4886\
        );

    \I__621\ : Odrv4
    port map (
            O => \N__4889\,
            I => \U712_CHIP_RAM.N_389\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__4886\,
            I => \U712_CHIP_RAM.N_389\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__4881\,
            I => \N__4878\
        );

    \I__618\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4875\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__4875\,
            I => \N__4872\
        );

    \I__616\ : Odrv12
    port map (
            O => \N__4872\,
            I => \U712_CHIP_RAM.N_300\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__4869\,
            I => \U712_REG_SM.N_277_cascade_\
        );

    \I__614\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4862\
        );

    \I__613\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4859\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4862\,
            I => \U712_REG_SM.N_236\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__4859\,
            I => \U712_REG_SM.N_236\
        );

    \I__610\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4851\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__4851\,
            I => \U712_REG_SM.N_277\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__4848\,
            I => \U712_REG_SM.N_236_cascade_\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__4845\,
            I => \U712_CHIP_RAM.N_374_cascade_\
        );

    \I__606\ : InMux
    port map (
            O => \N__4842\,
            I => \N__4835\
        );

    \I__605\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4835\
        );

    \I__604\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4832\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__4835\,
            I => \U712_CHIP_RAM.N_418\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4832\,
            I => \U712_CHIP_RAM.N_418\
        );

    \I__601\ : InMux
    port map (
            O => \N__4827\,
            I => \N__4824\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__4824\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__4821\,
            I => \U712_CHIP_RAM.N_418_cascade_\
        );

    \I__598\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4815\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4815\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_0_a2_1_a2_0\
        );

    \I__596\ : InMux
    port map (
            O => \N__4812\,
            I => \N__4809\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4809\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__594\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4798\
        );

    \I__593\ : InMux
    port map (
            O => \N__4805\,
            I => \N__4798\
        );

    \I__592\ : InMux
    port map (
            O => \N__4804\,
            I => \N__4793\
        );

    \I__591\ : InMux
    port map (
            O => \N__4803\,
            I => \N__4793\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__4798\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4793\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__588\ : InMux
    port map (
            O => \N__4788\,
            I => \N__4781\
        );

    \I__587\ : InMux
    port map (
            O => \N__4787\,
            I => \N__4781\
        );

    \I__586\ : InMux
    port map (
            O => \N__4786\,
            I => \N__4778\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__4781\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4778\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__583\ : InMux
    port map (
            O => \N__4773\,
            I => \N__4769\
        );

    \I__582\ : InMux
    port map (
            O => \N__4772\,
            I => \N__4766\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__4769\,
            I => \U712_CHIP_RAM.N_229\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4766\,
            I => \U712_CHIP_RAM.N_229\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__4761\,
            I => \U712_CHIP_RAM.N_389_cascade_\
        );

    \I__578\ : InMux
    port map (
            O => \N__4758\,
            I => \N__4755\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__4755\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__576\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4749\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4749\,
            I => \U712_CHIP_RAM.REFRESH5lto7_0\
        );

    \I__574\ : CascadeMux
    port map (
            O => \N__4746\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_0_0_1_cascade_\
        );

    \I__573\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4740\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4740\,
            I => \N__4737\
        );

    \I__571\ : Span4Mux_h
    port map (
            O => \N__4737\,
            I => \N__4734\
        );

    \I__570\ : Sp12to4
    port map (
            O => \N__4734\,
            I => \N__4731\
        );

    \I__569\ : Span12Mux_v
    port map (
            O => \N__4731\,
            I => \N__4728\
        );

    \I__568\ : Odrv12
    port map (
            O => \N__4728\,
            I => \A_c_20\
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__4725\,
            I => \U712_CHIP_RAM.N_323_cascade_\
        );

    \I__566\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4718\
        );

    \I__565\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4715\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4718\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4715\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\
        );

    \I__562\ : IoInMux
    port map (
            O => \N__4710\,
            I => \N__4707\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__4707\,
            I => \N__4704\
        );

    \I__560\ : Span4Mux_s3_v
    port map (
            O => \N__4704\,
            I => \N__4701\
        );

    \I__559\ : Span4Mux_v
    port map (
            O => \N__4701\,
            I => \N__4698\
        );

    \I__558\ : Span4Mux_h
    port map (
            O => \N__4698\,
            I => \N__4695\
        );

    \I__557\ : Odrv4
    port map (
            O => \N__4695\,
            I => \BANK0_c\
        );

    \I__556\ : CEMux
    port map (
            O => \N__4692\,
            I => \N__4689\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4689\,
            I => \N__4686\
        );

    \I__554\ : Span4Mux_h
    port map (
            O => \N__4686\,
            I => \N__4683\
        );

    \I__553\ : Odrv4
    port map (
            O => \N__4683\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0\
        );

    \I__552\ : CascadeMux
    port map (
            O => \N__4680\,
            I => \U712_CHIP_RAM.N_367_cascade_\
        );

    \I__551\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4674\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4674\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a3_0\
        );

    \I__549\ : InMux
    port map (
            O => \N__4671\,
            I => \N__4668\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4668\,
            I => \N__4664\
        );

    \I__547\ : IoInMux
    port map (
            O => \N__4667\,
            I => \N__4661\
        );

    \I__546\ : Span4Mux_v
    port map (
            O => \N__4664\,
            I => \N__4658\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__4661\,
            I => \N__4655\
        );

    \I__544\ : Sp12to4
    port map (
            O => \N__4658\,
            I => \N__4652\
        );

    \I__543\ : IoSpan4Mux
    port map (
            O => \N__4655\,
            I => \N__4649\
        );

    \I__542\ : Span12Mux_h
    port map (
            O => \N__4652\,
            I => \N__4646\
        );

    \I__541\ : IoSpan4Mux
    port map (
            O => \N__4649\,
            I => \N__4643\
        );

    \I__540\ : Span12Mux_v
    port map (
            O => \N__4646\,
            I => \N__4640\
        );

    \I__539\ : IoSpan4Mux
    port map (
            O => \N__4643\,
            I => \N__4637\
        );

    \I__538\ : Odrv12
    port map (
            O => \N__4640\,
            I => \C1_c\
        );

    \I__537\ : Odrv4
    port map (
            O => \N__4637\,
            I => \C1_c\
        );

    \I__536\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4629\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4629\,
            I => \N__4626\
        );

    \I__534\ : Odrv4
    port map (
            O => \N__4626\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__533\ : CascadeMux
    port map (
            O => \N__4623\,
            I => \N__4620\
        );

    \I__532\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4617\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__4617\,
            I => \N__4614\
        );

    \I__530\ : Span4Mux_v
    port map (
            O => \N__4614\,
            I => \N__4610\
        );

    \I__529\ : InMux
    port map (
            O => \N__4613\,
            I => \N__4607\
        );

    \I__528\ : Sp12to4
    port map (
            O => \N__4610\,
            I => \N__4602\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4607\,
            I => \N__4602\
        );

    \I__526\ : Span12Mux_h
    port map (
            O => \N__4602\,
            I => \N__4599\
        );

    \I__525\ : Span12Mux_v
    port map (
            O => \N__4599\,
            I => \N__4596\
        );

    \I__524\ : Odrv12
    port map (
            O => \N__4596\,
            I => \TSn_c\
        );

    \I__523\ : InMux
    port map (
            O => \N__4593\,
            I => \N__4590\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4590\,
            I => \N__4587\
        );

    \I__521\ : Span12Mux_v
    port map (
            O => \N__4587\,
            I => \N__4584\
        );

    \I__520\ : Odrv12
    port map (
            O => \N__4584\,
            I => \RAMSPACEn_c\
        );

    \I__519\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4578\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4578\,
            I => \N__4575\
        );

    \I__517\ : Span12Mux_v
    port map (
            O => \N__4575\,
            I => \N__4572\
        );

    \I__516\ : Odrv12
    port map (
            O => \N__4572\,
            I => \U712_CHIP_RAM.N_360\
        );

    \I__515\ : IoInMux
    port map (
            O => \N__4569\,
            I => \N__4566\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__4566\,
            I => \N__4563\
        );

    \I__513\ : Span12Mux_s8_v
    port map (
            O => \N__4563\,
            I => \N__4560\
        );

    \I__512\ : Odrv12
    port map (
            O => \N__4560\,
            I => \VBENn_c\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__4557\,
            I => \U712_CHIP_RAM.N_239_cascade_\
        );

    \I__510\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4550\
        );

    \I__509\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4547\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4550\,
            I => \LATCH_REG\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__4547\,
            I => \LATCH_REG\
        );

    \I__506\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4539\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4539\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__504\ : InMux
    port map (
            O => \N__4536\,
            I => \N__4533\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4533\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_0\
        );

    \I__502\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4521\
        );

    \I__501\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4521\
        );

    \I__500\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4521\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4521\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_1\
        );

    \I__498\ : IoInMux
    port map (
            O => \N__4518\,
            I => \N__4515\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4515\,
            I => \N__4512\
        );

    \I__496\ : IoSpan4Mux
    port map (
            O => \N__4512\,
            I => \N__4509\
        );

    \I__495\ : Span4Mux_s3_v
    port map (
            O => \N__4509\,
            I => \N__4506\
        );

    \I__494\ : Sp12to4
    port map (
            O => \N__4506\,
            I => \N__4503\
        );

    \I__493\ : Span12Mux_v
    port map (
            O => \N__4503\,
            I => \N__4499\
        );

    \I__492\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4496\
        );

    \I__491\ : Odrv12
    port map (
            O => \N__4499\,
            I => \REGENn_c\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4496\,
            I => \REGENn_c\
        );

    \I__489\ : IoInMux
    port map (
            O => \N__4491\,
            I => \N__4488\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4488\,
            I => \N__4485\
        );

    \I__487\ : Span4Mux_s2_v
    port map (
            O => \N__4485\,
            I => \N__4482\
        );

    \I__486\ : Span4Mux_h
    port map (
            O => \N__4482\,
            I => \N__4479\
        );

    \I__485\ : Span4Mux_h
    port map (
            O => \N__4479\,
            I => \N__4476\
        );

    \I__484\ : Span4Mux_v
    port map (
            O => \N__4476\,
            I => \N__4473\
        );

    \I__483\ : Sp12to4
    port map (
            O => \N__4473\,
            I => \N__4470\
        );

    \I__482\ : Span12Mux_v
    port map (
            O => \N__4470\,
            I => \N__4466\
        );

    \I__481\ : InMux
    port map (
            O => \N__4469\,
            I => \N__4463\
        );

    \I__480\ : Odrv12
    port map (
            O => \N__4466\,
            I => \ASn_c\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4463\,
            I => \ASn_c\
        );

    \I__478\ : InMux
    port map (
            O => \N__4458\,
            I => \N__4455\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4455\,
            I => \N__4452\
        );

    \I__476\ : Span4Mux_v
    port map (
            O => \N__4452\,
            I => \N__4449\
        );

    \I__475\ : Span4Mux_h
    port map (
            O => \N__4449\,
            I => \N__4446\
        );

    \I__474\ : Sp12to4
    port map (
            O => \N__4446\,
            I => \N__4443\
        );

    \I__473\ : Span12Mux_v
    port map (
            O => \N__4443\,
            I => \N__4440\
        );

    \I__472\ : Odrv12
    port map (
            O => \N__4440\,
            I => \REGSPACEn_c\
        );

    \I__471\ : InMux
    port map (
            O => \N__4437\,
            I => \N__4431\
        );

    \I__470\ : InMux
    port map (
            O => \N__4436\,
            I => \N__4431\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4431\,
            I => \U712_REG_SM.CYCLE_RUNZ0\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__4428\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_\
        );

    \I__467\ : IoInMux
    port map (
            O => \N__4425\,
            I => \N__4422\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4422\,
            I => \N__4419\
        );

    \I__465\ : Span12Mux_s4_v
    port map (
            O => \N__4419\,
            I => \N__4415\
        );

    \I__464\ : InMux
    port map (
            O => \N__4418\,
            I => \N__4412\
        );

    \I__463\ : Odrv12
    port map (
            O => \N__4415\,
            I => \DBDIR_c\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4412\,
            I => \DBDIR_c\
        );

    \I__461\ : InMux
    port map (
            O => \N__4407\,
            I => \N__4404\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4404\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0\
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__4401\,
            I => \U712_CHIP_RAM.DBENn_8_0_cascade_\
        );

    \I__458\ : CascadeMux
    port map (
            O => \N__4398\,
            I => \N__4395\
        );

    \I__457\ : InMux
    port map (
            O => \N__4395\,
            I => \N__4392\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__4392\,
            I => \U712_CHIP_RAM.N_316\
        );

    \I__455\ : InMux
    port map (
            O => \N__4389\,
            I => \N__4386\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__4386\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\
        );

    \I__453\ : InMux
    port map (
            O => \N__4383\,
            I => \N__4379\
        );

    \I__452\ : InMux
    port map (
            O => \N__4382\,
            I => \N__4376\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__4379\,
            I => \N__4373\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4376\,
            I => \N__4370\
        );

    \I__449\ : Span4Mux_v
    port map (
            O => \N__4373\,
            I => \N__4364\
        );

    \I__448\ : Span4Mux_v
    port map (
            O => \N__4370\,
            I => \N__4364\
        );

    \I__447\ : InMux
    port map (
            O => \N__4369\,
            I => \N__4361\
        );

    \I__446\ : Sp12to4
    port map (
            O => \N__4364\,
            I => \N__4356\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4361\,
            I => \N__4356\
        );

    \I__444\ : Span12Mux_h
    port map (
            O => \N__4356\,
            I => \N__4353\
        );

    \I__443\ : Span12Mux_v
    port map (
            O => \N__4353\,
            I => \N__4350\
        );

    \I__442\ : Odrv12
    port map (
            O => \N__4350\,
            I => \DBRn_c\
        );

    \I__441\ : CascadeMux
    port map (
            O => \N__4347\,
            I => \U712_CHIP_RAM.N_229_cascade_\
        );

    \I__440\ : InMux
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4341\,
            I => \U712_CHIP_RAM.N_345_1\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__4338\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_\
        );

    \I__437\ : InMux
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4332\,
            I => \N__4328\
        );

    \I__435\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4325\
        );

    \I__434\ : Odrv4
    port map (
            O => \N__4328\,
            I => \LATCH_RAM\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__4325\,
            I => \LATCH_RAM\
        );

    \I__432\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4317\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__4317\,
            I => \U712_CHIP_RAM.N_379\
        );

    \I__430\ : CascadeMux
    port map (
            O => \N__4314\,
            I => \U712_CHIP_RAM.N_316_cascade_\
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__4311\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_\
        );

    \I__428\ : IoInMux
    port map (
            O => \N__4308\,
            I => \N__4305\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__4305\,
            I => \N__4302\
        );

    \I__426\ : IoSpan4Mux
    port map (
            O => \N__4302\,
            I => \N__4299\
        );

    \I__425\ : Span4Mux_s3_h
    port map (
            O => \N__4299\,
            I => \N__4296\
        );

    \I__424\ : Span4Mux_h
    port map (
            O => \N__4296\,
            I => \N__4292\
        );

    \I__423\ : InMux
    port map (
            O => \N__4295\,
            I => \N__4289\
        );

    \I__422\ : Span4Mux_h
    port map (
            O => \N__4292\,
            I => \N__4286\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__4289\,
            I => \N__4283\
        );

    \I__420\ : Span4Mux_h
    port map (
            O => \N__4286\,
            I => \N__4280\
        );

    \I__419\ : Span4Mux_v
    port map (
            O => \N__4283\,
            I => \N__4277\
        );

    \I__418\ : Sp12to4
    port map (
            O => \N__4280\,
            I => \N__4272\
        );

    \I__417\ : Sp12to4
    port map (
            O => \N__4277\,
            I => \N__4272\
        );

    \I__416\ : Span12Mux_h
    port map (
            O => \N__4272\,
            I => \N__4269\
        );

    \I__415\ : Span12Mux_v
    port map (
            O => \N__4269\,
            I => \N__4266\
        );

    \I__414\ : Odrv12
    port map (
            O => \N__4266\,
            I => \C3_c\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__4263\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_\
        );

    \I__412\ : CascadeMux
    port map (
            O => \N__4260\,
            I => \U712_CHIP_RAM.N_390_cascade_\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__4257\,
            I => \N__4254\
        );

    \I__410\ : InMux
    port map (
            O => \N__4254\,
            I => \N__4251\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__4251\,
            I => \U712_CHIP_RAM.N_346\
        );

    \I__408\ : InMux
    port map (
            O => \N__4248\,
            I => \N__4242\
        );

    \I__407\ : InMux
    port map (
            O => \N__4247\,
            I => \N__4242\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__4242\,
            I => \U712_CHIP_RAM.N_319\
        );

    \I__405\ : IoInMux
    port map (
            O => \N__4239\,
            I => \N__4236\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4236\,
            I => \N__4232\
        );

    \I__403\ : IoInMux
    port map (
            O => \N__4235\,
            I => \N__4229\
        );

    \I__402\ : Span12Mux_s0_v
    port map (
            O => \N__4232\,
            I => \N__4225\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__4229\,
            I => \N__4222\
        );

    \I__400\ : IoInMux
    port map (
            O => \N__4228\,
            I => \N__4219\
        );

    \I__399\ : Span12Mux_v
    port map (
            O => \N__4225\,
            I => \N__4216\
        );

    \I__398\ : Span12Mux_s6_v
    port map (
            O => \N__4222\,
            I => \N__4213\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__4219\,
            I => \N__4210\
        );

    \I__396\ : Span12Mux_h
    port map (
            O => \N__4216\,
            I => \N__4207\
        );

    \I__395\ : Span12Mux_h
    port map (
            O => \N__4213\,
            I => \N__4204\
        );

    \I__394\ : Span4Mux_s3_h
    port map (
            O => \N__4210\,
            I => \N__4201\
        );

    \I__393\ : Span12Mux_h
    port map (
            O => \N__4207\,
            I => \N__4198\
        );

    \I__392\ : Span12Mux_h
    port map (
            O => \N__4204\,
            I => \N__4195\
        );

    \I__391\ : Span4Mux_v
    port map (
            O => \N__4201\,
            I => \N__4192\
        );

    \I__390\ : Odrv12
    port map (
            O => \N__4198\,
            I => \CLK40_PLL_iso_i\
        );

    \I__389\ : Odrv12
    port map (
            O => \N__4195\,
            I => \CLK40_PLL_iso_i\
        );

    \I__388\ : Odrv4
    port map (
            O => \N__4192\,
            I => \CLK40_PLL_iso_i\
        );

    \I__387\ : IoInMux
    port map (
            O => \N__4185\,
            I => \N__4182\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__4182\,
            I => \N__4179\
        );

    \I__385\ : Span4Mux_s1_h
    port map (
            O => \N__4179\,
            I => \N__4176\
        );

    \I__384\ : Span4Mux_h
    port map (
            O => \N__4176\,
            I => \N__4173\
        );

    \I__383\ : Odrv4
    port map (
            O => \N__4173\,
            I => \DBRn_c_i_0\
        );

    \I__382\ : IoInMux
    port map (
            O => \N__4170\,
            I => \N__4167\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__4167\,
            I => \N__4164\
        );

    \I__380\ : Span4Mux_s3_h
    port map (
            O => \N__4164\,
            I => \N__4161\
        );

    \I__379\ : Span4Mux_v
    port map (
            O => \N__4161\,
            I => \N__4158\
        );

    \I__378\ : Odrv4
    port map (
            O => \N__4158\,
            I => \N_929_i\
        );

    \I__377\ : IoInMux
    port map (
            O => \N__4155\,
            I => \N__4152\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__4152\,
            I => \N__4149\
        );

    \I__375\ : Span4Mux_s2_v
    port map (
            O => \N__4149\,
            I => \N__4146\
        );

    \I__374\ : Span4Mux_v
    port map (
            O => \N__4146\,
            I => \N__4143\
        );

    \I__373\ : Span4Mux_h
    port map (
            O => \N__4143\,
            I => \N__4140\
        );

    \I__372\ : Odrv4
    port map (
            O => \N__4140\,
            I => \CLK80_PLL_i_i\
        );

    \I__371\ : IoInMux
    port map (
            O => \N__4137\,
            I => \N__4134\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__4134\,
            I => \N__4131\
        );

    \I__369\ : IoSpan4Mux
    port map (
            O => \N__4131\,
            I => \N__4128\
        );

    \I__368\ : Sp12to4
    port map (
            O => \N__4128\,
            I => \N__4125\
        );

    \I__367\ : Span12Mux_v
    port map (
            O => \N__4125\,
            I => \N__4122\
        );

    \I__366\ : Odrv12
    port map (
            O => \N__4122\,
            I => \LATCH_CLK_0_i\
        );

    \I__365\ : IoInMux
    port map (
            O => \N__4119\,
            I => \N__4116\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__4116\,
            I => \N__4113\
        );

    \I__363\ : Span4Mux_s0_v
    port map (
            O => \N__4113\,
            I => \N__4110\
        );

    \I__362\ : Span4Mux_v
    port map (
            O => \N__4110\,
            I => \N__4107\
        );

    \I__361\ : Sp12to4
    port map (
            O => \N__4107\,
            I => \N__4104\
        );

    \I__360\ : Span12Mux_h
    port map (
            O => \N__4104\,
            I => \N__4101\
        );

    \I__359\ : Span12Mux_v
    port map (
            O => \N__4101\,
            I => \N__4098\
        );

    \I__358\ : Odrv12
    port map (
            O => \N__4098\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__5075\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__5072\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__5073\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__5074\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__5070\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__5071\
        );

    \INVU712_REG_SM.LDSnC\ : INV
    port map (
            O => \INVU712_REG_SM.LDSnC_net\,
            I => \N__6528\
        );

    \INVU712_REG_SM.STATE_COUNTER_5C\ : INV
    port map (
            O => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            I => \N__6530\
        );

    \INVU712_REG_SM.C1_SYNC_0C\ : INV
    port map (
            O => \INVU712_REG_SM.C1_SYNC_0C_net\,
            I => \N__6527\
        );

    \INVU712_REG_SM.C3_SYNC_1C\ : INV
    port map (
            O => \INVU712_REG_SM.C3_SYNC_1C_net\,
            I => \N__6529\
        );

    \INVU712_REG_SM.C1_SYNC_1C\ : INV
    port map (
            O => \INVU712_REG_SM.C1_SYNC_1C_net\,
            I => \N__6532\
        );

    \INVU712_REG_SM.C3_SYNC_0C\ : INV
    port map (
            O => \INVU712_REG_SM.C3_SYNC_0C_net\,
            I => \N__6531\
        );

    \IN_MUX_bfv_9_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_4_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_6_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4667\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \CLK40_PLL_derived_clock_RNIIOT\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7828\,
            GLOBALBUFFEROUTPUT => \CLK40_PLL_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8154\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4185\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4308\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLK40_PLL_derived_clock_RNIIOT_0_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6543\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_iso_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11253\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8894\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6765\,
            lcout => \N_929_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10683\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4369\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.LATCH_CLK_0_i_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__4335\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4554\,
            lcout => \LATCH_CLK_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4295\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_0C_net\,
            ce => 'H',
            sr => \N__11204\
        );

    \U712_REG_SM.DBR_SYNC_0_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4382\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_0C_net\,
            ce => 'H',
            sr => \N__11204\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__5899\,
            in1 => \N__4247\,
            in2 => \N__4257\,
            in3 => \N__4344\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11252\,
            in1 => \_gnd_net_\,
            in2 => \N__4263\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_5_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7291\,
            in2 => \_gnd_net_\,
            in3 => \N__6636\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_390_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_4_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8471\,
            in1 => \N__5386\,
            in2 => \N__4260\,
            in3 => \N__5898\,
            lcout => \U712_CHIP_RAM.N_346\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001000"
        )
    port map (
            in0 => \N__4248\,
            in1 => \N__4721\,
            in2 => \N__7171\,
            in3 => \N__10767\,
            lcout => \CPU_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10665\,
            ce => 'H',
            sr => \N__11224\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__4804\,
            in1 => \N__8289\,
            in2 => \N__10848\,
            in3 => \N__4581\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10670\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__7282\,
            in1 => \N__6314\,
            in2 => \_gnd_net_\,
            in3 => \N__4840\,
            lcout => \U712_CHIP_RAM.N_319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_0_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__4803\,
            in1 => \N__4786\,
            in2 => \N__5264\,
            in3 => \N__5343\,
            lcout => \U712_CHIP_RAM.N_229\,
            ltout => \U712_CHIP_RAM.N_229_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7366\,
            in2 => \N__4347\,
            in3 => \N__5387\,
            lcout => \U712_CHIP_RAM.N_345_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5388\,
            in1 => \N__7380\,
            in2 => \N__7173\,
            in3 => \N__4773\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8293\,
            in1 => \N__4905\,
            in2 => \N__4338\,
            in3 => \N__6315\,
            lcout => \WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10670\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIC9HD1_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6635\,
            in1 => \N__7281\,
            in2 => \_gnd_net_\,
            in3 => \N__5342\,
            lcout => \U712_CHIP_RAM.N_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_RAM_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011000000"
        )
    port map (
            in0 => \N__5223\,
            in1 => \N__4331\,
            in2 => \N__8302\,
            in3 => \N__4389\,
            lcout => \LATCH_RAM\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10670\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKV5I5_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__5415\,
            in1 => \N__5389\,
            in2 => \N__7172\,
            in3 => \N__4320\,
            lcout => \U712_CHIP_RAM.N_316\,
            ltout => \U712_CHIP_RAM.N_316_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNICBGO9_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__7289\,
            in1 => \N__6329\,
            in2 => \N__4314\,
            in3 => \N__4841\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4311\,
            in3 => \N__11251\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5349\,
            in1 => \N__7164\,
            in2 => \N__5401\,
            in3 => \N__7386\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBDIR_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101111101010000"
        )
    port map (
            in0 => \N__4925\,
            in1 => \_gnd_net_\,
            in2 => \N__4428\,
            in3 => \N__4418\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10674\,
            ce => 'H',
            sr => \N__11216\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5393\,
            in1 => \N__7385\,
            in2 => \_gnd_net_\,
            in3 => \N__9906\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.DBENn_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4407\,
            in2 => \N__4401\,
            in3 => \N__8350\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10674\,
            ce => 'H',
            sr => \N__11216\
        );

    \U712_CHIP_RAM.LATCH_RAM_RNO_1_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__7290\,
            in1 => \N__4842\,
            in2 => \N__4398\,
            in3 => \N__6330\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_0_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4383\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10677\,
            ce => 'H',
            sr => \N__11211\
        );

    \U712_REG_SM.C1_SYNC_1_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4632\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C1_SYNC_1C_net\,
            ce => 'H',
            sr => \N__11205\
        );

    \U712_REG_SM.REG_CYCLE_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__10987\,
            in1 => \N__6008\,
            in2 => \_gnd_net_\,
            in3 => \N__5957\,
            lcout => \REG_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C1_SYNC_1C_net\,
            ce => 'H',
            sr => \N__11205\
        );

    \U712_REG_SM.STATE_COUNTER_0_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__5955\,
            in1 => \N__6140\,
            in2 => \_gnd_net_\,
            in3 => \N__6185\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C1_SYNC_1C_net\,
            ce => 'H',
            sr => \N__11205\
        );

    \U712_REG_SM.STATE_COUNTER_3_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6097\,
            in1 => \N__5609\,
            in2 => \N__5661\,
            in3 => \N__5049\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C1_SYNC_1C_net\,
            ce => 'H',
            sr => \N__11205\
        );

    \U712_REG_SM.LATCH_REG_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010111000000"
        )
    port map (
            in0 => \N__5956\,
            in1 => \N__6043\,
            in2 => \N__5843\,
            in3 => \N__4553\,
            lcout => \LATCH_REG\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C1_SYNC_1C_net\,
            ce => 'H',
            sr => \N__11205\
        );

    \U712_REG_SM.C3_SYNC_1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4542\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_1C_net\,
            ce => 'H',
            sr => \N__11197\
        );

    \U712_REG_SM.STATE_COUNTER_1_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__6184\,
            in1 => \N__6138\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_1C_net\,
            ce => 'H',
            sr => \N__11197\
        );

    \U712_REG_SM.STATE_COUNTER_2_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011011100"
        )
    port map (
            in0 => \N__5048\,
            in1 => \N__4530\,
            in2 => \N__6099\,
            in3 => \N__4866\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_1C_net\,
            ce => 'H',
            sr => \N__11197\
        );

    \U712_REG_SM.CYCLE_RUN_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100110000"
        )
    port map (
            in0 => \N__4528\,
            in1 => \N__6139\,
            in2 => \N__6197\,
            in3 => \N__4436\,
            lcout => \U712_REG_SM.CYCLE_RUNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_1C_net\,
            ce => 'H',
            sr => \N__11197\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4536\,
            lcout => \U712_REG_SM.DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_1C_net\,
            ce => 'H',
            sr => \N__11197\
        );

    \U712_REG_SM.REGENn_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__4529\,
            in1 => \N__5966\,
            in2 => \_gnd_net_\,
            in3 => \N__4502\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_1C_net\,
            ce => 'H',
            sr => \N__11197\
        );

    \U712_REG_SM.ASn_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__5013\,
            in1 => \N__5659\,
            in2 => \N__5967\,
            in3 => \N__4469\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_1C_net\,
            ce => 'H',
            sr => \N__11197\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__4458\,
            in1 => \N__4437\,
            in2 => \N__4623\,
            in3 => \N__5028\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_1C_net\,
            ce => 'H',
            sr => \N__11197\
        );

    \U712_REG_SM.C1_SYNC_0_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4671\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C1_SYNC_0C_net\,
            ce => 'H',
            sr => \N__11192\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4613\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4593\,
            lcout => \U712_CHIP_RAM.N_360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__5153\,
            in1 => \N__5168\,
            in2 => \N__5139\,
            in3 => \N__5183\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5685\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10771\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5105\,
            in2 => \_gnd_net_\,
            in3 => \N__5120\,
            lcout => \U712_CHIP_RAM.REFRESH5lto7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__7096\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6968\,
            lcout => \U712_CHIP_RAM.N_300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAQ_4_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7017\,
            in2 => \_gnd_net_\,
            in3 => \N__7095\,
            lcout => \U712_CHIP_RAM.N_239\,
            ltout => \U712_CHIP_RAM.N_239_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI4LVP1_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000101"
        )
    port map (
            in0 => \N__6612\,
            in1 => \N__8459\,
            in2 => \N__4557\,
            in3 => \N__7272\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7271\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6611\,
            lcout => \U712_CHIP_RAM.N_228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__5088\,
            in1 => \N__4758\,
            in2 => \N__8304\,
            in3 => \N__4752\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10659\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJHLS1_1_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101001111"
        )
    port map (
            in0 => \N__7270\,
            in1 => \N__6610\,
            in2 => \N__8303\,
            in3 => \N__6466\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNINIA74_1_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__6467\,
            in1 => \N__6892\,
            in2 => \N__4746\,
            in3 => \N__6262\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110001000"
        )
    port map (
            in0 => \N__8295\,
            in1 => \N__7923\,
            in2 => \N__8470\,
            in3 => \N__5336\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10659\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIURFN4_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4818\,
            in1 => \N__7364\,
            in2 => \_gnd_net_\,
            in3 => \N__5402\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7365\,
            in1 => \N__5335\,
            in2 => \N__5406\,
            in3 => \N__8871\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__10140\,
            in1 => \N__4743\,
            in2 => \N__4725\,
            in3 => \N__4722\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10666\,
            ce => \N__4692\,
            sr => \N__11217\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_1_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6934\,
            in1 => \N__6469\,
            in2 => \_gnd_net_\,
            in3 => \N__6261\,
            lcout => \U712_CHIP_RAM.N_367\,
            ltout => \U712_CHIP_RAM.N_367_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNITGCI5_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101110101"
        )
    port map (
            in0 => \N__8240\,
            in1 => \N__7363\,
            in2 => \N__4680\,
            in3 => \N__4677\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_1_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6613\,
            in1 => \N__6468\,
            in2 => \_gnd_net_\,
            in3 => \N__6260\,
            lcout => \U712_CHIP_RAM.N_374\,
            ltout => \U712_CHIP_RAM.N_374_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5897\,
            in2 => \N__4845\,
            in3 => \N__6935\,
            lcout => \U712_CHIP_RAM.N_418\,
            ltout => \U712_CHIP_RAM.N_418_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIQG71D_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__6341\,
            in1 => \N__4827\,
            in2 => \N__4821\,
            in3 => \N__5232\,
            lcout => \U712_CHIP_RAM.N_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_1_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__4788\,
            in1 => \N__5263\,
            in2 => \N__5348\,
            in3 => \N__4806\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_0_a2_1_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_1_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4812\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10671\,
            ce => 'H',
            sr => \N__11212\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__4805\,
            in1 => \N__4787\,
            in2 => \N__5265\,
            in3 => \N__5337\,
            lcout => \U712_CHIP_RAM.N_278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFMOI5_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4772\,
            in1 => \N__4892\,
            in2 => \_gnd_net_\,
            in3 => \N__7149\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_1_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8288\,
            in1 => \N__7384\,
            in2 => \_gnd_net_\,
            in3 => \N__5394\,
            lcout => \U712_CHIP_RAM.N_389\,
            ltout => \U712_CHIP_RAM.N_389_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIGGM16_4_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100111111"
        )
    port map (
            in0 => \N__7418\,
            in1 => \N__7028\,
            in2 => \N__4761\,
            in3 => \N__7148\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__7509\,
            in1 => \N__7570\,
            in2 => \N__7683\,
            in3 => \N__7649\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10675\,
            ce => 'H',
            sr => \N__11206\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110001100"
        )
    port map (
            in0 => \N__7833\,
            in1 => \N__4943\,
            in2 => \N__7572\,
            in3 => \N__7530\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10675\,
            ce => 'H',
            sr => \N__11206\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__5344\,
            in1 => \N__4932\,
            in2 => \_gnd_net_\,
            in3 => \N__6237\,
            lcout => \U712_CHIP_RAM.N_276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5833\,
            in1 => \N__6118\,
            in2 => \_gnd_net_\,
            in3 => \N__5562\,
            lcout => \U712_REG_SM.un15_0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__6822\,
            in1 => \N__4896\,
            in2 => \N__4881\,
            in3 => \N__5499\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10678\,
            ce => \N__5442\,
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_RNI5J3V_7_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__6229\,
            in1 => \N__5557\,
            in2 => \_gnd_net_\,
            in3 => \N__6177\,
            lcout => \U712_REG_SM.N_277\,
            ltout => \U712_REG_SM.N_277_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_RNO_1_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5707\,
            in1 => \N__4865\,
            in2 => \N__4869\,
            in3 => \N__6092\,
            lcout => \U712_REG_SM.UDSn_7_iv_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5610\,
            in2 => \_gnd_net_\,
            in3 => \N__5648\,
            lcout => \U712_REG_SM.N_236\,
            ltout => \U712_REG_SM.N_236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_1_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__4854\,
            in1 => \N__5773\,
            in2 => \N__4848\,
            in3 => \N__6093\,
            lcout => \U712_REG_SM.LDSn_7_iv_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_RNIELLV_7_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5611\,
            in1 => \N__5558\,
            in2 => \_gnd_net_\,
            in3 => \N__5649\,
            lcout => \U712_REG_SM.LATCH_REG_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_RNO_0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__9776\,
            in1 => \N__5004\,
            in2 => \N__6203\,
            in3 => \N__9667\,
            lcout => \U712_REG_SM.N_337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNIPBK41_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__5652\,
            in1 => \N__5605\,
            in2 => \_gnd_net_\,
            in3 => \N__5027\,
            lcout => \U712_REG_SM.N_255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6086\,
            in1 => \N__5047\,
            in2 => \N__5612\,
            in3 => \N__5650\,
            lcout => \U712_REG_SM.STATE_COUNTERc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_2_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5772\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6087\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_437_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__9775\,
            in1 => \N__9666\,
            in2 => \N__5031\,
            in3 => \N__6199\,
            lcout => \U712_REG_SM.N_339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNIGHT91_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__6198\,
            in1 => \N__5604\,
            in2 => \N__5567\,
            in3 => \N__5026\,
            lcout => \U712_REG_SM.N_244\,
            ltout => \U712_REG_SM.N_244_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI5ITS1_1_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111010"
        )
    port map (
            in0 => \N__6088\,
            in1 => \_gnd_net_\,
            in2 => \N__5007\,
            in3 => \N__5651\,
            lcout => \U712_REG_SM.N_169\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_RNO_2_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5706\,
            in2 => \_gnd_net_\,
            in3 => \N__6085\,
            lcout => \U712_REG_SM.N_434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DMA_LATCH_EN_1_i_m2_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__6045\,
            in1 => \N__10994\,
            in2 => \_gnd_net_\,
            in3 => \N__6348\,
            lcout => \N_275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5193\,
            in2 => \_gnd_net_\,
            in3 => \N__5187\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_9_4_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__5076\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5184\,
            in2 => \_gnd_net_\,
            in3 => \N__5172\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__5076\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5169\,
            in2 => \_gnd_net_\,
            in3 => \N__5157\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__5076\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5154\,
            in2 => \_gnd_net_\,
            in3 => \N__5142\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__5076\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5138\,
            in2 => \_gnd_net_\,
            in3 => \N__5124\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__5076\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5121\,
            in2 => \_gnd_net_\,
            in3 => \N__5109\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__5076\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5106\,
            in2 => \_gnd_net_\,
            in3 => \N__5094\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__5076\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5087\,
            in2 => \_gnd_net_\,
            in3 => \N__5091\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5076\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_RNIRILU_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__5331\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5259\,
            lcout => \U712_CHIP_RAM.N_263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5453\,
            in1 => \N__5513\,
            in2 => \_gnd_net_\,
            in3 => \N__5528\,
            lcout => \U712_CHIP_RAM.N_57\,
            ltout => \U712_CHIP_RAM.N_57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__6937\,
            in1 => \N__6624\,
            in2 => \N__5235\,
            in3 => \N__7108\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_4_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__7435\,
            in1 => \N__7022\,
            in2 => \_gnd_net_\,
            in3 => \N__6364\,
            lcout => \U712_CHIP_RAM.N_436\,
            ltout => \U712_CHIP_RAM.N_436_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__8294\,
            in1 => \_gnd_net_\,
            in2 => \N__5226\,
            in3 => \N__7109\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10656\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110111"
        )
    port map (
            in0 => \N__8455\,
            in1 => \N__6936\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_83\,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__5211\,
            in1 => \N__6486\,
            in2 => \N__5497\,
            in3 => \N__5214\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__10660\,
            ce => \N__5438\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__5210\,
            in1 => \N__7269\,
            in2 => \N__5498\,
            in3 => \N__5199\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \N__10660\,
            ce => \N__5438\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5486\,
            in1 => \N__6630\,
            in2 => \_gnd_net_\,
            in3 => \N__5196\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__10660\,
            ce => \N__5438\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5492\,
            in1 => \N__7030\,
            in2 => \_gnd_net_\,
            in3 => \N__5532\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__10660\,
            ce => \N__5438\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5487\,
            in1 => \N__5529\,
            in2 => \_gnd_net_\,
            in3 => \N__5517\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__10660\,
            ce => \N__5438\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5493\,
            in1 => \N__5514\,
            in2 => \_gnd_net_\,
            in3 => \N__5502\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__10660\,
            ce => \N__5438\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5488\,
            in1 => \N__5454\,
            in2 => \_gnd_net_\,
            in3 => \N__5457\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10660\,
            ce => \N__5438\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI94JE1_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7253\,
            in1 => \N__7020\,
            in2 => \N__6634\,
            in3 => \N__8448\,
            lcout => \U712_CHIP_RAM.N_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7388\,
            in1 => \N__5400\,
            in2 => \N__7166\,
            in3 => \N__5341\,
            lcout => \DMA_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10667\,
            ce => \N__5280\,
            sr => \N__11207\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7141\,
            in1 => \N__7387\,
            in2 => \_gnd_net_\,
            in3 => \N__7021\,
            lcout => \U712_CHIP_RAM.N_283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001010"
        )
    port map (
            in0 => \N__7254\,
            in1 => \N__6470\,
            in2 => \N__6939\,
            in3 => \N__6627\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_237_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIGRU43_1_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100001111"
        )
    port map (
            in0 => \N__6471\,
            in1 => \N__6919\,
            in2 => \N__5268\,
            in3 => \N__7140\,
            lcout => \U712_CHIP_RAM.N_281\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101110100101"
        )
    port map (
            in0 => \N__6472\,
            in1 => \N__6920\,
            in2 => \N__7165\,
            in3 => \N__7255\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_5_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5987\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__11198\
        );

    \U712_REG_SM.STATE_COUNTER_4_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5844\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__11198\
        );

    \U712_REG_SM.STATE_COUNTER_6_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5817\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__11198\
        );

    \U712_REG_SM.LDSn_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__5736\,
            in1 => \N__5811\,
            in2 => \N__5805\,
            in3 => \N__5774\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.LDSnC_net\,
            ce => 'H',
            sr => \N__11193\
        );

    \U712_REG_SM.UDSn_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__5751\,
            in1 => \N__5708\,
            in2 => \N__5745\,
            in3 => \N__5735\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.LDSnC_net\,
            ce => 'H',
            sr => \N__11193\
        );

    \U712_REG_SM.REG_CPU_CYCLE_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000100100001"
        )
    port map (
            in0 => \N__5986\,
            in1 => \N__5566\,
            in2 => \N__5934\,
            in3 => \N__5678\,
            lcout => \REG_CPU_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.LDSnC_net\,
            ce => 'H',
            sr => \N__11193\
        );

    \U712_REG_SM.REG_TACK_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__6051\,
            in1 => \N__6009\,
            in2 => \N__7662\,
            in3 => \N__5667\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.LDSnC_net\,
            ce => 'H',
            sr => \N__11193\
        );

    \U712_REG_SM.STATE_COUNTER_7_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__6119\,
            in1 => \N__5660\,
            in2 => \N__5568\,
            in3 => \N__5616\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.LDSnC_net\,
            ce => 'H',
            sr => \N__11193\
        );

    \U712_REG_SM.REG_WRITE_CYCLE_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110001011100"
        )
    port map (
            in0 => \N__6233\,
            in1 => \N__6044\,
            in2 => \N__6204\,
            in3 => \N__6141\,
            lcout => \REG_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.LDSnC_net\,
            ce => 'H',
            sr => \N__11193\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6120\,
            in1 => \N__6032\,
            in2 => \_gnd_net_\,
            in3 => \N__6098\,
            lcout => \U712_REG_SM.N_274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010011"
        )
    port map (
            in0 => \N__6033\,
            in1 => \N__6007\,
            in2 => \N__5991\,
            in3 => \N__5954\,
            lcout => \U712_REG_SM.REG_CPU_CYCLE_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6891\,
            in1 => \N__5910\,
            in2 => \_gnd_net_\,
            in3 => \N__6375\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNIK9021_0_3_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9454\,
            in1 => \N__9201\,
            in2 => \N__9407\,
            in3 => \N__9241\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__6938\,
            in1 => \N__6396\,
            in2 => \N__6491\,
            in3 => \N__6266\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__7437\,
            in1 => \N__6629\,
            in2 => \N__5913\,
            in3 => \N__5906\,
            lcout => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5874\,
            in1 => \N__5859\,
            in2 => \_gnd_net_\,
            in3 => \N__9362\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__7247\,
            in1 => \N__6334\,
            in2 => \N__6944\,
            in3 => \N__6625\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111011101110"
        )
    port map (
            in0 => \N__6390\,
            in1 => \N__6933\,
            in2 => \N__6347\,
            in3 => \N__7249\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIBKQ41_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__10811\,
            in1 => \N__7248\,
            in2 => \N__6346\,
            in3 => \N__6932\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CLK_EN_5_0_i_i_a2_0_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJIDU3_4_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7029\,
            in2 => \N__6378\,
            in3 => \N__6371\,
            lcout => \U712_CHIP_RAM.N_130\,
            ltout => \U712_CHIP_RAM.N_130_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__6626\,
            in1 => \N__6342\,
            in2 => \N__6285\,
            in3 => \N__10833\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_60_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__6282\,
            in1 => \N__8287\,
            in2 => \N__6276\,
            in3 => \N__7601\,
            lcout => \CPU_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_0_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7246\,
            in2 => \_gnd_net_\,
            in3 => \N__6928\,
            lcout => \U712_CHIP_RAM.N_248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001010"
        )
    port map (
            in0 => \N__6628\,
            in1 => \N__7019\,
            in2 => \N__6492\,
            in3 => \N__6273\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI52LA2_0_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__7267\,
            in1 => \N__6940\,
            in2 => \_gnd_net_\,
            in3 => \N__6267\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDs_0_6\,
            ltout => \U712_CHIP_RAM.SDRAM_CMDs_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__7742\,
            in1 => \N__7268\,
            in2 => \N__6642\,
            in3 => \N__6487\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__7775\,
            in1 => \N__7310\,
            in2 => \N__6639\,
            in3 => \N__9450\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10661\,
            ce => 'H',
            sr => \N__11199\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI0BPC1_4_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__7245\,
            in1 => \N__6617\,
            in2 => \_gnd_net_\,
            in3 => \N__7018\,
            lcout => \U712_CHIP_RAM.N_377\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_3_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6488\,
            in1 => \N__7292\,
            in2 => \_gnd_net_\,
            in3 => \N__7153\,
            lcout => \U712_CHIP_RAM.N_311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101111111"
        )
    port map (
            in0 => \N__6542\,
            in1 => \N__8261\,
            in2 => \N__7571\,
            in3 => \N__7708\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.TACK_STATE_r_sx_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__7604\,
            in1 => \N__7564\,
            in2 => \N__6501\,
            in3 => \N__7650\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10668\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIFCQ24_4_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__6489\,
            in1 => \N__6498\,
            in2 => \_gnd_net_\,
            in3 => \N__7042\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDs_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__7043\,
            in1 => \N__6490\,
            in2 => \N__6945\,
            in3 => \N__6417\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__7314\,
            in1 => \N__6411\,
            in2 => \N__9200\,
            in3 => \N__6405\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10672\,
            ce => 'H',
            sr => \N__11185\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__6740\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6924\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__6776\,
            in1 => \N__6813\,
            in2 => \_gnd_net_\,
            in3 => \N__6807\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10676\,
            ce => 'H',
            sr => \N__11179\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011011111111111"
        )
    port map (
            in0 => \N__7605\,
            in1 => \N__7713\,
            in2 => \N__7661\,
            in3 => \N__8208\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10679\,
            ce => \N__7902\,
            sr => \N__11178\
        );

    \CONSTANT_ONE_LUT4_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__9363\,
            in1 => \N__7443\,
            in2 => \N__9057\,
            in3 => \N__10795\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6717\,
            in1 => \N__10794\,
            in2 => \_gnd_net_\,
            in3 => \N__10497\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_292_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8769\,
            in2 => \N__6696\,
            in3 => \N__9364\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_207_i_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111110101"
        )
    port map (
            in0 => \N__8019\,
            in1 => \N__7893\,
            in2 => \N__8398\,
            in3 => \N__10796\,
            lcout => \N_207_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6681\,
            in1 => \N__6663\,
            in2 => \_gnd_net_\,
            in3 => \N__9338\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_205_i_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__7884\,
            in1 => \N__10862\,
            in2 => \N__8018\,
            in3 => \N__8375\,
            lcout => \N_205_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7476\,
            in1 => \N__7455\,
            in2 => \_gnd_net_\,
            in3 => \N__9337\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__9448\,
            in1 => \N__9336\,
            in2 => \_gnd_net_\,
            in3 => \N__9194\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN91M2_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__7741\,
            in1 => \N__7436\,
            in2 => \_gnd_net_\,
            in3 => \N__7160\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI8N6A9_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__7419\,
            in1 => \N__7404\,
            in2 => \N__7392\,
            in3 => \N__7389\,
            lcout => \U712_CHIP_RAM.N_50\,
            ltout => \U712_CHIP_RAM.N_50_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111100000"
        )
    port map (
            in0 => \N__7323\,
            in1 => \N__6951\,
            in2 => \N__7317\,
            in3 => \N__9358\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10658\,
            ce => 'H',
            sr => \N__11194\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_3_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11250\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7309\,
            lcout => \U712_CHIP_RAM.N_50_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__7293\,
            in1 => \N__7167\,
            in2 => \N__7044\,
            in3 => \N__6972\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_280_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6954\,
            in3 => \N__7757\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDsr_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8260\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7526\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8259\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7617\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNIK9021_3_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000111"
        )
    port map (
            in0 => \N__9449\,
            in1 => \N__9330\,
            in2 => \N__9240\,
            in3 => \N__9175\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8258\,
            in1 => \N__7829\,
            in2 => \_gnd_net_\,
            in3 => \N__7565\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10662\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_3_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7782\,
            in1 => \N__7776\,
            in2 => \N__7764\,
            in3 => \N__7746\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10669\,
            ce => \N__7725\,
            sr => \N__11180\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8265\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7712\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_252_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__7676\,
            in1 => \N__7602\,
            in2 => \N__7665\,
            in3 => \N__7654\,
            lcout => \U712_CYCLE_TERM.N_252_i_0_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7616\,
            in1 => \N__7603\,
            in2 => \N__7566\,
            in3 => \N__7525\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8322\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8242\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10673\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7929\,
            in2 => \_gnd_net_\,
            in3 => \N__8321\,
            lcout => \U712_CHIP_RAM.un3_DMA_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__8150\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7908\,
            lcout => \U712_CYCLE_TERM.N_252_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_i_o3_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011010101"
        )
    port map (
            in0 => \N__9797\,
            in1 => \N__9873\,
            in2 => \N__9713\,
            in3 => \N__9630\,
            lcout => \U712_BYTE_ENABLE.N_257\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_i_o3_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101101110101"
        )
    port map (
            in0 => \N__9798\,
            in1 => \N__9877\,
            in2 => \N__9714\,
            in3 => \N__9631\,
            lcout => \U712_BYTE_ENABLE.N_258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LMBE_i_o3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111111001"
        )
    port map (
            in0 => \N__9809\,
            in1 => \N__9632\,
            in2 => \N__9879\,
            in3 => \N__9699\,
            lcout => \U712_BYTE_ENABLE.N_259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8661\,
            in1 => \N__8130\,
            in2 => \_gnd_net_\,
            in3 => \N__7875\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10644\,
            ce => \N__10557\,
            sr => \N__11203\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8820\,
            in1 => \N__8697\,
            in2 => \N__8787\,
            in3 => \N__8523\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10644\,
            ce => \N__10557\,
            sr => \N__11203\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9463\,
            in2 => \_gnd_net_\,
            in3 => \N__9202\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011110000"
        )
    port map (
            in0 => \N__10804\,
            in1 => \N__9120\,
            in2 => \N__8133\,
            in3 => \N__9396\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8097\,
            in1 => \N__8025\,
            in2 => \_gnd_net_\,
            in3 => \N__8124\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10646\,
            ce => \N__10564\,
            sr => \N__11196\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110111011"
        )
    port map (
            in0 => \N__9981\,
            in1 => \N__10909\,
            in2 => \N__8052\,
            in3 => \N__10849\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_222_i_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111110101"
        )
    port map (
            in0 => \N__8415\,
            in1 => \N__8091\,
            in2 => \N__8399\,
            in3 => \N__10854\,
            lcout => \N_222_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__10853\,
            in1 => \N__8058\,
            in2 => \N__9387\,
            in3 => \N__9033\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__10908\,
            in1 => \N__8048\,
            in2 => \N__10867\,
            in3 => \N__9980\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0_0_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__11079\,
            in1 => \N__8469\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8001\,
            in1 => \N__7980\,
            in2 => \_gnd_net_\,
            in3 => \N__9333\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7965\,
            in1 => \N__7947\,
            in2 => \_gnd_net_\,
            in3 => \N__9332\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9334\,
            in1 => \N__8559\,
            in2 => \_gnd_net_\,
            in3 => \N__8541\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__10865\,
            in1 => \N__9042\,
            in2 => \N__8526\,
            in3 => \N__9335\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_ess_RNIAJSH1_3_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11249\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8514\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8508\,
            in1 => \N__8487\,
            in2 => \_gnd_net_\,
            in3 => \N__9331\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_0_0_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8472\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11043\,
            lcout => \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_0Z0Z_0\,
            ltout => \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_203_i_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__10866\,
            in1 => \N__8313\,
            in2 => \N__8406\,
            in3 => \N__8394\,
            lcout => \N_203_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__11042\,
            in1 => \N__11075\,
            in2 => \_gnd_net_\,
            in3 => \N__8241\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10664\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_i_o3_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100011111"
        )
    port map (
            in0 => \N__9878\,
            in1 => \N__9703\,
            in2 => \N__9636\,
            in3 => \N__9810\,
            lcout => \U712_BYTE_ENABLE.N_260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8212\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8816\,
            in1 => \N__8706\,
            in2 => \N__8788\,
            in3 => \N__8913\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10647\,
            ce => \N__10566\,
            sr => \N__11213\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__10843\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9391\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__8670\,
            in1 => \N__10844\,
            in2 => \N__9408\,
            in3 => \N__9093\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111011"
        )
    port map (
            in0 => \N__10842\,
            in1 => \N__9392\,
            in2 => \N__9119\,
            in3 => \N__8768\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8817\,
            in1 => \N__9126\,
            in2 => \N__8789\,
            in3 => \N__8655\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10650\,
            ce => \N__10565\,
            sr => \N__11200\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__10855\,
            in1 => \N__8628\,
            in2 => \N__9411\,
            in3 => \N__8904\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__8819\,
            in1 => \N__8783\,
            in2 => \N__8616\,
            in3 => \N__9099\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10650\,
            ce => \N__10565\,
            sr => \N__11200\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__8782\,
            in1 => \N__8818\,
            in2 => \N__10308\,
            in3 => \N__8565\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10650\,
            ce => \N__10565\,
            sr => \N__11200\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__9383\,
            in1 => \N__8571\,
            in2 => \N__9021\,
            in3 => \N__10864\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__10863\,
            in1 => \N__8919\,
            in2 => \N__9403\,
            in3 => \N__8925\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10283\,
            in1 => \N__10485\,
            in2 => \_gnd_net_\,
            in3 => \N__10133\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__9935\,
            sr => \N__11186\
        );

    \U712_CHIP_RAM.DMA_A20_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__10132\,
            in1 => \N__8895\,
            in2 => \N__10284\,
            in3 => \N__8864\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__11181\
        );

    \U712_BYTE_ENABLE.N_260_i_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001001000"
        )
    port map (
            in0 => \N__9806\,
            in1 => \N__9870\,
            in2 => \N__9629\,
            in3 => \N__9707\,
            lcout => \N_260_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_259_i_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111000100"
        )
    port map (
            in0 => \N__9869\,
            in1 => \N__9805\,
            in2 => \N__9715\,
            in3 => \N__9612\,
            lcout => \N_259_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8815\,
            in1 => \N__10362\,
            in2 => \N__8790\,
            in3 => \N__8730\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10651\,
            ce => \N__10570\,
            sr => \N__11214\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10103\,
            in1 => \N__9011\,
            in2 => \_gnd_net_\,
            in3 => \N__9084\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9969\,
            ce => \N__9941\,
            sr => \N__11208\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9012\,
            in1 => \N__8966\,
            in2 => \_gnd_net_\,
            in3 => \N__10104\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9969\,
            ce => \N__9941\,
            sr => \N__11208\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__8967\,
            in1 => \_gnd_net_\,
            in2 => \N__10129\,
            in3 => \N__10227\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9969\,
            ce => \N__9941\,
            sr => \N__11208\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9083\,
            in1 => \N__10434\,
            in2 => \_gnd_net_\,
            in3 => \N__10102\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9969\,
            ce => \N__9941\,
            sr => \N__11208\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10350\,
            in1 => \N__10484\,
            in2 => \_gnd_net_\,
            in3 => \N__10108\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9969\,
            ce => \N__9941\,
            sr => \N__11208\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9081\,
            in1 => \N__10069\,
            in2 => \_gnd_net_\,
            in3 => \N__10433\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9939\,
            sr => \N__11201\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9005\,
            in1 => \N__9082\,
            in2 => \_gnd_net_\,
            in3 => \N__10070\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9939\,
            sr => \N__11201\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10225\,
            in1 => \N__8965\,
            in2 => \_gnd_net_\,
            in3 => \N__10071\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9939\,
            sr => \N__11201\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10072\,
            in1 => \N__10226\,
            in2 => \_gnd_net_\,
            in3 => \N__10187\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9939\,
            sr => \N__11201\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10073\,
            in1 => \N__10345\,
            in2 => \_gnd_net_\,
            in3 => \N__10483\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9939\,
            sr => \N__11201\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8998\,
            in1 => \N__8956\,
            in2 => \_gnd_net_\,
            in3 => \N__10112\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__9938\,
            sr => \N__11195\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10389\,
            in1 => \N__10419\,
            in2 => \_gnd_net_\,
            in3 => \N__10110\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__9936\,
            sr => \N__11187\
        );

    \U712_BYTE_ENABLE.N_257_i_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101001100"
        )
    port map (
            in0 => \N__9871\,
            in1 => \N__9807\,
            in2 => \N__9722\,
            in3 => \N__9616\,
            lcout => \N_257_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_258_i_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001100"
        )
    port map (
            in0 => \N__9872\,
            in1 => \N__9808\,
            in2 => \N__9723\,
            in3 => \N__9617\,
            lcout => \N_258_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CRCSn_LC_15_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9255\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10645\,
            ce => 'H',
            sr => \N__11233\
        );

    \U712_CHIP_RAM.RASn_LC_15_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9474\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10648\,
            ce => 'H',
            sr => \N__11232\
        );

    \U712_CHIP_RAM.CASn_LC_15_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9410\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10649\,
            ce => 'H',
            sr => \N__11225\
        );

    \U712_CHIP_RAM.WEn_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9210\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10649\,
            ce => 'H',
            sr => \N__11225\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9470\,
            in1 => \N__9409\,
            in2 => \N__9254\,
            in3 => \N__9209\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10652\,
            ce => \N__10571\,
            sr => \N__11222\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__10916\,
            in1 => \N__10956\,
            in2 => \N__10872\,
            in3 => \N__10443\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10663\,
            ce => \N__10572\,
            sr => \N__11215\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__10236\,
            in1 => \N__10917\,
            in2 => \N__10893\,
            in3 => \N__10871\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10663\,
            ce => \N__10572\,
            sr => \N__11215\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10338\,
            in1 => \N__10186\,
            in2 => \_gnd_net_\,
            in3 => \N__10068\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__9942\,
            sr => \N__11209\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10273\,
            in1 => \N__10482\,
            in2 => \_gnd_net_\,
            in3 => \N__10111\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9966\,
            ce => \N__9940\,
            sr => \N__11202\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10429\,
            in1 => \N__10382\,
            in2 => \_gnd_net_\,
            in3 => \N__10109\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9964\,
            ce => \N__9937\,
            sr => \N__11188\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10346\,
            in1 => \N__10188\,
            in2 => \_gnd_net_\,
            in3 => \N__10131\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9968\,
            ce => \N__9944\,
            sr => \N__11218\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10296\,
            in1 => \N__10272\,
            in2 => \_gnd_net_\,
            in3 => \N__10113\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9965\,
            ce => \N__9943\,
            sr => \N__11210\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10224\,
            in1 => \N__10176\,
            in2 => \_gnd_net_\,
            in3 => \N__10130\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9967\,
            ce => \N__9945\,
            sr => \N__11223\
        );

    \U712_BUFFERS.un1_DRDENn_0_a3_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__11060\,
            in1 => \N__11030\,
            in2 => \_gnd_net_\,
            in3 => \N__11001\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Feb 8 2025 11:14:35

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U109_TOP" view "INTERFACE"

module U109_TOP (
    AD0,
    AD2,
    DLL,
    DUU,
    AD1,
    AD3,
    DLM,
    DUM,
    PCICYCLEn,
    ADLATCH,
    PCI_DIR,
    ALATCH);

    output [7:0] AD0;
    output [7:0] AD2;
    input [7:0] DLL;
    input [7:0] DUU;
    output [7:0] AD1;
    output [7:0] AD3;
    input [7:0] DLM;
    input [7:0] DUM;
    output PCICYCLEn;
    output ADLATCH;
    output PCI_DIR;
    output ALATCH;

    wire N__2211;
    wire N__2210;
    wire N__2209;
    wire N__2202;
    wire N__2201;
    wire N__2200;
    wire N__2193;
    wire N__2192;
    wire N__2191;
    wire N__2184;
    wire N__2183;
    wire N__2182;
    wire N__2175;
    wire N__2174;
    wire N__2173;
    wire N__2166;
    wire N__2165;
    wire N__2164;
    wire N__2157;
    wire N__2156;
    wire N__2155;
    wire N__2148;
    wire N__2147;
    wire N__2146;
    wire N__2139;
    wire N__2138;
    wire N__2137;
    wire N__2130;
    wire N__2129;
    wire N__2128;
    wire N__2121;
    wire N__2120;
    wire N__2119;
    wire N__2112;
    wire N__2111;
    wire N__2110;
    wire N__2103;
    wire N__2102;
    wire N__2101;
    wire N__2094;
    wire N__2093;
    wire N__2092;
    wire N__2085;
    wire N__2084;
    wire N__2083;
    wire N__2076;
    wire N__2075;
    wire N__2074;
    wire N__2067;
    wire N__2066;
    wire N__2065;
    wire N__2058;
    wire N__2057;
    wire N__2056;
    wire N__2049;
    wire N__2048;
    wire N__2047;
    wire N__2040;
    wire N__2039;
    wire N__2038;
    wire N__2031;
    wire N__2030;
    wire N__2029;
    wire N__2022;
    wire N__2021;
    wire N__2020;
    wire N__2013;
    wire N__2012;
    wire N__2011;
    wire N__2004;
    wire N__2003;
    wire N__2002;
    wire N__1995;
    wire N__1994;
    wire N__1993;
    wire N__1986;
    wire N__1985;
    wire N__1984;
    wire N__1977;
    wire N__1976;
    wire N__1975;
    wire N__1968;
    wire N__1967;
    wire N__1966;
    wire N__1959;
    wire N__1958;
    wire N__1957;
    wire N__1950;
    wire N__1949;
    wire N__1948;
    wire N__1941;
    wire N__1940;
    wire N__1939;
    wire N__1932;
    wire N__1931;
    wire N__1930;
    wire N__1923;
    wire N__1922;
    wire N__1921;
    wire N__1914;
    wire N__1913;
    wire N__1912;
    wire N__1905;
    wire N__1904;
    wire N__1903;
    wire N__1896;
    wire N__1895;
    wire N__1894;
    wire N__1887;
    wire N__1886;
    wire N__1885;
    wire N__1878;
    wire N__1877;
    wire N__1876;
    wire N__1869;
    wire N__1868;
    wire N__1867;
    wire N__1860;
    wire N__1859;
    wire N__1858;
    wire N__1851;
    wire N__1850;
    wire N__1849;
    wire N__1842;
    wire N__1841;
    wire N__1840;
    wire N__1833;
    wire N__1832;
    wire N__1831;
    wire N__1824;
    wire N__1823;
    wire N__1822;
    wire N__1815;
    wire N__1814;
    wire N__1813;
    wire N__1806;
    wire N__1805;
    wire N__1804;
    wire N__1797;
    wire N__1796;
    wire N__1795;
    wire N__1788;
    wire N__1787;
    wire N__1786;
    wire N__1779;
    wire N__1778;
    wire N__1777;
    wire N__1770;
    wire N__1769;
    wire N__1768;
    wire N__1761;
    wire N__1760;
    wire N__1759;
    wire N__1752;
    wire N__1751;
    wire N__1750;
    wire N__1743;
    wire N__1742;
    wire N__1741;
    wire N__1734;
    wire N__1733;
    wire N__1732;
    wire N__1725;
    wire N__1724;
    wire N__1723;
    wire N__1716;
    wire N__1715;
    wire N__1714;
    wire N__1707;
    wire N__1706;
    wire N__1705;
    wire N__1698;
    wire N__1697;
    wire N__1696;
    wire N__1689;
    wire N__1688;
    wire N__1687;
    wire N__1680;
    wire N__1679;
    wire N__1678;
    wire N__1671;
    wire N__1670;
    wire N__1669;
    wire N__1662;
    wire N__1661;
    wire N__1660;
    wire N__1653;
    wire N__1652;
    wire N__1651;
    wire N__1644;
    wire N__1643;
    wire N__1642;
    wire N__1635;
    wire N__1634;
    wire N__1633;
    wire N__1626;
    wire N__1625;
    wire N__1624;
    wire N__1617;
    wire N__1616;
    wire N__1615;
    wire N__1608;
    wire N__1607;
    wire N__1606;
    wire N__1589;
    wire N__1586;
    wire N__1583;
    wire N__1580;
    wire N__1577;
    wire N__1574;
    wire N__1571;
    wire N__1568;
    wire N__1565;
    wire N__1562;
    wire N__1559;
    wire N__1556;
    wire N__1553;
    wire N__1550;
    wire N__1547;
    wire N__1544;
    wire N__1541;
    wire N__1538;
    wire N__1535;
    wire N__1532;
    wire N__1529;
    wire N__1526;
    wire N__1523;
    wire N__1520;
    wire N__1517;
    wire N__1514;
    wire N__1511;
    wire N__1508;
    wire N__1505;
    wire N__1502;
    wire N__1499;
    wire N__1496;
    wire N__1493;
    wire N__1490;
    wire N__1487;
    wire N__1484;
    wire N__1481;
    wire N__1478;
    wire N__1475;
    wire N__1472;
    wire N__1469;
    wire N__1466;
    wire N__1463;
    wire N__1460;
    wire N__1457;
    wire N__1454;
    wire N__1451;
    wire N__1448;
    wire N__1445;
    wire N__1442;
    wire N__1439;
    wire N__1436;
    wire N__1433;
    wire N__1430;
    wire N__1427;
    wire N__1424;
    wire N__1421;
    wire N__1418;
    wire N__1415;
    wire N__1412;
    wire N__1409;
    wire N__1406;
    wire N__1403;
    wire N__1400;
    wire N__1397;
    wire N__1394;
    wire N__1391;
    wire N__1388;
    wire N__1385;
    wire N__1382;
    wire N__1379;
    wire N__1376;
    wire N__1373;
    wire N__1370;
    wire N__1367;
    wire N__1364;
    wire N__1361;
    wire N__1358;
    wire N__1355;
    wire N__1352;
    wire N__1349;
    wire N__1346;
    wire N__1343;
    wire N__1340;
    wire N__1337;
    wire N__1334;
    wire N__1331;
    wire N__1328;
    wire N__1325;
    wire N__1322;
    wire N__1319;
    wire N__1316;
    wire N__1313;
    wire N__1310;
    wire N__1307;
    wire N__1304;
    wire N__1301;
    wire N__1298;
    wire N__1295;
    wire N__1292;
    wire N__1289;
    wire N__1286;
    wire N__1283;
    wire N__1280;
    wire N__1277;
    wire N__1274;
    wire N__1271;
    wire N__1268;
    wire N__1265;
    wire N__1262;
    wire N__1259;
    wire N__1256;
    wire N__1253;
    wire N__1250;
    wire N__1247;
    wire N__1244;
    wire N__1241;
    wire N__1238;
    wire N__1235;
    wire N__1232;
    wire N__1229;
    wire N__1226;
    wire N__1223;
    wire N__1220;
    wire N__1217;
    wire N__1214;
    wire N__1211;
    wire N__1208;
    wire N__1205;
    wire N__1202;
    wire N__1199;
    wire N__1196;
    wire N__1193;
    wire N__1190;
    wire N__1187;
    wire N__1184;
    wire N__1181;
    wire N__1178;
    wire N__1175;
    wire N__1172;
    wire N__1169;
    wire N__1166;
    wire N__1163;
    wire N__1160;
    wire N__1157;
    wire N__1154;
    wire N__1151;
    wire N__1148;
    wire N__1145;
    wire N__1142;
    wire N__1139;
    wire N__1136;
    wire N__1133;
    wire N__1130;
    wire N__1127;
    wire N__1124;
    wire N__1121;
    wire N__1118;
    wire N__1115;
    wire N__1112;
    wire N__1109;
    wire N__1106;
    wire N__1103;
    wire N__1100;
    wire N__1097;
    wire N__1094;
    wire N__1091;
    wire N__1088;
    wire N__1085;
    wire N__1082;
    wire N__1079;
    wire N__1076;
    wire N__1073;
    wire N__1070;
    wire N__1067;
    wire N__1064;
    wire N__1061;
    wire N__1058;
    wire N__1055;
    wire N__1052;
    wire N__1049;
    wire N__1046;
    wire N__1043;
    wire N__1040;
    wire N__1037;
    wire N__1034;
    wire N__1031;
    wire N__1028;
    wire N__1025;
    wire N__1022;
    wire N__1019;
    wire N__1016;
    wire N__1013;
    wire N__1010;
    wire N__1007;
    wire N__1004;
    wire N__1001;
    wire N__998;
    wire N__995;
    wire N__992;
    wire N__989;
    wire N__986;
    wire N__983;
    wire N__980;
    wire N__977;
    wire N__974;
    wire N__971;
    wire N__968;
    wire N__965;
    wire N__962;
    wire N__959;
    wire N__956;
    wire N__953;
    wire N__950;
    wire N__947;
    wire N__944;
    wire N__941;
    wire N__938;
    wire N__935;
    wire N__932;
    wire N__929;
    wire N__926;
    wire N__923;
    wire N__920;
    wire N__917;
    wire N__914;
    wire N__911;
    wire N__908;
    wire N__905;
    wire N__902;
    wire N__899;
    wire N__896;
    wire N__893;
    wire N__890;
    wire N__887;
    wire N__884;
    wire N__881;
    wire N__878;
    wire N__875;
    wire N__872;
    wire N__869;
    wire N__866;
    wire N__863;
    wire N__860;
    wire N__857;
    wire N__854;
    wire N__851;
    wire N__848;
    wire N__845;
    wire N__842;
    wire N__839;
    wire N__836;
    wire N__833;
    wire N__830;
    wire N__827;
    wire N__824;
    wire N__821;
    wire N__818;
    wire N__815;
    wire N__812;
    wire N__809;
    wire N__806;
    wire N__803;
    wire N__800;
    wire AD0_c_2;
    wire AD3_c_0;
    wire VCCG0;
    wire AD1_c_6;
    wire AD3_c_6;
    wire AD2_c_3;
    wire AD0_c_3;
    wire AD1_c_0;
    wire AD3_c_4;
    wire AD2_c_4;
    wire AD2_c_5;
    wire AD3_c_3;
    wire AD0_c_1;
    wire GNDG0;
    wire AD1_c_2;
    wire AD2_c_6;
    wire AD0_c_4;
    wire AD1_c_5;
    wire AD2_c_7;
    wire AD3_c_1;
    wire AD1_c_3;
    wire AD0_c_7;
    wire AD2_c_0;
    wire AD3_c_5;
    wire AD0_c_6;
    wire AD1_c_7;
    wire AD3_c_7;
    wire AD2_c_1;
    wire AD0_c_5;
    wire AD2_c_2;
    wire AD1_c_4;
    wire AD0_c_0;
    wire AD1_c_1;
    wire AD3_c_2;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    IO_PAD AD3_obuf_2_iopad (
            .OE(N__2211),
            .DIN(N__2210),
            .DOUT(N__2209),
            .PACKAGEPIN(AD3[2]));
    defparam AD3_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam AD3_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO AD3_obuf_2_preio (
            .PADOEN(N__2211),
            .PADOUT(N__2210),
            .PADIN(N__2209),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1562),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUM_ibuf_1_iopad (
            .OE(N__2202),
            .DIN(N__2201),
            .DOUT(N__2200),
            .PACKAGEPIN(DUM[1]));
    defparam DUM_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DUM_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DUM_ibuf_1_preio (
            .PADOEN(N__2202),
            .PADOUT(N__2201),
            .PADIN(N__2200),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD1_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUU_ibuf_0_iopad (
            .OE(N__2193),
            .DIN(N__2192),
            .DOUT(N__2191),
            .PACKAGEPIN(DUU[0]));
    defparam DUU_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DUU_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DUU_ibuf_0_preio (
            .PADOEN(N__2193),
            .PADOUT(N__2192),
            .PADIN(N__2191),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD0_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD1_obuf_4_iopad (
            .OE(N__2184),
            .DIN(N__2183),
            .DOUT(N__2182),
            .PACKAGEPIN(AD1[4]));
    defparam AD1_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam AD1_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO AD1_obuf_4_preio (
            .PADOEN(N__2184),
            .PADOUT(N__2183),
            .PADIN(N__2182),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1313),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLM_ibuf_2_iopad (
            .OE(N__2175),
            .DIN(N__2174),
            .DOUT(N__2173),
            .PACKAGEPIN(DLM[2]));
    defparam DLM_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DLM_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DLM_ibuf_2_preio (
            .PADOEN(N__2175),
            .PADOUT(N__2174),
            .PADIN(N__2173),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD2_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD0_obuf_5_iopad (
            .OE(N__2166),
            .DIN(N__2165),
            .DOUT(N__2164),
            .PACKAGEPIN(AD0[5]));
    defparam AD0_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam AD0_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO AD0_obuf_5_preio (
            .PADOEN(N__2166),
            .PADOUT(N__2165),
            .PADIN(N__2164),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1364),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD2_obuf_1_iopad (
            .OE(N__2157),
            .DIN(N__2156),
            .DOUT(N__2155),
            .PACKAGEPIN(AD2[1]));
    defparam AD2_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam AD2_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO AD2_obuf_1_preio (
            .PADOEN(N__2157),
            .PADOUT(N__2156),
            .PADIN(N__2155),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1391),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLL_ibuf_7_iopad (
            .OE(N__2148),
            .DIN(N__2147),
            .DOUT(N__2146),
            .PACKAGEPIN(DLL[7]));
    defparam DLL_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DLL_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DLL_ibuf_7_preio (
            .PADOEN(N__2148),
            .PADOUT(N__2147),
            .PADIN(N__2146),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD3_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUM_ibuf_7_iopad (
            .OE(N__2139),
            .DIN(N__2138),
            .DOUT(N__2137),
            .PACKAGEPIN(DUM[7]));
    defparam DUM_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DUM_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DUM_ibuf_7_preio (
            .PADOEN(N__2139),
            .PADOUT(N__2138),
            .PADIN(N__2137),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD1_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUU_ibuf_6_iopad (
            .OE(N__2130),
            .DIN(N__2129),
            .DOUT(N__2128),
            .PACKAGEPIN(DUU[6]));
    defparam DUU_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DUU_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DUU_ibuf_6_preio (
            .PADOEN(N__2130),
            .PADOUT(N__2129),
            .PADIN(N__2128),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD0_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD3_obuf_5_iopad (
            .OE(N__2121),
            .DIN(N__2120),
            .DOUT(N__2119),
            .PACKAGEPIN(AD3[5]));
    defparam AD3_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam AD3_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO AD3_obuf_5_preio (
            .PADOEN(N__2121),
            .PADOUT(N__2120),
            .PADIN(N__2119),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1478),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLM_ibuf_0_iopad (
            .OE(N__2112),
            .DIN(N__2111),
            .DOUT(N__2110),
            .PACKAGEPIN(DLM[0]));
    defparam DLM_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DLM_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DLM_ibuf_0_preio (
            .PADOEN(N__2112),
            .PADOUT(N__2111),
            .PADIN(N__2110),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD2_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD0_obuf_7_iopad (
            .OE(N__2103),
            .DIN(N__2102),
            .DOUT(N__2101),
            .PACKAGEPIN(AD0[7]));
    defparam AD0_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam AD0_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO AD0_obuf_7_preio (
            .PADOEN(N__2103),
            .PADOUT(N__2102),
            .PADIN(N__2101),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1526),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD1_obuf_3_iopad (
            .OE(N__2094),
            .DIN(N__2093),
            .DOUT(N__2092),
            .PACKAGEPIN(AD1[3]));
    defparam AD1_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam AD1_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO AD1_obuf_3_preio (
            .PADOEN(N__2094),
            .PADOUT(N__2093),
            .PADIN(N__2092),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1121),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLL_ibuf_1_iopad (
            .OE(N__2085),
            .DIN(N__2084),
            .DOUT(N__2083),
            .PACKAGEPIN(DLL[1]));
    defparam DLL_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DLL_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DLL_ibuf_1_preio (
            .PADOEN(N__2085),
            .PADOUT(N__2084),
            .PADIN(N__2083),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD3_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLM_ibuf_7_iopad (
            .OE(N__2076),
            .DIN(N__2075),
            .DOUT(N__2074),
            .PACKAGEPIN(DLM[7]));
    defparam DLM_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DLM_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DLM_ibuf_7_preio (
            .PADOEN(N__2076),
            .PADOUT(N__2075),
            .PADIN(N__2074),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD2_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUM_ibuf_5_iopad (
            .OE(N__2067),
            .DIN(N__2066),
            .DOUT(N__2065),
            .PACKAGEPIN(DUM[5]));
    defparam DUM_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DUM_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DUM_ibuf_5_preio (
            .PADOEN(N__2067),
            .PADOUT(N__2066),
            .PADIN(N__2065),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD1_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUU_ibuf_4_iopad (
            .OE(N__2058),
            .DIN(N__2057),
            .DOUT(N__2056),
            .PACKAGEPIN(DUU[4]));
    defparam DUU_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DUU_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DUU_ibuf_4_preio (
            .PADOEN(N__2058),
            .PADOUT(N__2057),
            .PADIN(N__2056),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD0_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD2_obuf_6_iopad (
            .OE(N__2049),
            .DIN(N__2048),
            .DOUT(N__2047),
            .PACKAGEPIN(AD2[6]));
    defparam AD2_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam AD2_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO AD2_obuf_6_preio (
            .PADOEN(N__2049),
            .PADOUT(N__2048),
            .PADIN(N__2047),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1238),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD3_obuf_7_iopad (
            .OE(N__2040),
            .DIN(N__2039),
            .DOUT(N__2038),
            .PACKAGEPIN(AD3[7]));
    defparam AD3_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam AD3_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO AD3_obuf_7_preio (
            .PADOEN(N__2040),
            .PADOUT(N__2039),
            .PADIN(N__2038),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1412),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUM_ibuf_2_iopad (
            .OE(N__2031),
            .DIN(N__2030),
            .DOUT(N__2029),
            .PACKAGEPIN(DUM[2]));
    defparam DUM_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DUM_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DUM_ibuf_2_preio (
            .PADOEN(N__2031),
            .PADOUT(N__2030),
            .PADIN(N__2029),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD1_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PCI_DIR_obuf_iopad (
            .OE(N__2022),
            .DIN(N__2021),
            .DOUT(N__2020),
            .PACKAGEPIN(PCI_DIR));
    defparam PCI_DIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PCI_DIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PCI_DIR_obuf_preio (
            .PADOEN(N__2022),
            .PADOUT(N__2021),
            .PADIN(N__2020),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD0_obuf_1_iopad (
            .OE(N__2013),
            .DIN(N__2012),
            .DOUT(N__2011),
            .PACKAGEPIN(AD0[1]));
    defparam AD0_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam AD0_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO AD0_obuf_1_preio (
            .PADOEN(N__2013),
            .PADOUT(N__2012),
            .PADIN(N__2011),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__941),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD1_obuf_1_iopad (
            .OE(N__2004),
            .DIN(N__2003),
            .DOUT(N__2002),
            .PACKAGEPIN(AD1[1]));
    defparam AD1_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam AD1_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO AD1_obuf_1_preio (
            .PADOEN(N__2004),
            .PADOUT(N__2003),
            .PADIN(N__2002),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1589),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLL_ibuf_3_iopad (
            .OE(N__1995),
            .DIN(N__1994),
            .DOUT(N__1993),
            .PACKAGEPIN(DLL[3]));
    defparam DLL_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DLL_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DLL_ibuf_3_preio (
            .PADOEN(N__1995),
            .PADOUT(N__1994),
            .PADIN(N__1993),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD3_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLM_ibuf_5_iopad (
            .OE(N__1986),
            .DIN(N__1985),
            .DOUT(N__1984),
            .PACKAGEPIN(DLM[5]));
    defparam DLM_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DLM_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DLM_ibuf_5_preio (
            .PADOEN(N__1986),
            .PADOUT(N__1985),
            .PADIN(N__1984),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD2_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD2_obuf_4_iopad (
            .OE(N__1977),
            .DIN(N__1976),
            .DOUT(N__1975),
            .PACKAGEPIN(AD2[4]));
    defparam AD2_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam AD2_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO AD2_obuf_4_preio (
            .PADOEN(N__1977),
            .PADOUT(N__1976),
            .PADIN(N__1975),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1019),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD3_obuf_1_iopad (
            .OE(N__1968),
            .DIN(N__1967),
            .DOUT(N__1966),
            .PACKAGEPIN(AD3[1]));
    defparam AD3_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam AD3_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO AD3_obuf_1_preio (
            .PADOEN(N__1968),
            .PADOUT(N__1967),
            .PADIN(N__1966),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1145),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLL_ibuf_4_iopad (
            .OE(N__1959),
            .DIN(N__1958),
            .DOUT(N__1957),
            .PACKAGEPIN(DLL[4]));
    defparam DLL_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DLL_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DLL_ibuf_4_preio (
            .PADOEN(N__1959),
            .PADOUT(N__1958),
            .PADIN(N__1957),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD3_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUM_ibuf_0_iopad (
            .OE(N__1950),
            .DIN(N__1949),
            .DOUT(N__1948),
            .PACKAGEPIN(DUM[0]));
    defparam DUM_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DUM_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DUM_ibuf_0_preio (
            .PADOEN(N__1950),
            .PADOUT(N__1949),
            .PADIN(N__1948),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD1_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUU_ibuf_3_iopad (
            .OE(N__1941),
            .DIN(N__1940),
            .DOUT(N__1939),
            .PACKAGEPIN(DUU[3]));
    defparam DUU_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DUU_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DUU_ibuf_3_preio (
            .PADOEN(N__1941),
            .PADOUT(N__1940),
            .PADIN(N__1939),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD0_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD0_obuf_3_iopad (
            .OE(N__1932),
            .DIN(N__1931),
            .DOUT(N__1930),
            .PACKAGEPIN(AD0[3]));
    defparam AD0_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam AD0_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO AD0_obuf_3_preio (
            .PADOEN(N__1932),
            .PADOUT(N__1931),
            .PADIN(N__1930),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1094),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD1_obuf_7_iopad (
            .OE(N__1923),
            .DIN(N__1922),
            .DOUT(N__1921),
            .PACKAGEPIN(AD1[7]));
    defparam AD1_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam AD1_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO AD1_obuf_7_preio (
            .PADOEN(N__1923),
            .PADOUT(N__1922),
            .PADIN(N__1921),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1427),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLM_ibuf_3_iopad (
            .OE(N__1914),
            .DIN(N__1913),
            .DOUT(N__1912),
            .PACKAGEPIN(DLM[3]));
    defparam DLM_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DLM_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DLM_ibuf_3_preio (
            .PADOEN(N__1914),
            .PADOUT(N__1913),
            .PADIN(N__1912),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD2_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD2_obuf_2_iopad (
            .OE(N__1905),
            .DIN(N__1904),
            .DOUT(N__1903),
            .PACKAGEPIN(AD2[2]));
    defparam AD2_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam AD2_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO AD2_obuf_2_preio (
            .PADOEN(N__1905),
            .PADOUT(N__1904),
            .PADIN(N__1903),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1340),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD3_obuf_3_iopad (
            .OE(N__1896),
            .DIN(N__1895),
            .DOUT(N__1894),
            .PACKAGEPIN(AD3[3]));
    defparam AD3_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam AD3_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO AD3_obuf_3_preio (
            .PADOEN(N__1896),
            .PADOUT(N__1895),
            .PADIN(N__1894),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__968),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLL_ibuf_6_iopad (
            .OE(N__1887),
            .DIN(N__1886),
            .DOUT(N__1885),
            .PACKAGEPIN(DLL[6]));
    defparam DLL_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DLL_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DLL_ibuf_6_preio (
            .PADOEN(N__1887),
            .PADOUT(N__1886),
            .PADIN(N__1885),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD3_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUM_ibuf_6_iopad (
            .OE(N__1878),
            .DIN(N__1877),
            .DOUT(N__1876),
            .PACKAGEPIN(DUM[6]));
    defparam DUM_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DUM_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DUM_ibuf_6_preio (
            .PADOEN(N__1878),
            .PADOUT(N__1877),
            .PADIN(N__1876),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD1_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUU_ibuf_1_iopad (
            .OE(N__1869),
            .DIN(N__1868),
            .DOUT(N__1867),
            .PACKAGEPIN(DUU[1]));
    defparam DUU_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DUU_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DUU_ibuf_1_preio (
            .PADOEN(N__1869),
            .PADOUT(N__1868),
            .PADIN(N__1867),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD0_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD1_obuf_5_iopad (
            .OE(N__1860),
            .DIN(N__1859),
            .DOUT(N__1858),
            .PACKAGEPIN(AD1[5]));
    defparam AD1_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam AD1_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO AD1_obuf_5_preio (
            .PADOEN(N__1860),
            .PADOUT(N__1859),
            .PADIN(N__1858),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1190),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD3_obuf_4_iopad (
            .OE(N__1851),
            .DIN(N__1850),
            .DOUT(N__1849),
            .PACKAGEPIN(AD3[4]));
    defparam AD3_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam AD3_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO AD3_obuf_4_preio (
            .PADOEN(N__1851),
            .PADOUT(N__1850),
            .PADIN(N__1849),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1049),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ADLATCH_obuf_iopad (
            .OE(N__1842),
            .DIN(N__1841),
            .DOUT(N__1840),
            .PACKAGEPIN(ADLATCH));
    defparam ADLATCH_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ADLATCH_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ADLATCH_obuf_preio (
            .PADOEN(N__1842),
            .PADOUT(N__1841),
            .PADIN(N__1840),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLM_ibuf_1_iopad (
            .OE(N__1833),
            .DIN(N__1832),
            .DOUT(N__1831),
            .PACKAGEPIN(DLM[1]));
    defparam DLM_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DLM_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DLM_ibuf_1_preio (
            .PADOEN(N__1833),
            .PADOUT(N__1832),
            .PADIN(N__1831),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD2_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD0_obuf_4_iopad (
            .OE(N__1824),
            .DIN(N__1823),
            .DOUT(N__1822),
            .PACKAGEPIN(AD0[4]));
    defparam AD0_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam AD0_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO AD0_obuf_4_preio (
            .PADOEN(N__1824),
            .PADOUT(N__1823),
            .PADIN(N__1822),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1214),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD1_obuf_2_iopad (
            .OE(N__1815),
            .DIN(N__1814),
            .DOUT(N__1813),
            .PACKAGEPIN(AD1[2]));
    defparam AD1_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam AD1_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO AD1_obuf_2_preio (
            .PADOEN(N__1815),
            .PADOUT(N__1814),
            .PADIN(N__1813),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1265),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD2_obuf_0_iopad (
            .OE(N__1806),
            .DIN(N__1805),
            .DOUT(N__1804),
            .PACKAGEPIN(AD2[0]));
    defparam AD2_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam AD2_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO AD2_obuf_0_preio (
            .PADOEN(N__1806),
            .PADOUT(N__1805),
            .PADIN(N__1804),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1499),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ALATCH_obuf_iopad (
            .OE(N__1797),
            .DIN(N__1796),
            .DOUT(N__1795),
            .PACKAGEPIN(ALATCH));
    defparam ALATCH_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ALATCH_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ALATCH_obuf_preio (
            .PADOEN(N__1797),
            .PADOUT(N__1796),
            .PADIN(N__1795),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLL_ibuf_0_iopad (
            .OE(N__1788),
            .DIN(N__1787),
            .DOUT(N__1786),
            .PACKAGEPIN(DLL[0]));
    defparam DLL_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DLL_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DLL_ibuf_0_preio (
            .PADOEN(N__1788),
            .PADOUT(N__1787),
            .PADIN(N__1786),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD3_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUM_ibuf_4_iopad (
            .OE(N__1779),
            .DIN(N__1778),
            .DOUT(N__1777),
            .PACKAGEPIN(DUM[4]));
    defparam DUM_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DUM_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DUM_ibuf_4_preio (
            .PADOEN(N__1779),
            .PADOUT(N__1778),
            .PADIN(N__1777),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD1_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUU_ibuf_7_iopad (
            .OE(N__1770),
            .DIN(N__1769),
            .DOUT(N__1768),
            .PACKAGEPIN(DUU[7]));
    defparam DUU_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DUU_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DUU_ibuf_7_preio (
            .PADOEN(N__1770),
            .PADOUT(N__1769),
            .PADIN(N__1768),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD0_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD2_obuf_7_iopad (
            .OE(N__1761),
            .DIN(N__1760),
            .DOUT(N__1759),
            .PACKAGEPIN(AD2[7]));
    defparam AD2_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam AD2_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO AD2_obuf_7_preio (
            .PADOEN(N__1761),
            .PADOUT(N__1760),
            .PADIN(N__1759),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1169),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD3_obuf_6_iopad (
            .OE(N__1752),
            .DIN(N__1751),
            .DOUT(N__1750),
            .PACKAGEPIN(AD3[6]));
    defparam AD3_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam AD3_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO AD3_obuf_6_preio (
            .PADOEN(N__1752),
            .PADOUT(N__1751),
            .PADIN(N__1750),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__893),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD0_obuf_6_iopad (
            .OE(N__1743),
            .DIN(N__1742),
            .DOUT(N__1741),
            .PACKAGEPIN(AD0[6]));
    defparam AD0_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam AD0_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO AD0_obuf_6_preio (
            .PADOEN(N__1743),
            .PADOUT(N__1742),
            .PADIN(N__1741),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1448),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD1_obuf_0_iopad (
            .OE(N__1734),
            .DIN(N__1733),
            .DOUT(N__1732),
            .PACKAGEPIN(AD1[0]));
    defparam AD1_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam AD1_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO AD1_obuf_0_preio (
            .PADOEN(N__1734),
            .PADOUT(N__1733),
            .PADIN(N__1732),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1076),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLL_ibuf_2_iopad (
            .OE(N__1725),
            .DIN(N__1724),
            .DOUT(N__1723),
            .PACKAGEPIN(DLL[2]));
    defparam DLL_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DLL_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DLL_ibuf_2_preio (
            .PADOEN(N__1725),
            .PADOUT(N__1724),
            .PADIN(N__1723),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD3_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLM_ibuf_6_iopad (
            .OE(N__1716),
            .DIN(N__1715),
            .DOUT(N__1714),
            .PACKAGEPIN(DLM[6]));
    defparam DLM_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DLM_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DLM_ibuf_6_preio (
            .PADOEN(N__1716),
            .PADOUT(N__1715),
            .PADIN(N__1714),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD2_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUU_ibuf_5_iopad (
            .OE(N__1707),
            .DIN(N__1706),
            .DOUT(N__1705),
            .PACKAGEPIN(DUU[5]));
    defparam DUU_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DUU_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DUU_ibuf_5_preio (
            .PADOEN(N__1707),
            .PADOUT(N__1706),
            .PADIN(N__1705),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD0_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD2_obuf_5_iopad (
            .OE(N__1698),
            .DIN(N__1697),
            .DOUT(N__1696),
            .PACKAGEPIN(AD2[5]));
    defparam AD2_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam AD2_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO AD2_obuf_5_preio (
            .PADOEN(N__1698),
            .PADOUT(N__1697),
            .PADIN(N__1696),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__995),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD3_obuf_0_iopad (
            .OE(N__1689),
            .DIN(N__1688),
            .DOUT(N__1687),
            .PACKAGEPIN(AD3[0]));
    defparam AD3_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam AD3_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO AD3_obuf_0_preio (
            .PADOEN(N__1689),
            .PADOUT(N__1688),
            .PADIN(N__1687),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__845),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUM_ibuf_3_iopad (
            .OE(N__1680),
            .DIN(N__1679),
            .DOUT(N__1678),
            .PACKAGEPIN(DUM[3]));
    defparam DUM_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DUM_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DUM_ibuf_3_preio (
            .PADOEN(N__1680),
            .PADOUT(N__1679),
            .PADIN(N__1678),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD1_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DUU_ibuf_2_iopad (
            .OE(N__1671),
            .DIN(N__1670),
            .DOUT(N__1669),
            .PACKAGEPIN(DUU[2]));
    defparam DUU_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DUU_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DUU_ibuf_2_preio (
            .PADOEN(N__1671),
            .PADOUT(N__1670),
            .PADIN(N__1669),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD0_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PCICYCLEn_obuf_iopad (
            .OE(N__1662),
            .DIN(N__1661),
            .DOUT(N__1660),
            .PACKAGEPIN(PCICYCLEn));
    defparam PCICYCLEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PCICYCLEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PCICYCLEn_obuf_preio (
            .PADOEN(N__1662),
            .PADOUT(N__1661),
            .PADIN(N__1660),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1538),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD0_obuf_0_iopad (
            .OE(N__1653),
            .DIN(N__1652),
            .DOUT(N__1651),
            .PACKAGEPIN(AD0[0]));
    defparam AD0_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam AD0_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO AD0_obuf_0_preio (
            .PADOEN(N__1653),
            .PADOUT(N__1652),
            .PADIN(N__1651),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1292),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD1_obuf_6_iopad (
            .OE(N__1644),
            .DIN(N__1643),
            .DOUT(N__1642),
            .PACKAGEPIN(AD1[6]));
    defparam AD1_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam AD1_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO AD1_obuf_6_preio (
            .PADOEN(N__1644),
            .PADOUT(N__1643),
            .PADIN(N__1642),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__914),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLM_ibuf_4_iopad (
            .OE(N__1635),
            .DIN(N__1634),
            .DOUT(N__1633),
            .PACKAGEPIN(DLM[4]));
    defparam DLM_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DLM_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DLM_ibuf_4_preio (
            .PADOEN(N__1635),
            .PADOUT(N__1634),
            .PADIN(N__1633),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD2_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD2_obuf_3_iopad (
            .OE(N__1626),
            .DIN(N__1625),
            .DOUT(N__1624),
            .PACKAGEPIN(AD2[3]));
    defparam AD2_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam AD2_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO AD2_obuf_3_preio (
            .PADOEN(N__1626),
            .PADOUT(N__1625),
            .PADIN(N__1624),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__863),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DLL_ibuf_5_iopad (
            .OE(N__1617),
            .DIN(N__1616),
            .DOUT(N__1615),
            .PACKAGEPIN(DLL[5]));
    defparam DLL_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DLL_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DLL_ibuf_5_preio (
            .PADOEN(N__1617),
            .PADOUT(N__1616),
            .PADIN(N__1615),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AD3_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AD0_obuf_2_iopad (
            .OE(N__1608),
            .DIN(N__1607),
            .DOUT(N__1606),
            .PACKAGEPIN(AD0[2]));
    defparam AD0_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam AD0_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO AD0_obuf_2_preio (
            .PADOEN(N__1608),
            .PADOUT(N__1607),
            .PADIN(N__1606),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__821),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__335 (
            .O(N__1589),
            .I(N__1586));
    LocalMux I__334 (
            .O(N__1586),
            .I(N__1583));
    Span4Mux_s1_v I__333 (
            .O(N__1583),
            .I(N__1580));
    Span4Mux_v I__332 (
            .O(N__1580),
            .I(N__1577));
    Sp12to4 I__331 (
            .O(N__1577),
            .I(N__1574));
    Span12Mux_h I__330 (
            .O(N__1574),
            .I(N__1571));
    Span12Mux_v I__329 (
            .O(N__1571),
            .I(N__1568));
    Span12Mux_h I__328 (
            .O(N__1568),
            .I(N__1565));
    Odrv12 I__327 (
            .O(N__1565),
            .I(AD1_c_1));
    IoInMux I__326 (
            .O(N__1562),
            .I(N__1559));
    LocalMux I__325 (
            .O(N__1559),
            .I(N__1556));
    IoSpan4Mux I__324 (
            .O(N__1556),
            .I(N__1553));
    Span4Mux_s3_h I__323 (
            .O(N__1553),
            .I(N__1550));
    Sp12to4 I__322 (
            .O(N__1550),
            .I(N__1547));
    Span12Mux_v I__321 (
            .O(N__1547),
            .I(N__1544));
    Span12Mux_v I__320 (
            .O(N__1544),
            .I(N__1541));
    Odrv12 I__319 (
            .O(N__1541),
            .I(AD3_c_2));
    IoInMux I__318 (
            .O(N__1538),
            .I(N__1535));
    LocalMux I__317 (
            .O(N__1535),
            .I(N__1532));
    Span4Mux_s3_h I__316 (
            .O(N__1532),
            .I(N__1529));
    Odrv4 I__315 (
            .O(N__1529),
            .I(CONSTANT_ONE_NET));
    IoInMux I__314 (
            .O(N__1526),
            .I(N__1523));
    LocalMux I__313 (
            .O(N__1523),
            .I(N__1520));
    IoSpan4Mux I__312 (
            .O(N__1520),
            .I(N__1517));
    Span4Mux_s2_v I__311 (
            .O(N__1517),
            .I(N__1514));
    Span4Mux_v I__310 (
            .O(N__1514),
            .I(N__1511));
    Sp12to4 I__309 (
            .O(N__1511),
            .I(N__1508));
    Span12Mux_v I__308 (
            .O(N__1508),
            .I(N__1505));
    Span12Mux_v I__307 (
            .O(N__1505),
            .I(N__1502));
    Odrv12 I__306 (
            .O(N__1502),
            .I(AD0_c_7));
    IoInMux I__305 (
            .O(N__1499),
            .I(N__1496));
    LocalMux I__304 (
            .O(N__1496),
            .I(N__1493));
    Span12Mux_s4_v I__303 (
            .O(N__1493),
            .I(N__1490));
    Span12Mux_h I__302 (
            .O(N__1490),
            .I(N__1487));
    Span12Mux_v I__301 (
            .O(N__1487),
            .I(N__1484));
    Span12Mux_v I__300 (
            .O(N__1484),
            .I(N__1481));
    Odrv12 I__299 (
            .O(N__1481),
            .I(AD2_c_0));
    IoInMux I__298 (
            .O(N__1478),
            .I(N__1475));
    LocalMux I__297 (
            .O(N__1475),
            .I(N__1472));
    IoSpan4Mux I__296 (
            .O(N__1472),
            .I(N__1469));
    Span4Mux_s3_h I__295 (
            .O(N__1469),
            .I(N__1466));
    Sp12to4 I__294 (
            .O(N__1466),
            .I(N__1463));
    Span12Mux_v I__293 (
            .O(N__1463),
            .I(N__1460));
    Span12Mux_v I__292 (
            .O(N__1460),
            .I(N__1457));
    Span12Mux_h I__291 (
            .O(N__1457),
            .I(N__1454));
    Span12Mux_h I__290 (
            .O(N__1454),
            .I(N__1451));
    Odrv12 I__289 (
            .O(N__1451),
            .I(AD3_c_5));
    IoInMux I__288 (
            .O(N__1448),
            .I(N__1445));
    LocalMux I__287 (
            .O(N__1445),
            .I(N__1442));
    Span4Mux_s2_v I__286 (
            .O(N__1442),
            .I(N__1439));
    Sp12to4 I__285 (
            .O(N__1439),
            .I(N__1436));
    Span12Mux_h I__284 (
            .O(N__1436),
            .I(N__1433));
    Span12Mux_h I__283 (
            .O(N__1433),
            .I(N__1430));
    Odrv12 I__282 (
            .O(N__1430),
            .I(AD0_c_6));
    IoInMux I__281 (
            .O(N__1427),
            .I(N__1424));
    LocalMux I__280 (
            .O(N__1424),
            .I(N__1421));
    Span12Mux_s11_v I__279 (
            .O(N__1421),
            .I(N__1418));
    Span12Mux_h I__278 (
            .O(N__1418),
            .I(N__1415));
    Odrv12 I__277 (
            .O(N__1415),
            .I(AD1_c_7));
    IoInMux I__276 (
            .O(N__1412),
            .I(N__1409));
    LocalMux I__275 (
            .O(N__1409),
            .I(N__1406));
    Span12Mux_s9_h I__274 (
            .O(N__1406),
            .I(N__1403));
    Span12Mux_v I__273 (
            .O(N__1403),
            .I(N__1400));
    Span12Mux_v I__272 (
            .O(N__1400),
            .I(N__1397));
    Span12Mux_h I__271 (
            .O(N__1397),
            .I(N__1394));
    Odrv12 I__270 (
            .O(N__1394),
            .I(AD3_c_7));
    IoInMux I__269 (
            .O(N__1391),
            .I(N__1388));
    LocalMux I__268 (
            .O(N__1388),
            .I(N__1385));
    IoSpan4Mux I__267 (
            .O(N__1385),
            .I(N__1382));
    Span4Mux_s2_v I__266 (
            .O(N__1382),
            .I(N__1379));
    Span4Mux_v I__265 (
            .O(N__1379),
            .I(N__1376));
    Sp12to4 I__264 (
            .O(N__1376),
            .I(N__1373));
    Span12Mux_v I__263 (
            .O(N__1373),
            .I(N__1370));
    Span12Mux_v I__262 (
            .O(N__1370),
            .I(N__1367));
    Odrv12 I__261 (
            .O(N__1367),
            .I(AD2_c_1));
    IoInMux I__260 (
            .O(N__1364),
            .I(N__1361));
    LocalMux I__259 (
            .O(N__1361),
            .I(N__1358));
    IoSpan4Mux I__258 (
            .O(N__1358),
            .I(N__1355));
    Span4Mux_s2_v I__257 (
            .O(N__1355),
            .I(N__1352));
    Sp12to4 I__256 (
            .O(N__1352),
            .I(N__1349));
    Span12Mux_h I__255 (
            .O(N__1349),
            .I(N__1346));
    Span12Mux_h I__254 (
            .O(N__1346),
            .I(N__1343));
    Odrv12 I__253 (
            .O(N__1343),
            .I(AD0_c_5));
    IoInMux I__252 (
            .O(N__1340),
            .I(N__1337));
    LocalMux I__251 (
            .O(N__1337),
            .I(N__1334));
    IoSpan4Mux I__250 (
            .O(N__1334),
            .I(N__1331));
    Span4Mux_s1_v I__249 (
            .O(N__1331),
            .I(N__1328));
    Span4Mux_v I__248 (
            .O(N__1328),
            .I(N__1325));
    Sp12to4 I__247 (
            .O(N__1325),
            .I(N__1322));
    Span12Mux_v I__246 (
            .O(N__1322),
            .I(N__1319));
    Span12Mux_v I__245 (
            .O(N__1319),
            .I(N__1316));
    Odrv12 I__244 (
            .O(N__1316),
            .I(AD2_c_2));
    IoInMux I__243 (
            .O(N__1313),
            .I(N__1310));
    LocalMux I__242 (
            .O(N__1310),
            .I(N__1307));
    Span12Mux_s3_v I__241 (
            .O(N__1307),
            .I(N__1304));
    Span12Mux_v I__240 (
            .O(N__1304),
            .I(N__1301));
    Span12Mux_h I__239 (
            .O(N__1301),
            .I(N__1298));
    Span12Mux_h I__238 (
            .O(N__1298),
            .I(N__1295));
    Odrv12 I__237 (
            .O(N__1295),
            .I(AD1_c_4));
    IoInMux I__236 (
            .O(N__1292),
            .I(N__1289));
    LocalMux I__235 (
            .O(N__1289),
            .I(N__1286));
    IoSpan4Mux I__234 (
            .O(N__1286),
            .I(N__1283));
    Span4Mux_s1_h I__233 (
            .O(N__1283),
            .I(N__1280));
    Sp12to4 I__232 (
            .O(N__1280),
            .I(N__1277));
    Span12Mux_s11_v I__231 (
            .O(N__1277),
            .I(N__1274));
    Span12Mux_h I__230 (
            .O(N__1274),
            .I(N__1271));
    Span12Mux_h I__229 (
            .O(N__1271),
            .I(N__1268));
    Odrv12 I__228 (
            .O(N__1268),
            .I(AD0_c_0));
    IoInMux I__227 (
            .O(N__1265),
            .I(N__1262));
    LocalMux I__226 (
            .O(N__1262),
            .I(N__1259));
    Span4Mux_s0_v I__225 (
            .O(N__1259),
            .I(N__1256));
    Span4Mux_v I__224 (
            .O(N__1256),
            .I(N__1253));
    Sp12to4 I__223 (
            .O(N__1253),
            .I(N__1250));
    Span12Mux_h I__222 (
            .O(N__1250),
            .I(N__1247));
    Span12Mux_v I__221 (
            .O(N__1247),
            .I(N__1244));
    Span12Mux_h I__220 (
            .O(N__1244),
            .I(N__1241));
    Odrv12 I__219 (
            .O(N__1241),
            .I(AD1_c_2));
    IoInMux I__218 (
            .O(N__1238),
            .I(N__1235));
    LocalMux I__217 (
            .O(N__1235),
            .I(N__1232));
    IoSpan4Mux I__216 (
            .O(N__1232),
            .I(N__1229));
    Span4Mux_s2_v I__215 (
            .O(N__1229),
            .I(N__1226));
    Sp12to4 I__214 (
            .O(N__1226),
            .I(N__1223));
    Span12Mux_s10_v I__213 (
            .O(N__1223),
            .I(N__1220));
    Span12Mux_v I__212 (
            .O(N__1220),
            .I(N__1217));
    Odrv12 I__211 (
            .O(N__1217),
            .I(AD2_c_6));
    IoInMux I__210 (
            .O(N__1214),
            .I(N__1211));
    LocalMux I__209 (
            .O(N__1211),
            .I(N__1208));
    IoSpan4Mux I__208 (
            .O(N__1208),
            .I(N__1205));
    Span4Mux_s3_v I__207 (
            .O(N__1205),
            .I(N__1202));
    Sp12to4 I__206 (
            .O(N__1202),
            .I(N__1199));
    Span12Mux_h I__205 (
            .O(N__1199),
            .I(N__1196));
    Span12Mux_h I__204 (
            .O(N__1196),
            .I(N__1193));
    Odrv12 I__203 (
            .O(N__1193),
            .I(AD0_c_4));
    IoInMux I__202 (
            .O(N__1190),
            .I(N__1187));
    LocalMux I__201 (
            .O(N__1187),
            .I(N__1184));
    Span4Mux_s1_v I__200 (
            .O(N__1184),
            .I(N__1181));
    Sp12to4 I__199 (
            .O(N__1181),
            .I(N__1178));
    Span12Mux_h I__198 (
            .O(N__1178),
            .I(N__1175));
    Span12Mux_v I__197 (
            .O(N__1175),
            .I(N__1172));
    Odrv12 I__196 (
            .O(N__1172),
            .I(AD1_c_5));
    IoInMux I__195 (
            .O(N__1169),
            .I(N__1166));
    LocalMux I__194 (
            .O(N__1166),
            .I(N__1163));
    Span4Mux_s3_v I__193 (
            .O(N__1163),
            .I(N__1160));
    IoSpan4Mux I__192 (
            .O(N__1160),
            .I(N__1157));
    IoSpan4Mux I__191 (
            .O(N__1157),
            .I(N__1154));
    IoSpan4Mux I__190 (
            .O(N__1154),
            .I(N__1151));
    IoSpan4Mux I__189 (
            .O(N__1151),
            .I(N__1148));
    Odrv4 I__188 (
            .O(N__1148),
            .I(AD2_c_7));
    IoInMux I__187 (
            .O(N__1145),
            .I(N__1142));
    LocalMux I__186 (
            .O(N__1142),
            .I(N__1139));
    Span4Mux_s3_v I__185 (
            .O(N__1139),
            .I(N__1136));
    Sp12to4 I__184 (
            .O(N__1136),
            .I(N__1133));
    Span12Mux_s3_h I__183 (
            .O(N__1133),
            .I(N__1130));
    Span12Mux_v I__182 (
            .O(N__1130),
            .I(N__1127));
    Span12Mux_v I__181 (
            .O(N__1127),
            .I(N__1124));
    Odrv12 I__180 (
            .O(N__1124),
            .I(AD3_c_1));
    IoInMux I__179 (
            .O(N__1121),
            .I(N__1118));
    LocalMux I__178 (
            .O(N__1118),
            .I(N__1115));
    IoSpan4Mux I__177 (
            .O(N__1115),
            .I(N__1112));
    Span4Mux_s2_v I__176 (
            .O(N__1112),
            .I(N__1109));
    Span4Mux_v I__175 (
            .O(N__1109),
            .I(N__1106));
    Sp12to4 I__174 (
            .O(N__1106),
            .I(N__1103));
    Span12Mux_v I__173 (
            .O(N__1103),
            .I(N__1100));
    Span12Mux_h I__172 (
            .O(N__1100),
            .I(N__1097));
    Odrv12 I__171 (
            .O(N__1097),
            .I(AD1_c_3));
    IoInMux I__170 (
            .O(N__1094),
            .I(N__1091));
    LocalMux I__169 (
            .O(N__1091),
            .I(N__1088));
    Span12Mux_s4_v I__168 (
            .O(N__1088),
            .I(N__1085));
    Span12Mux_h I__167 (
            .O(N__1085),
            .I(N__1082));
    Span12Mux_h I__166 (
            .O(N__1082),
            .I(N__1079));
    Odrv12 I__165 (
            .O(N__1079),
            .I(AD0_c_3));
    IoInMux I__164 (
            .O(N__1076),
            .I(N__1073));
    LocalMux I__163 (
            .O(N__1073),
            .I(N__1070));
    IoSpan4Mux I__162 (
            .O(N__1070),
            .I(N__1067));
    Span4Mux_s3_h I__161 (
            .O(N__1067),
            .I(N__1064));
    Sp12to4 I__160 (
            .O(N__1064),
            .I(N__1061));
    Span12Mux_v I__159 (
            .O(N__1061),
            .I(N__1058));
    Span12Mux_h I__158 (
            .O(N__1058),
            .I(N__1055));
    Span12Mux_h I__157 (
            .O(N__1055),
            .I(N__1052));
    Odrv12 I__156 (
            .O(N__1052),
            .I(AD1_c_0));
    IoInMux I__155 (
            .O(N__1049),
            .I(N__1046));
    LocalMux I__154 (
            .O(N__1046),
            .I(N__1043));
    IoSpan4Mux I__153 (
            .O(N__1043),
            .I(N__1040));
    Span4Mux_s2_h I__152 (
            .O(N__1040),
            .I(N__1037));
    Sp12to4 I__151 (
            .O(N__1037),
            .I(N__1034));
    Span12Mux_h I__150 (
            .O(N__1034),
            .I(N__1031));
    Span12Mux_v I__149 (
            .O(N__1031),
            .I(N__1028));
    Span12Mux_v I__148 (
            .O(N__1028),
            .I(N__1025));
    Span12Mux_h I__147 (
            .O(N__1025),
            .I(N__1022));
    Odrv12 I__146 (
            .O(N__1022),
            .I(AD3_c_4));
    IoInMux I__145 (
            .O(N__1019),
            .I(N__1016));
    LocalMux I__144 (
            .O(N__1016),
            .I(N__1013));
    IoSpan4Mux I__143 (
            .O(N__1013),
            .I(N__1010));
    Span4Mux_s2_v I__142 (
            .O(N__1010),
            .I(N__1007));
    Sp12to4 I__141 (
            .O(N__1007),
            .I(N__1004));
    Span12Mux_v I__140 (
            .O(N__1004),
            .I(N__1001));
    Span12Mux_v I__139 (
            .O(N__1001),
            .I(N__998));
    Odrv12 I__138 (
            .O(N__998),
            .I(AD2_c_4));
    IoInMux I__137 (
            .O(N__995),
            .I(N__992));
    LocalMux I__136 (
            .O(N__992),
            .I(N__989));
    IoSpan4Mux I__135 (
            .O(N__989),
            .I(N__986));
    Span4Mux_s0_v I__134 (
            .O(N__986),
            .I(N__983));
    Span4Mux_v I__133 (
            .O(N__983),
            .I(N__980));
    Sp12to4 I__132 (
            .O(N__980),
            .I(N__977));
    Span12Mux_v I__131 (
            .O(N__977),
            .I(N__974));
    Span12Mux_v I__130 (
            .O(N__974),
            .I(N__971));
    Odrv12 I__129 (
            .O(N__971),
            .I(AD2_c_5));
    IoInMux I__128 (
            .O(N__968),
            .I(N__965));
    LocalMux I__127 (
            .O(N__965),
            .I(N__962));
    Span4Mux_s3_v I__126 (
            .O(N__962),
            .I(N__959));
    Span4Mux_v I__125 (
            .O(N__959),
            .I(N__956));
    Sp12to4 I__124 (
            .O(N__956),
            .I(N__953));
    Span12Mux_s0_h I__123 (
            .O(N__953),
            .I(N__950));
    Span12Mux_v I__122 (
            .O(N__950),
            .I(N__947));
    Span12Mux_v I__121 (
            .O(N__947),
            .I(N__944));
    Odrv12 I__120 (
            .O(N__944),
            .I(AD3_c_3));
    IoInMux I__119 (
            .O(N__941),
            .I(N__938));
    LocalMux I__118 (
            .O(N__938),
            .I(N__935));
    IoSpan4Mux I__117 (
            .O(N__935),
            .I(N__932));
    IoSpan4Mux I__116 (
            .O(N__932),
            .I(N__929));
    Span4Mux_s2_h I__115 (
            .O(N__929),
            .I(N__926));
    Sp12to4 I__114 (
            .O(N__926),
            .I(N__923));
    Span12Mux_h I__113 (
            .O(N__923),
            .I(N__920));
    Span12Mux_h I__112 (
            .O(N__920),
            .I(N__917));
    Odrv12 I__111 (
            .O(N__917),
            .I(AD0_c_1));
    IoInMux I__110 (
            .O(N__914),
            .I(N__911));
    LocalMux I__109 (
            .O(N__911),
            .I(N__908));
    Span4Mux_s0_v I__108 (
            .O(N__908),
            .I(N__905));
    Sp12to4 I__107 (
            .O(N__905),
            .I(N__902));
    Span12Mux_h I__106 (
            .O(N__902),
            .I(N__899));
    Span12Mux_v I__105 (
            .O(N__899),
            .I(N__896));
    Odrv12 I__104 (
            .O(N__896),
            .I(AD1_c_6));
    IoInMux I__103 (
            .O(N__893),
            .I(N__890));
    LocalMux I__102 (
            .O(N__890),
            .I(N__887));
    IoSpan4Mux I__101 (
            .O(N__887),
            .I(N__884));
    Span4Mux_s2_h I__100 (
            .O(N__884),
            .I(N__881));
    Sp12to4 I__99 (
            .O(N__881),
            .I(N__878));
    Span12Mux_h I__98 (
            .O(N__878),
            .I(N__875));
    Span12Mux_v I__97 (
            .O(N__875),
            .I(N__872));
    Span12Mux_v I__96 (
            .O(N__872),
            .I(N__869));
    Span12Mux_h I__95 (
            .O(N__869),
            .I(N__866));
    Odrv12 I__94 (
            .O(N__866),
            .I(AD3_c_6));
    IoInMux I__93 (
            .O(N__863),
            .I(N__860));
    LocalMux I__92 (
            .O(N__860),
            .I(N__857));
    Span12Mux_s3_v I__91 (
            .O(N__857),
            .I(N__854));
    Span12Mux_v I__90 (
            .O(N__854),
            .I(N__851));
    Span12Mux_v I__89 (
            .O(N__851),
            .I(N__848));
    Odrv12 I__88 (
            .O(N__848),
            .I(AD2_c_3));
    IoInMux I__87 (
            .O(N__845),
            .I(N__842));
    LocalMux I__86 (
            .O(N__842),
            .I(N__839));
    IoSpan4Mux I__85 (
            .O(N__839),
            .I(N__836));
    Span4Mux_s3_v I__84 (
            .O(N__836),
            .I(N__833));
    Sp12to4 I__83 (
            .O(N__833),
            .I(N__830));
    Span12Mux_s11_v I__82 (
            .O(N__830),
            .I(N__827));
    Span12Mux_v I__81 (
            .O(N__827),
            .I(N__824));
    Odrv12 I__80 (
            .O(N__824),
            .I(AD3_c_0));
    IoInMux I__79 (
            .O(N__821),
            .I(N__818));
    LocalMux I__78 (
            .O(N__818),
            .I(N__815));
    Span4Mux_s1_v I__77 (
            .O(N__815),
            .I(N__812));
    Span4Mux_v I__76 (
            .O(N__812),
            .I(N__809));
    Sp12to4 I__75 (
            .O(N__809),
            .I(N__806));
    Span12Mux_h I__74 (
            .O(N__806),
            .I(N__803));
    Span12Mux_h I__73 (
            .O(N__803),
            .I(N__800));
    Odrv12 I__72 (
            .O(N__800),
            .I(AD0_c_2));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_1_11_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_11_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_11_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U109_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 28 2025 22:04:17

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    CMA : out std_logic_vector(10 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__11817\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \N_996_i\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \U712_CHIP_RAM.N_186_cascade_\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_i_i_a2_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_a2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_265_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_265\ : std_logic;
signal \U712_CHIP_RAM.N_236_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_426_cascade_\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_350_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_350\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_287\ : std_logic;
signal \U712_CHIP_RAM.un3_DMA_CYCLE_START\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_300_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_301\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_esr_RNIULZ0Z431\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_1\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_236\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_348\ : std_logic;
signal \U712_CHIP_RAM.N_437\ : std_logic;
signal \U712_CHIP_RAM.N_426\ : std_logic;
signal \U712_CHIP_RAM.N_76_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_328\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \U712_CHIP_RAM.N_438_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_336\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_438\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_247\ : std_logic;
signal \U712_CHIP_RAM.N_247_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_244\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_0\ : std_logic;
signal \C3_c\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.BANK0_9_u_0_0_a2_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_269_i_0_en_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_269_i_0_en_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \N_249_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1_tz_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_325_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_325\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_241_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_388_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_325_1\ : std_logic;
signal \U712_CHIP_RAM.N_381\ : std_logic;
signal \U712_CHIP_RAM.N_386\ : std_logic;
signal \U712_CHIP_RAM.N_434_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_439\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_335\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_1\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.N_351_cascade_\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.m17_i_0_o2_1_cascade_\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_REG_SM.C3_SYNC_RNI7UAPZ0Z_1_cascade_\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.m15_i_0_a2_0_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_289\ : std_logic;
signal \U712_REG_SM.N_358_cascade_\ : std_logic;
signal \U712_REG_SM.N_360\ : std_logic;
signal \U712_REG_SM.N_359\ : std_logic;
signal \U712_REG_SM.N_270_i\ : std_logic;
signal \U712_REG_SM.REG_TACK_7\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.N_340_cascade_\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_345\ : std_logic;
signal \U712_BYTE_ENABLE.N_374_cascade_\ : std_logic;
signal \N_51_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_10\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_322_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\ : std_logic;
signal \U712_CHIP_RAM.N_388\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_271_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_2_1\ : std_logic;
signal \U712_CHIP_RAM.N_317\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_434\ : std_logic;
signal \U712_CHIP_RAM.N_13\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_300\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_241\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.N_360_1_cascade_\ : std_logic;
signal \U712_REG_SM.C3_SYNC_RNI7UAPZ0Z_1\ : std_logic;
signal \U712_REG_SM.m17_i_0_o2_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_RNOZ0Z_0_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \U712_REG_SM.m17_i_0_o2_1\ : std_logic;
signal \U712_REG_SM.N_435\ : std_logic;
signal \U712_REG_SM.N_435_cascade_\ : std_logic;
signal \U712_REG_SM.N_363\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.ASn_0_sqmuxa\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.m17_i_0_o2\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \RnW_c\ : std_logic;
signal \WRITE_CYCLEm\ : std_logic;
signal \N_276\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_5_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_112\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_392\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \U712_BYTE_ENABLE.N_370\ : std_logic;
signal \U712_BYTE_ENABLE.N_369_cascade_\ : std_logic;
signal \N_55_i\ : std_logic;
signal \WEn_c\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0\ : std_logic;
signal \N_53_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_303\ : std_logic;
signal \UMBE_0_o2_i\ : std_logic;
signal \U712_BYTE_ENABLE_UUBE_i\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1Z0Z_0\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \N_57_i\ : std_logic;
signal \U712_BYTE_ENABLE.UUBE\ : std_logic;
signal \N_185\ : std_logic;
signal \N_44\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \N_303_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \DS_ENm\ : std_logic;
signal \A_c_0\ : std_logic;
signal \N_337_i\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    RAMENn <= \RAMENn_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__3986\,
            RESETB => \N__5729\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11817\,
            DIN => \N__11816\,
            DOUT => \N__11815\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11817\,
            PADOUT => \N__11816\,
            PADIN => \N__11815\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5501\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11808\,
            DIN => \N__11807\,
            DOUT => \N__11806\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11808\,
            PADOUT => \N__11807\,
            PADIN => \N__11806\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11799\,
            DIN => \N__11798\,
            DOUT => \N__11797\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11799\,
            PADOUT => \N__11798\,
            PADIN => \N__11797\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9209\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11790\,
            DIN => \N__11789\,
            DOUT => \N__11788\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11790\,
            PADOUT => \N__11789\,
            PADIN => \N__11788\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6803\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11781\,
            DIN => \N__11780\,
            DOUT => \N__11779\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11781\,
            PADOUT => \N__11780\,
            PADIN => \N__11779\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11772\,
            DIN => \N__11771\,
            DOUT => \N__11770\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11772\,
            PADOUT => \N__11771\,
            PADIN => \N__11770\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11763\,
            DIN => \N__11762\,
            DOUT => \N__11761\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11763\,
            PADOUT => \N__11762\,
            PADIN => \N__11761\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11754\,
            DIN => \N__11753\,
            DOUT => \N__11752\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11754\,
            PADOUT => \N__11753\,
            PADIN => \N__11752\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11745\,
            DIN => \N__11744\,
            DOUT => \N__11743\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11745\,
            PADOUT => \N__11744\,
            PADIN => \N__11743\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11736\,
            DIN => \N__11735\,
            DOUT => \N__11734\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11736\,
            PADOUT => \N__11735\,
            PADIN => \N__11734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11727\,
            DIN => \N__11726\,
            DOUT => \N__11725\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11727\,
            PADOUT => \N__11726\,
            PADIN => \N__11725\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8915\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11718\,
            DIN => \N__11717\,
            DOUT => \N__11716\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11718\,
            PADOUT => \N__11717\,
            PADIN => \N__11716\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8285\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11709\,
            DIN => \N__11708\,
            DOUT => \N__11707\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11709\,
            PADOUT => \N__11708\,
            PADIN => \N__11707\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11700\,
            DIN => \N__11699\,
            DOUT => \N__11698\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11700\,
            PADOUT => \N__11699\,
            PADIN => \N__11698\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11691\,
            DIN => \N__11690\,
            DOUT => \N__11689\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11691\,
            PADOUT => \N__11690\,
            PADIN => \N__11689\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11682\,
            DIN => \N__11681\,
            DOUT => \N__11680\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11682\,
            PADOUT => \N__11681\,
            PADIN => \N__11680\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4295\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11673\,
            DIN => \N__11672\,
            DOUT => \N__11671\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11673\,
            PADOUT => \N__11672\,
            PADIN => \N__11671\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11664\,
            DIN => \N__11663\,
            DOUT => \N__11662\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11664\,
            PADOUT => \N__11663\,
            PADIN => \N__11662\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11655\,
            DIN => \N__11654\,
            DOUT => \N__11653\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11655\,
            PADOUT => \N__11654\,
            PADIN => \N__11653\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8789\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11646\,
            DIN => \N__11645\,
            DOUT => \N__11644\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11646\,
            PADOUT => \N__11645\,
            PADIN => \N__11644\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11637\,
            DIN => \N__11636\,
            DOUT => \N__11635\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11637\,
            PADOUT => \N__11636\,
            PADIN => \N__11635\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7901\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11628\,
            DIN => \N__11627\,
            DOUT => \N__11626\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11628\,
            PADOUT => \N__11627\,
            PADIN => \N__11626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11619\,
            DIN => \N__11618\,
            DOUT => \N__11617\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11619\,
            PADOUT => \N__11618\,
            PADIN => \N__11617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9242\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11610\,
            DIN => \N__11609\,
            DOUT => \N__11608\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11610\,
            PADOUT => \N__11609\,
            PADIN => \N__11608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11601\,
            DIN => \N__11600\,
            DOUT => \N__11599\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11601\,
            PADOUT => \N__11600\,
            PADIN => \N__11599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11592\,
            DIN => \N__11591\,
            DOUT => \N__11590\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11592\,
            PADOUT => \N__11591\,
            PADIN => \N__11590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11583\,
            DIN => \N__11582\,
            DOUT => \N__11581\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11583\,
            PADOUT => \N__11582\,
            PADIN => \N__11581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11574\,
            DIN => \N__11573\,
            DOUT => \N__11572\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11574\,
            PADOUT => \N__11573\,
            PADIN => \N__11572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11565\,
            DIN => \N__11564\,
            DOUT => \N__11563\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11565\,
            PADOUT => \N__11564\,
            PADIN => \N__11563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4838\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11556\,
            DIN => \N__11555\,
            DOUT => \N__11554\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11556\,
            PADOUT => \N__11555\,
            PADIN => \N__11554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11547\,
            DIN => \N__11546\,
            DOUT => \N__11545\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11547\,
            PADOUT => \N__11546\,
            PADIN => \N__11545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11538\,
            DIN => \N__11537\,
            DOUT => \N__11536\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11538\,
            PADOUT => \N__11537\,
            PADIN => \N__11536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11529\,
            DIN => \N__11528\,
            DOUT => \N__11527\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11529\,
            PADOUT => \N__11528\,
            PADIN => \N__11527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11520\,
            DIN => \N__11519\,
            DOUT => \N__11518\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11520\,
            PADOUT => \N__11519\,
            PADIN => \N__11518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11511\,
            DIN => \N__11510\,
            DOUT => \N__11509\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11511\,
            PADOUT => \N__11510\,
            PADIN => \N__11509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7883\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11502\,
            DIN => \N__11501\,
            DOUT => \N__11500\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11502\,
            PADOUT => \N__11501\,
            PADIN => \N__11500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11493\,
            DIN => \N__11492\,
            DOUT => \N__11491\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11493\,
            PADOUT => \N__11492\,
            PADIN => \N__11491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4172\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11484\,
            DIN => \N__11483\,
            DOUT => \N__11482\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11484\,
            PADOUT => \N__11483\,
            PADIN => \N__11482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4093\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11475\,
            DIN => \N__11474\,
            DOUT => \N__11473\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11475\,
            PADOUT => \N__11474\,
            PADIN => \N__11473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4004\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11466\,
            DIN => \N__11465\,
            DOUT => \N__11464\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11466\,
            PADOUT => \N__11465\,
            PADIN => \N__11464\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11457\,
            DIN => \N__11456\,
            DOUT => \N__11455\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11457\,
            PADOUT => \N__11456\,
            PADIN => \N__11455\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7112\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11448\,
            DIN => \N__11447\,
            DOUT => \N__11446\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11448\,
            PADOUT => \N__11447\,
            PADIN => \N__11446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8081\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11439\,
            DIN => \N__11438\,
            DOUT => \N__11437\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11439\,
            PADOUT => \N__11438\,
            PADIN => \N__11437\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11430\,
            DIN => \N__11429\,
            DOUT => \N__11428\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11430\,
            PADOUT => \N__11429\,
            PADIN => \N__11428\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11421\,
            DIN => \N__11420\,
            DOUT => \N__11419\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11421\,
            PADOUT => \N__11420\,
            PADIN => \N__11419\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11412\,
            DIN => \N__11411\,
            DOUT => \N__11410\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11412\,
            PADOUT => \N__11411\,
            PADIN => \N__11410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11403\,
            DIN => \N__11402\,
            DOUT => \N__11401\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11403\,
            PADOUT => \N__11402\,
            PADIN => \N__11401\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11394\,
            DIN => \N__11393\,
            DOUT => \N__11392\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11394\,
            PADOUT => \N__11393\,
            PADIN => \N__11392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8138\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11385\,
            DIN => \N__11384\,
            DOUT => \N__11383\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11385\,
            PADOUT => \N__11384\,
            PADIN => \N__11383\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11376\,
            DIN => \N__11375\,
            DOUT => \N__11374\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11376\,
            PADOUT => \N__11375\,
            PADIN => \N__11374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4081\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11367\,
            DIN => \N__11366\,
            DOUT => \N__11365\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11367\,
            PADOUT => \N__11366\,
            PADIN => \N__11365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9182\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11358\,
            DIN => \N__11357\,
            DOUT => \N__11356\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11358\,
            PADOUT => \N__11357\,
            PADIN => \N__11356\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10649\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11349\,
            DIN => \N__11348\,
            DOUT => \N__11347\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11349\,
            PADOUT => \N__11348\,
            PADIN => \N__11347\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5750\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11340\,
            DIN => \N__11339\,
            DOUT => \N__11338\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11340\,
            PADOUT => \N__11339\,
            PADIN => \N__11338\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8717\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11331\,
            DIN => \N__11330\,
            DOUT => \N__11329\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11331\,
            PADOUT => \N__11330\,
            PADIN => \N__11329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7111\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11322\,
            DIN => \N__11321\,
            DOUT => \N__11320\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11322\,
            PADOUT => \N__11321\,
            PADIN => \N__11320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11313\,
            DIN => \N__11312\,
            DOUT => \N__11311\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11313\,
            PADOUT => \N__11312\,
            PADIN => \N__11311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11304\,
            DIN => \N__11303\,
            DOUT => \N__11302\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11304\,
            PADOUT => \N__11303\,
            PADIN => \N__11302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8330\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11295\,
            DIN => \N__11294\,
            DOUT => \N__11293\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11295\,
            PADOUT => \N__11294\,
            PADIN => \N__11293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7919\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11286\,
            DIN => \N__11285\,
            DOUT => \N__11284\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11286\,
            PADOUT => \N__11285\,
            PADIN => \N__11284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4142\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11277\,
            DIN => \N__11276\,
            DOUT => \N__11275\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11277\,
            PADOUT => \N__11276\,
            PADIN => \N__11275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7943\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11268\,
            DIN => \N__11267\,
            DOUT => \N__11266\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11268\,
            PADOUT => \N__11267\,
            PADIN => \N__11266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11259\,
            DIN => \N__11258\,
            DOUT => \N__11257\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11259\,
            PADOUT => \N__11258\,
            PADIN => \N__11257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11250\,
            DIN => \N__11249\,
            DOUT => \N__11248\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11250\,
            PADOUT => \N__11249\,
            PADIN => \N__11248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11241\,
            DIN => \N__11240\,
            DOUT => \N__11239\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11241\,
            PADOUT => \N__11240\,
            PADIN => \N__11239\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11232\,
            DIN => \N__11231\,
            DOUT => \N__11230\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11232\,
            PADOUT => \N__11231\,
            PADIN => \N__11230\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7307\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11223\,
            DIN => \N__11222\,
            DOUT => \N__11221\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11223\,
            PADOUT => \N__11222\,
            PADIN => \N__11221\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10388\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11214\,
            DIN => \N__11213\,
            DOUT => \N__11212\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11214\,
            PADOUT => \N__11213\,
            PADIN => \N__11212\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11205\,
            DIN => \N__11204\,
            DOUT => \N__11203\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11205\,
            PADOUT => \N__11204\,
            PADIN => \N__11203\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9272\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11196\,
            DIN => \N__11195\,
            DOUT => \N__11194\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11196\,
            PADOUT => \N__11195\,
            PADIN => \N__11194\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4022\,
            DIN0 => OPEN,
            DOUT0 => \N__4121\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11187\,
            DIN => \N__11186\,
            DOUT => \N__11185\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11187\,
            PADOUT => \N__11186\,
            PADIN => \N__11185\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8093\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11178\,
            DIN => \N__11177\,
            DOUT => \N__11176\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11178\,
            PADOUT => \N__11177\,
            PADIN => \N__11176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11169\,
            DIN => \N__11168\,
            DOUT => \N__11167\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11169\,
            PADOUT => \N__11168\,
            PADIN => \N__11167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11160\,
            DIN => \N__11159\,
            DOUT => \N__11158\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11160\,
            PADOUT => \N__11159\,
            PADIN => \N__11158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9140\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11151\,
            DIN => \N__11150\,
            DOUT => \N__11149\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11151\,
            PADOUT => \N__11150\,
            PADIN => \N__11149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11142\,
            DIN => \N__11141\,
            DOUT => \N__11140\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11142\,
            PADOUT => \N__11141\,
            PADIN => \N__11140\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11133\,
            DIN => \N__11132\,
            DOUT => \N__11131\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11133\,
            PADOUT => \N__11132\,
            PADIN => \N__11131\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11124\,
            DIN => \N__11123\,
            DOUT => \N__11122\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11124\,
            PADOUT => \N__11123\,
            PADIN => \N__11122\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11115\,
            DIN => \N__11114\,
            DOUT => \N__11113\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11115\,
            PADOUT => \N__11114\,
            PADIN => \N__11113\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7769\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11106\,
            DIN => \N__11105\,
            DOUT => \N__11104\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11106\,
            PADOUT => \N__11105\,
            PADIN => \N__11104\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10082\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11097\,
            DIN => \N__11096\,
            DOUT => \N__11095\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11097\,
            PADOUT => \N__11096\,
            PADIN => \N__11095\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8303\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11088\,
            DIN => \N__11087\,
            DOUT => \N__11086\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11088\,
            PADOUT => \N__11087\,
            PADIN => \N__11086\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7232\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11079\,
            DIN => \N__11078\,
            DOUT => \N__11077\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11079\,
            PADOUT => \N__11078\,
            PADIN => \N__11077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11070\,
            DIN => \N__11069\,
            DOUT => \N__11068\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11070\,
            PADOUT => \N__11069\,
            PADIN => \N__11068\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11061\,
            DIN => \N__11060\,
            DOUT => \N__11059\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11061\,
            PADOUT => \N__11060\,
            PADIN => \N__11059\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8939\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11052\,
            DIN => \N__11051\,
            DOUT => \N__11050\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11052\,
            PADOUT => \N__11051\,
            PADIN => \N__11050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11043\,
            DIN => \N__11042\,
            DOUT => \N__11041\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11043\,
            PADOUT => \N__11042\,
            PADIN => \N__11041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11034\,
            DIN => \N__11033\,
            DOUT => \N__11032\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11034\,
            PADOUT => \N__11033\,
            PADIN => \N__11032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4643\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11025\,
            DIN => \N__11024\,
            DOUT => \N__11023\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11025\,
            PADOUT => \N__11024\,
            PADIN => \N__11023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9227\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11016\,
            DIN => \N__11015\,
            DOUT => \N__11014\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11016\,
            PADOUT => \N__11015\,
            PADIN => \N__11014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4097\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2687\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10991\
        );

    \I__2686\ : InMux
    port map (
            O => \N__10996\,
            I => \N__10988\
        );

    \I__2685\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10985\
        );

    \I__2684\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10982\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__10991\,
            I => \N__10979\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__10988\,
            I => \N__10969\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__10985\,
            I => \N__10959\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__10982\,
            I => \N__10946\
        );

    \I__2679\ : Glb2LocalMux
    port map (
            O => \N__10979\,
            I => \N__10853\
        );

    \I__2678\ : SRMux
    port map (
            O => \N__10978\,
            I => \N__10853\
        );

    \I__2677\ : SRMux
    port map (
            O => \N__10977\,
            I => \N__10853\
        );

    \I__2676\ : SRMux
    port map (
            O => \N__10976\,
            I => \N__10853\
        );

    \I__2675\ : SRMux
    port map (
            O => \N__10975\,
            I => \N__10853\
        );

    \I__2674\ : SRMux
    port map (
            O => \N__10974\,
            I => \N__10853\
        );

    \I__2673\ : SRMux
    port map (
            O => \N__10973\,
            I => \N__10853\
        );

    \I__2672\ : SRMux
    port map (
            O => \N__10972\,
            I => \N__10853\
        );

    \I__2671\ : Glb2LocalMux
    port map (
            O => \N__10969\,
            I => \N__10853\
        );

    \I__2670\ : SRMux
    port map (
            O => \N__10968\,
            I => \N__10853\
        );

    \I__2669\ : SRMux
    port map (
            O => \N__10967\,
            I => \N__10853\
        );

    \I__2668\ : SRMux
    port map (
            O => \N__10966\,
            I => \N__10853\
        );

    \I__2667\ : SRMux
    port map (
            O => \N__10965\,
            I => \N__10853\
        );

    \I__2666\ : SRMux
    port map (
            O => \N__10964\,
            I => \N__10853\
        );

    \I__2665\ : SRMux
    port map (
            O => \N__10963\,
            I => \N__10853\
        );

    \I__2664\ : SRMux
    port map (
            O => \N__10962\,
            I => \N__10853\
        );

    \I__2663\ : Glb2LocalMux
    port map (
            O => \N__10959\,
            I => \N__10853\
        );

    \I__2662\ : SRMux
    port map (
            O => \N__10958\,
            I => \N__10853\
        );

    \I__2661\ : SRMux
    port map (
            O => \N__10957\,
            I => \N__10853\
        );

    \I__2660\ : SRMux
    port map (
            O => \N__10956\,
            I => \N__10853\
        );

    \I__2659\ : SRMux
    port map (
            O => \N__10955\,
            I => \N__10853\
        );

    \I__2658\ : SRMux
    port map (
            O => \N__10954\,
            I => \N__10853\
        );

    \I__2657\ : SRMux
    port map (
            O => \N__10953\,
            I => \N__10853\
        );

    \I__2656\ : SRMux
    port map (
            O => \N__10952\,
            I => \N__10853\
        );

    \I__2655\ : SRMux
    port map (
            O => \N__10951\,
            I => \N__10853\
        );

    \I__2654\ : SRMux
    port map (
            O => \N__10950\,
            I => \N__10853\
        );

    \I__2653\ : SRMux
    port map (
            O => \N__10949\,
            I => \N__10853\
        );

    \I__2652\ : Glb2LocalMux
    port map (
            O => \N__10946\,
            I => \N__10853\
        );

    \I__2651\ : SRMux
    port map (
            O => \N__10945\,
            I => \N__10853\
        );

    \I__2650\ : SRMux
    port map (
            O => \N__10944\,
            I => \N__10853\
        );

    \I__2649\ : SRMux
    port map (
            O => \N__10943\,
            I => \N__10853\
        );

    \I__2648\ : SRMux
    port map (
            O => \N__10942\,
            I => \N__10853\
        );

    \I__2647\ : SRMux
    port map (
            O => \N__10941\,
            I => \N__10853\
        );

    \I__2646\ : SRMux
    port map (
            O => \N__10940\,
            I => \N__10853\
        );

    \I__2645\ : SRMux
    port map (
            O => \N__10939\,
            I => \N__10853\
        );

    \I__2644\ : SRMux
    port map (
            O => \N__10938\,
            I => \N__10853\
        );

    \I__2643\ : SRMux
    port map (
            O => \N__10937\,
            I => \N__10853\
        );

    \I__2642\ : SRMux
    port map (
            O => \N__10936\,
            I => \N__10853\
        );

    \I__2641\ : SRMux
    port map (
            O => \N__10935\,
            I => \N__10853\
        );

    \I__2640\ : SRMux
    port map (
            O => \N__10934\,
            I => \N__10853\
        );

    \I__2639\ : GlobalMux
    port map (
            O => \N__10853\,
            I => \N__10850\
        );

    \I__2638\ : gio2CtrlBuf
    port map (
            O => \N__10850\,
            I => \RESETn_c_i_g\
        );

    \I__2637\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10844\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__10844\,
            I => \N__10840\
        );

    \I__2635\ : InMux
    port map (
            O => \N__10843\,
            I => \N__10836\
        );

    \I__2634\ : Sp12to4
    port map (
            O => \N__10840\,
            I => \N__10833\
        );

    \I__2633\ : InMux
    port map (
            O => \N__10839\,
            I => \N__10830\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__10836\,
            I => \N__10827\
        );

    \I__2631\ : Span12Mux_v
    port map (
            O => \N__10833\,
            I => \N__10823\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__10830\,
            I => \N__10820\
        );

    \I__2629\ : Span4Mux_v
    port map (
            O => \N__10827\,
            I => \N__10817\
        );

    \I__2628\ : InMux
    port map (
            O => \N__10826\,
            I => \N__10813\
        );

    \I__2627\ : Span12Mux_h
    port map (
            O => \N__10823\,
            I => \N__10810\
        );

    \I__2626\ : Span12Mux_v
    port map (
            O => \N__10820\,
            I => \N__10807\
        );

    \I__2625\ : Span4Mux_v
    port map (
            O => \N__10817\,
            I => \N__10804\
        );

    \I__2624\ : InMux
    port map (
            O => \N__10816\,
            I => \N__10801\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__10813\,
            I => \N__10798\
        );

    \I__2622\ : Odrv12
    port map (
            O => \N__10810\,
            I => \REG_CYCLEm\
        );

    \I__2621\ : Odrv12
    port map (
            O => \N__10807\,
            I => \REG_CYCLEm\
        );

    \I__2620\ : Odrv4
    port map (
            O => \N__10804\,
            I => \REG_CYCLEm\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__10801\,
            I => \REG_CYCLEm\
        );

    \I__2618\ : Odrv4
    port map (
            O => \N__10798\,
            I => \REG_CYCLEm\
        );

    \I__2617\ : InMux
    port map (
            O => \N__10787\,
            I => \N__10784\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__10784\,
            I => \N__10781\
        );

    \I__2615\ : Span4Mux_h
    port map (
            O => \N__10781\,
            I => \N__10777\
        );

    \I__2614\ : InMux
    port map (
            O => \N__10780\,
            I => \N__10773\
        );

    \I__2613\ : Span4Mux_h
    port map (
            O => \N__10777\,
            I => \N__10769\
        );

    \I__2612\ : InMux
    port map (
            O => \N__10776\,
            I => \N__10765\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__10773\,
            I => \N__10762\
        );

    \I__2610\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10759\
        );

    \I__2609\ : Span4Mux_h
    port map (
            O => \N__10769\,
            I => \N__10756\
        );

    \I__2608\ : InMux
    port map (
            O => \N__10768\,
            I => \N__10753\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__10765\,
            I => \N__10750\
        );

    \I__2606\ : Sp12to4
    port map (
            O => \N__10762\,
            I => \N__10745\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__10759\,
            I => \N__10745\
        );

    \I__2604\ : Span4Mux_h
    port map (
            O => \N__10756\,
            I => \N__10740\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__10753\,
            I => \N__10740\
        );

    \I__2602\ : Span12Mux_h
    port map (
            O => \N__10750\,
            I => \N__10737\
        );

    \I__2601\ : Span12Mux_v
    port map (
            O => \N__10745\,
            I => \N__10734\
        );

    \I__2600\ : Span4Mux_h
    port map (
            O => \N__10740\,
            I => \N__10731\
        );

    \I__2599\ : Span12Mux_v
    port map (
            O => \N__10737\,
            I => \N__10728\
        );

    \I__2598\ : Span12Mux_h
    port map (
            O => \N__10734\,
            I => \N__10725\
        );

    \I__2597\ : Span4Mux_v
    port map (
            O => \N__10731\,
            I => \N__10722\
        );

    \I__2596\ : Odrv12
    port map (
            O => \N__10728\,
            I => \CASUn_c\
        );

    \I__2595\ : Odrv12
    port map (
            O => \N__10725\,
            I => \CASUn_c\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__10722\,
            I => \CASUn_c\
        );

    \I__2593\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10711\
        );

    \I__2592\ : InMux
    port map (
            O => \N__10714\,
            I => \N__10708\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__10711\,
            I => \N__10705\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__10708\,
            I => \N__10702\
        );

    \I__2589\ : Span4Mux_v
    port map (
            O => \N__10705\,
            I => \N__10695\
        );

    \I__2588\ : Span4Mux_v
    port map (
            O => \N__10702\,
            I => \N__10695\
        );

    \I__2587\ : InMux
    port map (
            O => \N__10701\,
            I => \N__10692\
        );

    \I__2586\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10689\
        );

    \I__2585\ : Sp12to4
    port map (
            O => \N__10695\,
            I => \N__10685\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__10692\,
            I => \N__10682\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__10689\,
            I => \N__10679\
        );

    \I__2582\ : InMux
    port map (
            O => \N__10688\,
            I => \N__10676\
        );

    \I__2581\ : Span12Mux_h
    port map (
            O => \N__10685\,
            I => \N__10673\
        );

    \I__2580\ : Span12Mux_v
    port map (
            O => \N__10682\,
            I => \N__10670\
        );

    \I__2579\ : Span12Mux_v
    port map (
            O => \N__10679\,
            I => \N__10667\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__10676\,
            I => \N__10664\
        );

    \I__2577\ : Span12Mux_v
    port map (
            O => \N__10673\,
            I => \N__10659\
        );

    \I__2576\ : Span12Mux_h
    port map (
            O => \N__10670\,
            I => \N__10659\
        );

    \I__2575\ : Span12Mux_h
    port map (
            O => \N__10667\,
            I => \N__10654\
        );

    \I__2574\ : Span12Mux_v
    port map (
            O => \N__10664\,
            I => \N__10654\
        );

    \I__2573\ : Odrv12
    port map (
            O => \N__10659\,
            I => \CASLn_c\
        );

    \I__2572\ : Odrv12
    port map (
            O => \N__10654\,
            I => \CASLn_c\
        );

    \I__2571\ : IoInMux
    port map (
            O => \N__10649\,
            I => \N__10646\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__10646\,
            I => \N__10643\
        );

    \I__2569\ : Span4Mux_s3_v
    port map (
            O => \N__10643\,
            I => \N__10640\
        );

    \I__2568\ : Span4Mux_v
    port map (
            O => \N__10640\,
            I => \N__10637\
        );

    \I__2567\ : Odrv4
    port map (
            O => \N__10637\,
            I => \DRDENn_c\
        );

    \I__2566\ : InMux
    port map (
            O => \N__10634\,
            I => \N__10629\
        );

    \I__2565\ : InMux
    port map (
            O => \N__10633\,
            I => \N__10625\
        );

    \I__2564\ : InMux
    port map (
            O => \N__10632\,
            I => \N__10622\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__10629\,
            I => \N__10616\
        );

    \I__2562\ : InMux
    port map (
            O => \N__10628\,
            I => \N__10613\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__10625\,
            I => \N__10610\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__10622\,
            I => \N__10607\
        );

    \I__2559\ : InMux
    port map (
            O => \N__10621\,
            I => \N__10602\
        );

    \I__2558\ : InMux
    port map (
            O => \N__10620\,
            I => \N__10602\
        );

    \I__2557\ : InMux
    port map (
            O => \N__10619\,
            I => \N__10599\
        );

    \I__2556\ : Span4Mux_v
    port map (
            O => \N__10616\,
            I => \N__10596\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__10613\,
            I => \N__10593\
        );

    \I__2554\ : Span4Mux_v
    port map (
            O => \N__10610\,
            I => \N__10590\
        );

    \I__2553\ : Span4Mux_v
    port map (
            O => \N__10607\,
            I => \N__10587\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10602\,
            I => \N__10584\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__10599\,
            I => \N__10580\
        );

    \I__2550\ : Span4Mux_v
    port map (
            O => \N__10596\,
            I => \N__10575\
        );

    \I__2549\ : Span4Mux_v
    port map (
            O => \N__10593\,
            I => \N__10575\
        );

    \I__2548\ : Span4Mux_v
    port map (
            O => \N__10590\,
            I => \N__10568\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__10587\,
            I => \N__10568\
        );

    \I__2546\ : Span4Mux_v
    port map (
            O => \N__10584\,
            I => \N__10568\
        );

    \I__2545\ : InMux
    port map (
            O => \N__10583\,
            I => \N__10565\
        );

    \I__2544\ : Span12Mux_v
    port map (
            O => \N__10580\,
            I => \N__10562\
        );

    \I__2543\ : Sp12to4
    port map (
            O => \N__10575\,
            I => \N__10555\
        );

    \I__2542\ : Sp12to4
    port map (
            O => \N__10568\,
            I => \N__10555\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__10565\,
            I => \N__10555\
        );

    \I__2540\ : Span12Mux_h
    port map (
            O => \N__10562\,
            I => \N__10552\
        );

    \I__2539\ : Span12Mux_h
    port map (
            O => \N__10555\,
            I => \N__10549\
        );

    \I__2538\ : Odrv12
    port map (
            O => \N__10552\,
            I => \A_c_1\
        );

    \I__2537\ : Odrv12
    port map (
            O => \N__10549\,
            I => \A_c_1\
        );

    \I__2536\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10541\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__10541\,
            I => \N__10535\
        );

    \I__2534\ : InMux
    port map (
            O => \N__10540\,
            I => \N__10532\
        );

    \I__2533\ : InMux
    port map (
            O => \N__10539\,
            I => \N__10529\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__10538\,
            I => \N__10525\
        );

    \I__2531\ : Span4Mux_v
    port map (
            O => \N__10535\,
            I => \N__10521\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__10532\,
            I => \N__10518\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__10529\,
            I => \N__10515\
        );

    \I__2528\ : InMux
    port map (
            O => \N__10528\,
            I => \N__10510\
        );

    \I__2527\ : InMux
    port map (
            O => \N__10525\,
            I => \N__10510\
        );

    \I__2526\ : InMux
    port map (
            O => \N__10524\,
            I => \N__10507\
        );

    \I__2525\ : Span4Mux_h
    port map (
            O => \N__10521\,
            I => \N__10502\
        );

    \I__2524\ : Span4Mux_v
    port map (
            O => \N__10518\,
            I => \N__10502\
        );

    \I__2523\ : Span4Mux_v
    port map (
            O => \N__10515\,
            I => \N__10495\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__10510\,
            I => \N__10495\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__10507\,
            I => \N__10495\
        );

    \I__2520\ : Span4Mux_v
    port map (
            O => \N__10502\,
            I => \N__10492\
        );

    \I__2519\ : Span4Mux_h
    port map (
            O => \N__10495\,
            I => \N__10489\
        );

    \I__2518\ : Span4Mux_v
    port map (
            O => \N__10492\,
            I => \N__10486\
        );

    \I__2517\ : Span4Mux_v
    port map (
            O => \N__10489\,
            I => \N__10483\
        );

    \I__2516\ : Sp12to4
    port map (
            O => \N__10486\,
            I => \N__10478\
        );

    \I__2515\ : Sp12to4
    port map (
            O => \N__10483\,
            I => \N__10478\
        );

    \I__2514\ : Span12Mux_h
    port map (
            O => \N__10478\,
            I => \N__10475\
        );

    \I__2513\ : Odrv12
    port map (
            O => \N__10475\,
            I => \SIZ_c_0\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__10472\,
            I => \N__10469\
        );

    \I__2511\ : InMux
    port map (
            O => \N__10469\,
            I => \N__10465\
        );

    \I__2510\ : InMux
    port map (
            O => \N__10468\,
            I => \N__10462\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__10465\,
            I => \N__10454\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10462\,
            I => \N__10454\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__10461\,
            I => \N__10448\
        );

    \I__2506\ : InMux
    port map (
            O => \N__10460\,
            I => \N__10443\
        );

    \I__2505\ : InMux
    port map (
            O => \N__10459\,
            I => \N__10443\
        );

    \I__2504\ : Span4Mux_v
    port map (
            O => \N__10454\,
            I => \N__10440\
        );

    \I__2503\ : InMux
    port map (
            O => \N__10453\,
            I => \N__10437\
        );

    \I__2502\ : InMux
    port map (
            O => \N__10452\,
            I => \N__10432\
        );

    \I__2501\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10432\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10448\,
            I => \N__10429\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__10443\,
            I => \N__10426\
        );

    \I__2498\ : Span4Mux_v
    port map (
            O => \N__10440\,
            I => \N__10423\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__10437\,
            I => \N__10416\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__10432\,
            I => \N__10416\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__10429\,
            I => \N__10416\
        );

    \I__2494\ : Sp12to4
    port map (
            O => \N__10426\,
            I => \N__10413\
        );

    \I__2493\ : Span4Mux_v
    port map (
            O => \N__10423\,
            I => \N__10410\
        );

    \I__2492\ : Sp12to4
    port map (
            O => \N__10416\,
            I => \N__10407\
        );

    \I__2491\ : Span12Mux_v
    port map (
            O => \N__10413\,
            I => \N__10404\
        );

    \I__2490\ : Sp12to4
    port map (
            O => \N__10410\,
            I => \N__10399\
        );

    \I__2489\ : Span12Mux_v
    port map (
            O => \N__10407\,
            I => \N__10399\
        );

    \I__2488\ : Span12Mux_h
    port map (
            O => \N__10404\,
            I => \N__10396\
        );

    \I__2487\ : Span12Mux_h
    port map (
            O => \N__10399\,
            I => \N__10393\
        );

    \I__2486\ : Odrv12
    port map (
            O => \N__10396\,
            I => \SIZ_c_1\
        );

    \I__2485\ : Odrv12
    port map (
            O => \N__10393\,
            I => \SIZ_c_1\
        );

    \I__2484\ : IoInMux
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__2482\ : Span4Mux_s2_v
    port map (
            O => \N__10382\,
            I => \N__10379\
        );

    \I__2481\ : Span4Mux_v
    port map (
            O => \N__10379\,
            I => \N__10376\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__10376\,
            I => \N_303_i\
        );

    \I__2479\ : InMux
    port map (
            O => \N__10373\,
            I => \N__10370\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__10370\,
            I => \N__10367\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__10367\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2476\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10358\
        );

    \I__2475\ : InMux
    port map (
            O => \N__10363\,
            I => \N__10355\
        );

    \I__2474\ : InMux
    port map (
            O => \N__10362\,
            I => \N__10352\
        );

    \I__2473\ : InMux
    port map (
            O => \N__10361\,
            I => \N__10349\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__10358\,
            I => \N__10340\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__10355\,
            I => \N__10340\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__10352\,
            I => \N__10340\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__10349\,
            I => \N__10340\
        );

    \I__2468\ : Span4Mux_v
    port map (
            O => \N__10340\,
            I => \N__10337\
        );

    \I__2467\ : Sp12to4
    port map (
            O => \N__10337\,
            I => \N__10334\
        );

    \I__2466\ : Span12Mux_h
    port map (
            O => \N__10334\,
            I => \N__10331\
        );

    \I__2465\ : Odrv12
    port map (
            O => \N__10331\,
            I => \DRA_c_8\
        );

    \I__2464\ : InMux
    port map (
            O => \N__10328\,
            I => \N__10325\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__10325\,
            I => \N__10322\
        );

    \I__2462\ : Span4Mux_h
    port map (
            O => \N__10322\,
            I => \N__10319\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__10319\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2460\ : InMux
    port map (
            O => \N__10316\,
            I => \N__10313\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__10313\,
            I => \N__10310\
        );

    \I__2458\ : Span12Mux_v
    port map (
            O => \N__10310\,
            I => \N__10307\
        );

    \I__2457\ : Odrv12
    port map (
            O => \N__10307\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2456\ : InMux
    port map (
            O => \N__10304\,
            I => \N__10301\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__10301\,
            I => \N__10296\
        );

    \I__2454\ : InMux
    port map (
            O => \N__10300\,
            I => \N__10293\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10299\,
            I => \N__10290\
        );

    \I__2452\ : Span4Mux_v
    port map (
            O => \N__10296\,
            I => \N__10285\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__10293\,
            I => \N__10285\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10290\,
            I => \N__10282\
        );

    \I__2449\ : Span4Mux_v
    port map (
            O => \N__10285\,
            I => \N__10278\
        );

    \I__2448\ : Span4Mux_v
    port map (
            O => \N__10282\,
            I => \N__10275\
        );

    \I__2447\ : InMux
    port map (
            O => \N__10281\,
            I => \N__10272\
        );

    \I__2446\ : Sp12to4
    port map (
            O => \N__10278\,
            I => \N__10269\
        );

    \I__2445\ : Sp12to4
    port map (
            O => \N__10275\,
            I => \N__10264\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__10272\,
            I => \N__10264\
        );

    \I__2443\ : Span12Mux_v
    port map (
            O => \N__10269\,
            I => \N__10261\
        );

    \I__2442\ : Span12Mux_h
    port map (
            O => \N__10264\,
            I => \N__10258\
        );

    \I__2441\ : Span12Mux_h
    port map (
            O => \N__10261\,
            I => \N__10253\
        );

    \I__2440\ : Span12Mux_v
    port map (
            O => \N__10258\,
            I => \N__10253\
        );

    \I__2439\ : Odrv12
    port map (
            O => \N__10253\,
            I => \DRA_c_1\
        );

    \I__2438\ : InMux
    port map (
            O => \N__10250\,
            I => \N__10247\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__10247\,
            I => \N__10243\
        );

    \I__2436\ : InMux
    port map (
            O => \N__10246\,
            I => \N__10240\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__10243\,
            I => \N__10235\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__10240\,
            I => \N__10235\
        );

    \I__2433\ : Sp12to4
    port map (
            O => \N__10235\,
            I => \N__10232\
        );

    \I__2432\ : Span12Mux_v
    port map (
            O => \N__10232\,
            I => \N__10229\
        );

    \I__2431\ : Span12Mux_h
    port map (
            O => \N__10229\,
            I => \N__10226\
        );

    \I__2430\ : Odrv12
    port map (
            O => \N__10226\,
            I => \DRA_c_0\
        );

    \I__2429\ : InMux
    port map (
            O => \N__10223\,
            I => \N__10220\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__10220\,
            I => \N__10217\
        );

    \I__2427\ : Odrv4
    port map (
            O => \N__10217\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2426\ : InMux
    port map (
            O => \N__10214\,
            I => \N__10211\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__10211\,
            I => \N__10207\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__10210\,
            I => \N__10204\
        );

    \I__2423\ : Span4Mux_h
    port map (
            O => \N__10207\,
            I => \N__10201\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10204\,
            I => \N__10198\
        );

    \I__2421\ : Sp12to4
    port map (
            O => \N__10201\,
            I => \N__10193\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__10198\,
            I => \N__10193\
        );

    \I__2419\ : Span12Mux_v
    port map (
            O => \N__10193\,
            I => \N__10189\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10192\,
            I => \N__10186\
        );

    \I__2417\ : Odrv12
    port map (
            O => \N__10189\,
            I => \DS_ENm\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__10186\,
            I => \DS_ENm\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__10181\,
            I => \N__10171\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10180\,
            I => \N__10165\
        );

    \I__2413\ : InMux
    port map (
            O => \N__10179\,
            I => \N__10165\
        );

    \I__2412\ : InMux
    port map (
            O => \N__10178\,
            I => \N__10162\
        );

    \I__2411\ : InMux
    port map (
            O => \N__10177\,
            I => \N__10158\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10176\,
            I => \N__10155\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10175\,
            I => \N__10150\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10174\,
            I => \N__10150\
        );

    \I__2407\ : InMux
    port map (
            O => \N__10171\,
            I => \N__10147\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__10170\,
            I => \N__10144\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__10165\,
            I => \N__10141\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10162\,
            I => \N__10138\
        );

    \I__2403\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10135\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__10158\,
            I => \N__10132\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__10155\,
            I => \N__10125\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__10150\,
            I => \N__10125\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__10147\,
            I => \N__10125\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10144\,
            I => \N__10122\
        );

    \I__2397\ : Span4Mux_v
    port map (
            O => \N__10141\,
            I => \N__10117\
        );

    \I__2396\ : Span4Mux_v
    port map (
            O => \N__10138\,
            I => \N__10117\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__10135\,
            I => \N__10114\
        );

    \I__2394\ : Span4Mux_v
    port map (
            O => \N__10132\,
            I => \N__10109\
        );

    \I__2393\ : Span4Mux_v
    port map (
            O => \N__10125\,
            I => \N__10109\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__10122\,
            I => \N__10106\
        );

    \I__2391\ : Sp12to4
    port map (
            O => \N__10117\,
            I => \N__10101\
        );

    \I__2390\ : Span12Mux_v
    port map (
            O => \N__10114\,
            I => \N__10101\
        );

    \I__2389\ : Sp12to4
    port map (
            O => \N__10109\,
            I => \N__10098\
        );

    \I__2388\ : Span4Mux_v
    port map (
            O => \N__10106\,
            I => \N__10095\
        );

    \I__2387\ : Span12Mux_h
    port map (
            O => \N__10101\,
            I => \N__10092\
        );

    \I__2386\ : Span12Mux_h
    port map (
            O => \N__10098\,
            I => \N__10087\
        );

    \I__2385\ : Sp12to4
    port map (
            O => \N__10095\,
            I => \N__10087\
        );

    \I__2384\ : Odrv12
    port map (
            O => \N__10092\,
            I => \A_c_0\
        );

    \I__2383\ : Odrv12
    port map (
            O => \N__10087\,
            I => \A_c_0\
        );

    \I__2382\ : IoInMux
    port map (
            O => \N__10082\,
            I => \N__10079\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__10079\,
            I => \N__10076\
        );

    \I__2380\ : Span4Mux_s3_v
    port map (
            O => \N__10076\,
            I => \N__10073\
        );

    \I__2379\ : Span4Mux_h
    port map (
            O => \N__10073\,
            I => \N__10070\
        );

    \I__2378\ : Span4Mux_h
    port map (
            O => \N__10070\,
            I => \N__10067\
        );

    \I__2377\ : Odrv4
    port map (
            O => \N__10067\,
            I => \N_337_i\
        );

    \I__2376\ : InMux
    port map (
            O => \N__10064\,
            I => \N__10061\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__10061\,
            I => \N__10058\
        );

    \I__2374\ : Span4Mux_v
    port map (
            O => \N__10058\,
            I => \N__10052\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10057\,
            I => \N__10049\
        );

    \I__2372\ : InMux
    port map (
            O => \N__10056\,
            I => \N__10046\
        );

    \I__2371\ : InMux
    port map (
            O => \N__10055\,
            I => \N__10043\
        );

    \I__2370\ : Span4Mux_v
    port map (
            O => \N__10052\,
            I => \N__10036\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__10049\,
            I => \N__10036\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__10046\,
            I => \N__10036\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10043\,
            I => \N__10033\
        );

    \I__2366\ : Span4Mux_h
    port map (
            O => \N__10036\,
            I => \N__10028\
        );

    \I__2365\ : Span4Mux_v
    port map (
            O => \N__10033\,
            I => \N__10028\
        );

    \I__2364\ : Span4Mux_v
    port map (
            O => \N__10028\,
            I => \N__10025\
        );

    \I__2363\ : Sp12to4
    port map (
            O => \N__10025\,
            I => \N__10022\
        );

    \I__2362\ : Odrv12
    port map (
            O => \N__10022\,
            I => \DRA_c_6\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__10019\,
            I => \N__10016\
        );

    \I__2360\ : InMux
    port map (
            O => \N__10016\,
            I => \N__10011\
        );

    \I__2359\ : InMux
    port map (
            O => \N__10015\,
            I => \N__10008\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10014\,
            I => \N__10005\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__10011\,
            I => \N__9997\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10008\,
            I => \N__9997\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__10005\,
            I => \N__9997\
        );

    \I__2354\ : InMux
    port map (
            O => \N__10004\,
            I => \N__9994\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__9997\,
            I => \N__9991\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__9994\,
            I => \N__9988\
        );

    \I__2351\ : Sp12to4
    port map (
            O => \N__9991\,
            I => \N__9983\
        );

    \I__2350\ : Span12Mux_v
    port map (
            O => \N__9988\,
            I => \N__9983\
        );

    \I__2349\ : Span12Mux_h
    port map (
            O => \N__9983\,
            I => \N__9980\
        );

    \I__2348\ : Odrv12
    port map (
            O => \N__9980\,
            I => \DRA_c_7\
        );

    \I__2347\ : InMux
    port map (
            O => \N__9977\,
            I => \N__9974\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__9974\,
            I => \N__9971\
        );

    \I__2345\ : Span4Mux_h
    port map (
            O => \N__9971\,
            I => \N__9968\
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__9968\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2343\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9960\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__9964\,
            I => \N__9954\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__9963\,
            I => \N__9951\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__9960\,
            I => \N__9941\
        );

    \I__2339\ : InMux
    port map (
            O => \N__9959\,
            I => \N__9936\
        );

    \I__2338\ : InMux
    port map (
            O => \N__9958\,
            I => \N__9936\
        );

    \I__2337\ : InMux
    port map (
            O => \N__9957\,
            I => \N__9933\
        );

    \I__2336\ : InMux
    port map (
            O => \N__9954\,
            I => \N__9926\
        );

    \I__2335\ : InMux
    port map (
            O => \N__9951\,
            I => \N__9926\
        );

    \I__2334\ : InMux
    port map (
            O => \N__9950\,
            I => \N__9926\
        );

    \I__2333\ : InMux
    port map (
            O => \N__9949\,
            I => \N__9921\
        );

    \I__2332\ : InMux
    port map (
            O => \N__9948\,
            I => \N__9921\
        );

    \I__2331\ : InMux
    port map (
            O => \N__9947\,
            I => \N__9918\
        );

    \I__2330\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9915\
        );

    \I__2329\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9912\
        );

    \I__2328\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9908\
        );

    \I__2327\ : Span4Mux_v
    port map (
            O => \N__9941\,
            I => \N__9900\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__9936\,
            I => \N__9887\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__9933\,
            I => \N__9887\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__9926\,
            I => \N__9887\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__9921\,
            I => \N__9887\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__9918\,
            I => \N__9887\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__9915\,
            I => \N__9887\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__9912\,
            I => \N__9884\
        );

    \I__2319\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9881\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__9908\,
            I => \N__9878\
        );

    \I__2317\ : InMux
    port map (
            O => \N__9907\,
            I => \N__9873\
        );

    \I__2316\ : InMux
    port map (
            O => \N__9906\,
            I => \N__9873\
        );

    \I__2315\ : InMux
    port map (
            O => \N__9905\,
            I => \N__9870\
        );

    \I__2314\ : InMux
    port map (
            O => \N__9904\,
            I => \N__9867\
        );

    \I__2313\ : InMux
    port map (
            O => \N__9903\,
            I => \N__9864\
        );

    \I__2312\ : Span4Mux_h
    port map (
            O => \N__9900\,
            I => \N__9857\
        );

    \I__2311\ : Span4Mux_v
    port map (
            O => \N__9887\,
            I => \N__9857\
        );

    \I__2310\ : Span4Mux_v
    port map (
            O => \N__9884\,
            I => \N__9852\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__9881\,
            I => \N__9852\
        );

    \I__2308\ : Span4Mux_v
    port map (
            O => \N__9878\,
            I => \N__9841\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__9873\,
            I => \N__9841\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__9870\,
            I => \N__9841\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__9867\,
            I => \N__9841\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__9864\,
            I => \N__9841\
        );

    \I__2303\ : InMux
    port map (
            O => \N__9863\,
            I => \N__9838\
        );

    \I__2302\ : InMux
    port map (
            O => \N__9862\,
            I => \N__9835\
        );

    \I__2301\ : Span4Mux_h
    port map (
            O => \N__9857\,
            I => \N__9830\
        );

    \I__2300\ : Span4Mux_v
    port map (
            O => \N__9852\,
            I => \N__9830\
        );

    \I__2299\ : Span4Mux_v
    port map (
            O => \N__9841\,
            I => \N__9827\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__9838\,
            I => \N__9822\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__9835\,
            I => \N__9822\
        );

    \I__2296\ : Sp12to4
    port map (
            O => \N__9830\,
            I => \N__9817\
        );

    \I__2295\ : Sp12to4
    port map (
            O => \N__9827\,
            I => \N__9817\
        );

    \I__2294\ : Span12Mux_h
    port map (
            O => \N__9822\,
            I => \N__9814\
        );

    \I__2293\ : Span12Mux_h
    port map (
            O => \N__9817\,
            I => \N__9811\
        );

    \I__2292\ : Span12Mux_v
    port map (
            O => \N__9814\,
            I => \N__9808\
        );

    \I__2291\ : Span12Mux_v
    port map (
            O => \N__9811\,
            I => \N__9805\
        );

    \I__2290\ : Odrv12
    port map (
            O => \N__9808\,
            I => \AGNUS_REV_c\
        );

    \I__2289\ : Odrv12
    port map (
            O => \N__9805\,
            I => \AGNUS_REV_c\
        );

    \I__2288\ : InMux
    port map (
            O => \N__9800\,
            I => \N__9797\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__9797\,
            I => \N__9794\
        );

    \I__2286\ : Span4Mux_v
    port map (
            O => \N__9794\,
            I => \N__9791\
        );

    \I__2285\ : Sp12to4
    port map (
            O => \N__9791\,
            I => \N__9788\
        );

    \I__2284\ : Odrv12
    port map (
            O => \N__9788\,
            I => \RAS0n_c\
        );

    \I__2283\ : InMux
    port map (
            O => \N__9785\,
            I => \N__9780\
        );

    \I__2282\ : InMux
    port map (
            O => \N__9784\,
            I => \N__9777\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__9783\,
            I => \N__9774\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__9780\,
            I => \N__9769\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__9777\,
            I => \N__9769\
        );

    \I__2278\ : InMux
    port map (
            O => \N__9774\,
            I => \N__9766\
        );

    \I__2277\ : Span4Mux_v
    port map (
            O => \N__9769\,
            I => \N__9762\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__9766\,
            I => \N__9759\
        );

    \I__2275\ : InMux
    port map (
            O => \N__9765\,
            I => \N__9756\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__9762\,
            I => \N__9753\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__9759\,
            I => \N__9750\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__9756\,
            I => \N__9747\
        );

    \I__2271\ : Sp12to4
    port map (
            O => \N__9753\,
            I => \N__9742\
        );

    \I__2270\ : Sp12to4
    port map (
            O => \N__9750\,
            I => \N__9742\
        );

    \I__2269\ : Sp12to4
    port map (
            O => \N__9747\,
            I => \N__9739\
        );

    \I__2268\ : Span12Mux_h
    port map (
            O => \N__9742\,
            I => \N__9736\
        );

    \I__2267\ : Span12Mux_v
    port map (
            O => \N__9739\,
            I => \N__9733\
        );

    \I__2266\ : Span12Mux_v
    port map (
            O => \N__9736\,
            I => \N__9730\
        );

    \I__2265\ : Span12Mux_v
    port map (
            O => \N__9733\,
            I => \N__9727\
        );

    \I__2264\ : Odrv12
    port map (
            O => \N__9730\,
            I => \DRA_c_9\
        );

    \I__2263\ : Odrv12
    port map (
            O => \N__9727\,
            I => \DRA_c_9\
        );

    \I__2262\ : InMux
    port map (
            O => \N__9722\,
            I => \N__9719\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__9719\,
            I => \N__9716\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__9716\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2259\ : ClkMux
    port map (
            O => \N__9713\,
            I => \N__9692\
        );

    \I__2258\ : ClkMux
    port map (
            O => \N__9712\,
            I => \N__9692\
        );

    \I__2257\ : ClkMux
    port map (
            O => \N__9711\,
            I => \N__9692\
        );

    \I__2256\ : ClkMux
    port map (
            O => \N__9710\,
            I => \N__9692\
        );

    \I__2255\ : ClkMux
    port map (
            O => \N__9709\,
            I => \N__9692\
        );

    \I__2254\ : ClkMux
    port map (
            O => \N__9708\,
            I => \N__9692\
        );

    \I__2253\ : ClkMux
    port map (
            O => \N__9707\,
            I => \N__9692\
        );

    \I__2252\ : GlobalMux
    port map (
            O => \N__9692\,
            I => \N__9689\
        );

    \I__2251\ : gio2CtrlBuf
    port map (
            O => \N__9689\,
            I => \C3_c_g\
        );

    \I__2250\ : CEMux
    port map (
            O => \N__9686\,
            I => \N__9644\
        );

    \I__2249\ : CEMux
    port map (
            O => \N__9685\,
            I => \N__9644\
        );

    \I__2248\ : CEMux
    port map (
            O => \N__9684\,
            I => \N__9644\
        );

    \I__2247\ : CEMux
    port map (
            O => \N__9683\,
            I => \N__9644\
        );

    \I__2246\ : CEMux
    port map (
            O => \N__9682\,
            I => \N__9644\
        );

    \I__2245\ : CEMux
    port map (
            O => \N__9681\,
            I => \N__9644\
        );

    \I__2244\ : CEMux
    port map (
            O => \N__9680\,
            I => \N__9644\
        );

    \I__2243\ : CEMux
    port map (
            O => \N__9679\,
            I => \N__9644\
        );

    \I__2242\ : CEMux
    port map (
            O => \N__9678\,
            I => \N__9644\
        );

    \I__2241\ : CEMux
    port map (
            O => \N__9677\,
            I => \N__9644\
        );

    \I__2240\ : CEMux
    port map (
            O => \N__9676\,
            I => \N__9644\
        );

    \I__2239\ : CEMux
    port map (
            O => \N__9675\,
            I => \N__9644\
        );

    \I__2238\ : CEMux
    port map (
            O => \N__9674\,
            I => \N__9644\
        );

    \I__2237\ : CEMux
    port map (
            O => \N__9673\,
            I => \N__9644\
        );

    \I__2236\ : GlobalMux
    port map (
            O => \N__9644\,
            I => \N__9641\
        );

    \I__2235\ : gio2CtrlBuf
    port map (
            O => \N__9641\,
            I => \DBRn_c_i_0_g\
        );

    \I__2234\ : InMux
    port map (
            O => \N__9638\,
            I => \N__9635\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__9635\,
            I => \N__9632\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__9632\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2231\ : InMux
    port map (
            O => \N__9629\,
            I => \N__9626\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__9626\,
            I => \N__9623\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__9623\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2228\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9617\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__9617\,
            I => \N__9611\
        );

    \I__2226\ : InMux
    port map (
            O => \N__9616\,
            I => \N__9606\
        );

    \I__2225\ : InMux
    port map (
            O => \N__9615\,
            I => \N__9606\
        );

    \I__2224\ : InMux
    port map (
            O => \N__9614\,
            I => \N__9603\
        );

    \I__2223\ : Span4Mux_h
    port map (
            O => \N__9611\,
            I => \N__9598\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__9606\,
            I => \N__9598\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__9603\,
            I => \N__9593\
        );

    \I__2220\ : Sp12to4
    port map (
            O => \N__9598\,
            I => \N__9593\
        );

    \I__2219\ : Span12Mux_v
    port map (
            O => \N__9593\,
            I => \N__9590\
        );

    \I__2218\ : Span12Mux_h
    port map (
            O => \N__9590\,
            I => \N__9587\
        );

    \I__2217\ : Odrv12
    port map (
            O => \N__9587\,
            I => \DRA_c_5\
        );

    \I__2216\ : InMux
    port map (
            O => \N__9584\,
            I => \N__9578\
        );

    \I__2215\ : InMux
    port map (
            O => \N__9583\,
            I => \N__9575\
        );

    \I__2214\ : InMux
    port map (
            O => \N__9582\,
            I => \N__9572\
        );

    \I__2213\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9569\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__9578\,
            I => \N__9564\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__9575\,
            I => \N__9564\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9572\,
            I => \N__9561\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__9569\,
            I => \N__9558\
        );

    \I__2208\ : Span4Mux_v
    port map (
            O => \N__9564\,
            I => \N__9555\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__9561\,
            I => \N__9552\
        );

    \I__2206\ : Span4Mux_h
    port map (
            O => \N__9558\,
            I => \N__9549\
        );

    \I__2205\ : Span4Mux_v
    port map (
            O => \N__9555\,
            I => \N__9546\
        );

    \I__2204\ : Span4Mux_v
    port map (
            O => \N__9552\,
            I => \N__9543\
        );

    \I__2203\ : Sp12to4
    port map (
            O => \N__9549\,
            I => \N__9540\
        );

    \I__2202\ : Sp12to4
    port map (
            O => \N__9546\,
            I => \N__9537\
        );

    \I__2201\ : Sp12to4
    port map (
            O => \N__9543\,
            I => \N__9532\
        );

    \I__2200\ : Span12Mux_v
    port map (
            O => \N__9540\,
            I => \N__9532\
        );

    \I__2199\ : Span12Mux_h
    port map (
            O => \N__9537\,
            I => \N__9529\
        );

    \I__2198\ : Span12Mux_h
    port map (
            O => \N__9532\,
            I => \N__9526\
        );

    \I__2197\ : Odrv12
    port map (
            O => \N__9529\,
            I => \DRA_c_4\
        );

    \I__2196\ : Odrv12
    port map (
            O => \N__9526\,
            I => \DRA_c_4\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9521\,
            I => \N__9518\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__9518\,
            I => \N__9515\
        );

    \I__2193\ : Odrv12
    port map (
            O => \N__9515\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9512\,
            I => \N__9509\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__9509\,
            I => \N__9506\
        );

    \I__2190\ : Span4Mux_h
    port map (
            O => \N__9506\,
            I => \N__9503\
        );

    \I__2189\ : Span4Mux_h
    port map (
            O => \N__9503\,
            I => \N__9500\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__9500\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9497\,
            I => \N__9493\
        );

    \I__2186\ : InMux
    port map (
            O => \N__9496\,
            I => \N__9490\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__9493\,
            I => \N__9487\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__9490\,
            I => \N__9484\
        );

    \I__2183\ : Span4Mux_h
    port map (
            O => \N__9487\,
            I => \N__9479\
        );

    \I__2182\ : Span4Mux_v
    port map (
            O => \N__9484\,
            I => \N__9479\
        );

    \I__2181\ : Odrv4
    port map (
            O => \N__9479\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1Z0Z_0\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__9476\,
            I => \N__9471\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__9475\,
            I => \N__9465\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__9474\,
            I => \N__9462\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9471\,
            I => \N__9457\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__9470\,
            I => \N__9449\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__9469\,
            I => \N__9444\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9468\,
            I => \N__9437\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9465\,
            I => \N__9434\
        );

    \I__2172\ : InMux
    port map (
            O => \N__9462\,
            I => \N__9431\
        );

    \I__2171\ : InMux
    port map (
            O => \N__9461\,
            I => \N__9426\
        );

    \I__2170\ : InMux
    port map (
            O => \N__9460\,
            I => \N__9426\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__9457\,
            I => \N__9423\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9456\,
            I => \N__9420\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9455\,
            I => \N__9417\
        );

    \I__2166\ : InMux
    port map (
            O => \N__9454\,
            I => \N__9414\
        );

    \I__2165\ : InMux
    port map (
            O => \N__9453\,
            I => \N__9410\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9452\,
            I => \N__9405\
        );

    \I__2163\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9405\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9448\,
            I => \N__9400\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9447\,
            I => \N__9400\
        );

    \I__2160\ : InMux
    port map (
            O => \N__9444\,
            I => \N__9397\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9443\,
            I => \N__9392\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9442\,
            I => \N__9392\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9441\,
            I => \N__9389\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9440\,
            I => \N__9386\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9437\,
            I => \N__9380\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9434\,
            I => \N__9380\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__9431\,
            I => \N__9375\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__9426\,
            I => \N__9375\
        );

    \I__2151\ : Span4Mux_v
    port map (
            O => \N__9423\,
            I => \N__9368\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__9420\,
            I => \N__9368\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__9417\,
            I => \N__9368\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9414\,
            I => \N__9365\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9362\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__9410\,
            I => \N__9355\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__9405\,
            I => \N__9355\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__9400\,
            I => \N__9355\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9397\,
            I => \N__9350\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9392\,
            I => \N__9350\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__9389\,
            I => \N__9345\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__9386\,
            I => \N__9345\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9385\,
            I => \N__9342\
        );

    \I__2138\ : Span4Mux_v
    port map (
            O => \N__9380\,
            I => \N__9334\
        );

    \I__2137\ : Span4Mux_v
    port map (
            O => \N__9375\,
            I => \N__9334\
        );

    \I__2136\ : Span4Mux_v
    port map (
            O => \N__9368\,
            I => \N__9325\
        );

    \I__2135\ : Span4Mux_v
    port map (
            O => \N__9365\,
            I => \N__9325\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9362\,
            I => \N__9325\
        );

    \I__2133\ : Span4Mux_h
    port map (
            O => \N__9355\,
            I => \N__9325\
        );

    \I__2132\ : Span4Mux_h
    port map (
            O => \N__9350\,
            I => \N__9322\
        );

    \I__2131\ : Span4Mux_v
    port map (
            O => \N__9345\,
            I => \N__9317\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__9342\,
            I => \N__9314\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9341\,
            I => \N__9311\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9340\,
            I => \N__9306\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9306\
        );

    \I__2126\ : Span4Mux_h
    port map (
            O => \N__9334\,
            I => \N__9303\
        );

    \I__2125\ : Span4Mux_h
    port map (
            O => \N__9325\,
            I => \N__9300\
        );

    \I__2124\ : Span4Mux_h
    port map (
            O => \N__9322\,
            I => \N__9297\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9321\,
            I => \N__9294\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9291\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__9317\,
            I => \CPU_CYCLEm\
        );

    \I__2120\ : Odrv12
    port map (
            O => \N__9314\,
            I => \CPU_CYCLEm\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__9311\,
            I => \CPU_CYCLEm\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9306\,
            I => \CPU_CYCLEm\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__9303\,
            I => \CPU_CYCLEm\
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__9300\,
            I => \CPU_CYCLEm\
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__9297\,
            I => \CPU_CYCLEm\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__9294\,
            I => \CPU_CYCLEm\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__9291\,
            I => \CPU_CYCLEm\
        );

    \I__2112\ : IoInMux
    port map (
            O => \N__9272\,
            I => \N__9269\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__9269\,
            I => \N__9266\
        );

    \I__2110\ : Span4Mux_s3_h
    port map (
            O => \N__9266\,
            I => \N__9263\
        );

    \I__2109\ : Span4Mux_v
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__2108\ : Span4Mux_v
    port map (
            O => \N__9260\,
            I => \N__9257\
        );

    \I__2107\ : Sp12to4
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__2106\ : Odrv12
    port map (
            O => \N__9254\,
            I => \N_57_i\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__9251\,
            I => \N__9248\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9245\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__9245\,
            I => \U712_BYTE_ENABLE.UUBE\
        );

    \I__2102\ : IoInMux
    port map (
            O => \N__9242\,
            I => \N__9239\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9239\,
            I => \N__9236\
        );

    \I__2100\ : Span4Mux_s3_v
    port map (
            O => \N__9236\,
            I => \N__9233\
        );

    \I__2099\ : Span4Mux_v
    port map (
            O => \N__9233\,
            I => \N__9230\
        );

    \I__2098\ : Odrv4
    port map (
            O => \N__9230\,
            I => \N_185\
        );

    \I__2097\ : IoInMux
    port map (
            O => \N__9227\,
            I => \N__9224\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__9224\,
            I => \N__9221\
        );

    \I__2095\ : Span4Mux_s3_v
    port map (
            O => \N__9221\,
            I => \N__9218\
        );

    \I__2094\ : Sp12to4
    port map (
            O => \N__9218\,
            I => \N__9215\
        );

    \I__2093\ : Span12Mux_h
    port map (
            O => \N__9215\,
            I => \N__9212\
        );

    \I__2092\ : Odrv12
    port map (
            O => \N__9212\,
            I => \N_44\
        );

    \I__2091\ : IoInMux
    port map (
            O => \N__9209\,
            I => \N__9206\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9206\,
            I => \N__9203\
        );

    \I__2089\ : IoSpan4Mux
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__2088\ : Span4Mux_s2_v
    port map (
            O => \N__9200\,
            I => \N__9197\
        );

    \I__2087\ : Span4Mux_v
    port map (
            O => \N__9197\,
            I => \N__9194\
        );

    \I__2086\ : Span4Mux_h
    port map (
            O => \N__9194\,
            I => \N__9191\
        );

    \I__2085\ : Odrv4
    port map (
            O => \N__9191\,
            I => \CASn_c\
        );

    \I__2084\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9185\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__9185\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__2082\ : IoInMux
    port map (
            O => \N__9182\,
            I => \N__9179\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__9179\,
            I => \N__9176\
        );

    \I__2080\ : IoSpan4Mux
    port map (
            O => \N__9176\,
            I => \N__9173\
        );

    \I__2079\ : Span4Mux_s3_h
    port map (
            O => \N__9173\,
            I => \N__9170\
        );

    \I__2078\ : Sp12to4
    port map (
            O => \N__9170\,
            I => \N__9167\
        );

    \I__2077\ : Span12Mux_h
    port map (
            O => \N__9167\,
            I => \N__9164\
        );

    \I__2076\ : Odrv12
    port map (
            O => \N__9164\,
            I => \CMA_c_4\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9161\,
            I => \N__9158\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__9158\,
            I => \N__9155\
        );

    \I__2073\ : Span4Mux_v
    port map (
            O => \N__9155\,
            I => \N__9152\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__9152\,
            I => \N__9149\
        );

    \I__2071\ : Sp12to4
    port map (
            O => \N__9149\,
            I => \N__9146\
        );

    \I__2070\ : Span12Mux_h
    port map (
            O => \N__9146\,
            I => \N__9143\
        );

    \I__2069\ : Odrv12
    port map (
            O => \N__9143\,
            I => \A_c_17\
        );

    \I__2068\ : IoInMux
    port map (
            O => \N__9140\,
            I => \N__9137\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__9137\,
            I => \N__9134\
        );

    \I__2066\ : Span12Mux_s2_h
    port map (
            O => \N__9134\,
            I => \N__9131\
        );

    \I__2065\ : Span12Mux_h
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__2064\ : Odrv12
    port map (
            O => \N__9128\,
            I => \CMA_c_8\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9125\,
            I => \N__9122\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__2061\ : Odrv12
    port map (
            O => \N__9119\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__9116\,
            I => \N__9108\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__9115\,
            I => \N__9105\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__9114\,
            I => \N__9099\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__9113\,
            I => \N__9096\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9112\,
            I => \N__9092\
        );

    \I__2055\ : InMux
    port map (
            O => \N__9111\,
            I => \N__9089\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9108\,
            I => \N__9084\
        );

    \I__2053\ : InMux
    port map (
            O => \N__9105\,
            I => \N__9084\
        );

    \I__2052\ : InMux
    port map (
            O => \N__9104\,
            I => \N__9079\
        );

    \I__2051\ : InMux
    port map (
            O => \N__9103\,
            I => \N__9079\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__9102\,
            I => \N__9075\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9070\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9066\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__9095\,
            I => \N__9063\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__9092\,
            I => \N__9055\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__9089\,
            I => \N__9050\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__9084\,
            I => \N__9045\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__9079\,
            I => \N__9045\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9078\,
            I => \N__9038\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9038\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9038\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9035\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__9070\,
            I => \N__9031\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9069\,
            I => \N__9028\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9066\,
            I => \N__9025\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9063\,
            I => \N__9020\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9020\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9061\,
            I => \N__9015\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9060\,
            I => \N__9015\
        );

    \I__2031\ : InMux
    port map (
            O => \N__9059\,
            I => \N__9010\
        );

    \I__2030\ : InMux
    port map (
            O => \N__9058\,
            I => \N__9010\
        );

    \I__2029\ : Span4Mux_v
    port map (
            O => \N__9055\,
            I => \N__9005\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9054\,
            I => \N__9002\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9053\,
            I => \N__8999\
        );

    \I__2026\ : Span4Mux_h
    port map (
            O => \N__9050\,
            I => \N__8990\
        );

    \I__2025\ : Span4Mux_v
    port map (
            O => \N__9045\,
            I => \N__8990\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9038\,
            I => \N__8990\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9035\,
            I => \N__8990\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9034\,
            I => \N__8987\
        );

    \I__2021\ : Span4Mux_h
    port map (
            O => \N__9031\,
            I => \N__8984\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__9028\,
            I => \N__8981\
        );

    \I__2019\ : Sp12to4
    port map (
            O => \N__9025\,
            I => \N__8972\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__9020\,
            I => \N__8972\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__9015\,
            I => \N__8972\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9010\,
            I => \N__8972\
        );

    \I__2015\ : InMux
    port map (
            O => \N__9009\,
            I => \N__8967\
        );

    \I__2014\ : InMux
    port map (
            O => \N__9008\,
            I => \N__8967\
        );

    \I__2013\ : Span4Mux_h
    port map (
            O => \N__9005\,
            I => \N__8960\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__9002\,
            I => \N__8960\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__8999\,
            I => \N__8960\
        );

    \I__2010\ : Span4Mux_h
    port map (
            O => \N__8990\,
            I => \N__8957\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__8987\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__8984\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__8981\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2006\ : Odrv12
    port map (
            O => \N__8972\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__8967\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__8960\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__8957\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__8942\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_\
        );

    \I__2001\ : IoInMux
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__8936\,
            I => \N__8933\
        );

    \I__1999\ : Span12Mux_s2_h
    port map (
            O => \N__8933\,
            I => \N__8930\
        );

    \I__1998\ : Span12Mux_h
    port map (
            O => \N__8930\,
            I => \N__8927\
        );

    \I__1997\ : Odrv12
    port map (
            O => \N__8927\,
            I => \CMA_c_6\
        );

    \I__1996\ : InMux
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__1994\ : Odrv12
    port map (
            O => \N__8918\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1993\ : IoInMux
    port map (
            O => \N__8915\,
            I => \N__8912\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__8912\,
            I => \N__8909\
        );

    \I__1991\ : Span12Mux_s2_h
    port map (
            O => \N__8909\,
            I => \N__8906\
        );

    \I__1990\ : Span12Mux_h
    port map (
            O => \N__8906\,
            I => \N__8903\
        );

    \I__1989\ : Odrv12
    port map (
            O => \N__8903\,
            I => \CMA_c_7\
        );

    \I__1988\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8892\
        );

    \I__1987\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8889\
        );

    \I__1986\ : InMux
    port map (
            O => \N__8898\,
            I => \N__8884\
        );

    \I__1985\ : InMux
    port map (
            O => \N__8897\,
            I => \N__8884\
        );

    \I__1984\ : InMux
    port map (
            O => \N__8896\,
            I => \N__8879\
        );

    \I__1983\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8879\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__8892\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__8889\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__8884\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__8879\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__8870\,
            I => \N__8864\
        );

    \I__1977\ : CascadeMux
    port map (
            O => \N__8869\,
            I => \N__8860\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__8868\,
            I => \N__8857\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__8867\,
            I => \N__8853\
        );

    \I__1974\ : InMux
    port map (
            O => \N__8864\,
            I => \N__8850\
        );

    \I__1973\ : InMux
    port map (
            O => \N__8863\,
            I => \N__8847\
        );

    \I__1972\ : InMux
    port map (
            O => \N__8860\,
            I => \N__8844\
        );

    \I__1971\ : InMux
    port map (
            O => \N__8857\,
            I => \N__8841\
        );

    \I__1970\ : InMux
    port map (
            O => \N__8856\,
            I => \N__8838\
        );

    \I__1969\ : InMux
    port map (
            O => \N__8853\,
            I => \N__8835\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__8850\,
            I => \N__8832\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__8847\,
            I => \N__8827\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__8844\,
            I => \N__8827\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__8841\,
            I => \N__8822\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__8838\,
            I => \N__8815\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__8835\,
            I => \N__8815\
        );

    \I__1962\ : Span4Mux_h
    port map (
            O => \N__8832\,
            I => \N__8815\
        );

    \I__1961\ : Span4Mux_h
    port map (
            O => \N__8827\,
            I => \N__8812\
        );

    \I__1960\ : InMux
    port map (
            O => \N__8826\,
            I => \N__8809\
        );

    \I__1959\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8806\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__8822\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__8815\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__8812\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__8809\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__8806\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1953\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8792\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__8792\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1951\ : IoInMux
    port map (
            O => \N__8789\,
            I => \N__8786\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__8786\,
            I => \N__8783\
        );

    \I__1949\ : Span4Mux_s3_v
    port map (
            O => \N__8783\,
            I => \N__8780\
        );

    \I__1948\ : Span4Mux_v
    port map (
            O => \N__8780\,
            I => \N__8777\
        );

    \I__1947\ : Span4Mux_v
    port map (
            O => \N__8777\,
            I => \N__8774\
        );

    \I__1946\ : Odrv4
    port map (
            O => \N__8774\,
            I => \CMA_c_0\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8771\,
            I => \N__8767\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8764\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__8767\,
            I => \N__8759\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__8764\,
            I => \N__8756\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8763\,
            I => \N__8751\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8762\,
            I => \N__8751\
        );

    \I__1939\ : Span4Mux_v
    port map (
            O => \N__8759\,
            I => \N__8746\
        );

    \I__1938\ : Span4Mux_v
    port map (
            O => \N__8756\,
            I => \N__8746\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__8751\,
            I => \N__8743\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__8746\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__8743\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1934\ : InMux
    port map (
            O => \N__8738\,
            I => \N__8735\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__8735\,
            I => \N__8732\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__8732\,
            I => \N__8729\
        );

    \I__1931\ : Sp12to4
    port map (
            O => \N__8729\,
            I => \N__8726\
        );

    \I__1930\ : Span12Mux_v
    port map (
            O => \N__8726\,
            I => \N__8723\
        );

    \I__1929\ : Span12Mux_h
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__1928\ : Odrv12
    port map (
            O => \N__8720\,
            I => \A_c_19\
        );

    \I__1927\ : IoInMux
    port map (
            O => \N__8717\,
            I => \N__8714\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__8714\,
            I => \N__8711\
        );

    \I__1925\ : IoSpan4Mux
    port map (
            O => \N__8711\,
            I => \N__8708\
        );

    \I__1924\ : IoSpan4Mux
    port map (
            O => \N__8708\,
            I => \N__8705\
        );

    \I__1923\ : Sp12to4
    port map (
            O => \N__8705\,
            I => \N__8702\
        );

    \I__1922\ : Span12Mux_s7_h
    port map (
            O => \N__8702\,
            I => \N__8699\
        );

    \I__1921\ : Odrv12
    port map (
            O => \N__8699\,
            I => \CMA_c_9\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8696\,
            I => \N__8693\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__8693\,
            I => \N__8662\
        );

    \I__1918\ : ClkMux
    port map (
            O => \N__8692\,
            I => \N__8579\
        );

    \I__1917\ : ClkMux
    port map (
            O => \N__8691\,
            I => \N__8579\
        );

    \I__1916\ : ClkMux
    port map (
            O => \N__8690\,
            I => \N__8579\
        );

    \I__1915\ : ClkMux
    port map (
            O => \N__8689\,
            I => \N__8579\
        );

    \I__1914\ : ClkMux
    port map (
            O => \N__8688\,
            I => \N__8579\
        );

    \I__1913\ : ClkMux
    port map (
            O => \N__8687\,
            I => \N__8579\
        );

    \I__1912\ : ClkMux
    port map (
            O => \N__8686\,
            I => \N__8579\
        );

    \I__1911\ : ClkMux
    port map (
            O => \N__8685\,
            I => \N__8579\
        );

    \I__1910\ : ClkMux
    port map (
            O => \N__8684\,
            I => \N__8579\
        );

    \I__1909\ : ClkMux
    port map (
            O => \N__8683\,
            I => \N__8579\
        );

    \I__1908\ : ClkMux
    port map (
            O => \N__8682\,
            I => \N__8579\
        );

    \I__1907\ : ClkMux
    port map (
            O => \N__8681\,
            I => \N__8579\
        );

    \I__1906\ : ClkMux
    port map (
            O => \N__8680\,
            I => \N__8579\
        );

    \I__1905\ : ClkMux
    port map (
            O => \N__8679\,
            I => \N__8579\
        );

    \I__1904\ : ClkMux
    port map (
            O => \N__8678\,
            I => \N__8579\
        );

    \I__1903\ : ClkMux
    port map (
            O => \N__8677\,
            I => \N__8579\
        );

    \I__1902\ : ClkMux
    port map (
            O => \N__8676\,
            I => \N__8579\
        );

    \I__1901\ : ClkMux
    port map (
            O => \N__8675\,
            I => \N__8579\
        );

    \I__1900\ : ClkMux
    port map (
            O => \N__8674\,
            I => \N__8579\
        );

    \I__1899\ : ClkMux
    port map (
            O => \N__8673\,
            I => \N__8579\
        );

    \I__1898\ : ClkMux
    port map (
            O => \N__8672\,
            I => \N__8579\
        );

    \I__1897\ : ClkMux
    port map (
            O => \N__8671\,
            I => \N__8579\
        );

    \I__1896\ : ClkMux
    port map (
            O => \N__8670\,
            I => \N__8579\
        );

    \I__1895\ : ClkMux
    port map (
            O => \N__8669\,
            I => \N__8579\
        );

    \I__1894\ : ClkMux
    port map (
            O => \N__8668\,
            I => \N__8579\
        );

    \I__1893\ : ClkMux
    port map (
            O => \N__8667\,
            I => \N__8579\
        );

    \I__1892\ : ClkMux
    port map (
            O => \N__8666\,
            I => \N__8579\
        );

    \I__1891\ : ClkMux
    port map (
            O => \N__8665\,
            I => \N__8579\
        );

    \I__1890\ : Glb2LocalMux
    port map (
            O => \N__8662\,
            I => \N__8579\
        );

    \I__1889\ : ClkMux
    port map (
            O => \N__8661\,
            I => \N__8579\
        );

    \I__1888\ : ClkMux
    port map (
            O => \N__8660\,
            I => \N__8579\
        );

    \I__1887\ : ClkMux
    port map (
            O => \N__8659\,
            I => \N__8579\
        );

    \I__1886\ : ClkMux
    port map (
            O => \N__8658\,
            I => \N__8579\
        );

    \I__1885\ : ClkMux
    port map (
            O => \N__8657\,
            I => \N__8579\
        );

    \I__1884\ : ClkMux
    port map (
            O => \N__8656\,
            I => \N__8579\
        );

    \I__1883\ : ClkMux
    port map (
            O => \N__8655\,
            I => \N__8579\
        );

    \I__1882\ : ClkMux
    port map (
            O => \N__8654\,
            I => \N__8579\
        );

    \I__1881\ : GlobalMux
    port map (
            O => \N__8579\,
            I => \CLK80_PLL\
        );

    \I__1880\ : CEMux
    port map (
            O => \N__8576\,
            I => \N__8573\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__8573\,
            I => \N__8567\
        );

    \I__1878\ : CEMux
    port map (
            O => \N__8572\,
            I => \N__8564\
        );

    \I__1877\ : CEMux
    port map (
            O => \N__8571\,
            I => \N__8560\
        );

    \I__1876\ : CEMux
    port map (
            O => \N__8570\,
            I => \N__8557\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__8567\,
            I => \N__8554\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__8564\,
            I => \N__8551\
        );

    \I__1873\ : CEMux
    port map (
            O => \N__8563\,
            I => \N__8548\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8560\,
            I => \N__8543\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8557\,
            I => \N__8540\
        );

    \I__1870\ : Span4Mux_h
    port map (
            O => \N__8554\,
            I => \N__8533\
        );

    \I__1869\ : Span4Mux_h
    port map (
            O => \N__8551\,
            I => \N__8533\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8548\,
            I => \N__8533\
        );

    \I__1867\ : CEMux
    port map (
            O => \N__8547\,
            I => \N__8530\
        );

    \I__1866\ : CEMux
    port map (
            O => \N__8546\,
            I => \N__8527\
        );

    \I__1865\ : Span4Mux_v
    port map (
            O => \N__8543\,
            I => \N__8522\
        );

    \I__1864\ : Span4Mux_v
    port map (
            O => \N__8540\,
            I => \N__8522\
        );

    \I__1863\ : Span4Mux_v
    port map (
            O => \N__8533\,
            I => \N__8517\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8530\,
            I => \N__8517\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8527\,
            I => \N__8514\
        );

    \I__1860\ : Span4Mux_h
    port map (
            O => \N__8522\,
            I => \N__8511\
        );

    \I__1859\ : Span4Mux_v
    port map (
            O => \N__8517\,
            I => \N__8508\
        );

    \I__1858\ : Odrv4
    port map (
            O => \N__8514\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__8511\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__8508\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__8501\,
            I => \N__8498\
        );

    \I__1854\ : InMux
    port map (
            O => \N__8498\,
            I => \N__8492\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8497\,
            I => \N__8492\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__8492\,
            I => \N__8489\
        );

    \I__1851\ : Span4Mux_v
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__8486\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1849\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8475\
        );

    \I__1848\ : InMux
    port map (
            O => \N__8482\,
            I => \N__8475\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8481\,
            I => \N__8472\
        );

    \I__1846\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8469\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8475\,
            I => \N__8462\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__8472\,
            I => \N__8462\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__8469\,
            I => \N__8462\
        );

    \I__1842\ : Span4Mux_v
    port map (
            O => \N__8462\,
            I => \N__8459\
        );

    \I__1841\ : Span4Mux_v
    port map (
            O => \N__8459\,
            I => \N__8456\
        );

    \I__1840\ : Sp12to4
    port map (
            O => \N__8456\,
            I => \N__8453\
        );

    \I__1839\ : Span12Mux_h
    port map (
            O => \N__8453\,
            I => \N__8450\
        );

    \I__1838\ : Odrv12
    port map (
            O => \N__8450\,
            I => \DRA_c_3\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__8447\,
            I => \N__8444\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8441\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8441\,
            I => \N__8438\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__8438\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8435\,
            I => \N__8432\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8432\,
            I => \N__8429\
        );

    \I__1831\ : Span4Mux_h
    port map (
            O => \N__8429\,
            I => \N__8426\
        );

    \I__1830\ : Odrv4
    port map (
            O => \N__8426\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8420\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__8420\,
            I => \N__8417\
        );

    \I__1827\ : Odrv4
    port map (
            O => \N__8417\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1826\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8409\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8413\,
            I => \N__8406\
        );

    \I__1824\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8403\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8409\,
            I => \N__8399\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__8406\,
            I => \N__8396\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8403\,
            I => \N__8393\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8402\,
            I => \N__8390\
        );

    \I__1819\ : Span4Mux_v
    port map (
            O => \N__8399\,
            I => \N__8387\
        );

    \I__1818\ : Span4Mux_h
    port map (
            O => \N__8396\,
            I => \N__8380\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__8393\,
            I => \N__8380\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8390\,
            I => \N__8380\
        );

    \I__1815\ : Sp12to4
    port map (
            O => \N__8387\,
            I => \N__8377\
        );

    \I__1814\ : Sp12to4
    port map (
            O => \N__8380\,
            I => \N__8374\
        );

    \I__1813\ : Span12Mux_h
    port map (
            O => \N__8377\,
            I => \N__8371\
        );

    \I__1812\ : Span12Mux_v
    port map (
            O => \N__8374\,
            I => \N__8368\
        );

    \I__1811\ : Span12Mux_v
    port map (
            O => \N__8371\,
            I => \N__8365\
        );

    \I__1810\ : Span12Mux_h
    port map (
            O => \N__8368\,
            I => \N__8362\
        );

    \I__1809\ : Odrv12
    port map (
            O => \N__8365\,
            I => \DRA_c_2\
        );

    \I__1808\ : Odrv12
    port map (
            O => \N__8362\,
            I => \DRA_c_2\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8354\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__8354\,
            I => \N__8351\
        );

    \I__1805\ : Odrv4
    port map (
            O => \N__8351\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8348\,
            I => \N__8345\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8345\,
            I => \N__8342\
        );

    \I__1802\ : Span4Mux_h
    port map (
            O => \N__8342\,
            I => \N__8338\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8341\,
            I => \N__8335\
        );

    \I__1800\ : Odrv4
    port map (
            O => \N__8338\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8335\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0\
        );

    \I__1798\ : IoInMux
    port map (
            O => \N__8330\,
            I => \N__8327\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8327\,
            I => \N__8324\
        );

    \I__1796\ : Span4Mux_s3_h
    port map (
            O => \N__8324\,
            I => \N__8321\
        );

    \I__1795\ : Sp12to4
    port map (
            O => \N__8321\,
            I => \N__8318\
        );

    \I__1794\ : Span12Mux_v
    port map (
            O => \N__8318\,
            I => \N__8315\
        );

    \I__1793\ : Span12Mux_h
    port map (
            O => \N__8315\,
            I => \N__8312\
        );

    \I__1792\ : Odrv12
    port map (
            O => \N__8312\,
            I => \N_53_i\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8309\,
            I => \N__8306\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8306\,
            I => \U712_BYTE_ENABLE.N_303\
        );

    \I__1789\ : IoInMux
    port map (
            O => \N__8303\,
            I => \N__8300\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8300\,
            I => \N__8297\
        );

    \I__1787\ : Span4Mux_s3_v
    port map (
            O => \N__8297\,
            I => \N__8294\
        );

    \I__1786\ : Span4Mux_h
    port map (
            O => \N__8294\,
            I => \N__8291\
        );

    \I__1785\ : Span4Mux_h
    port map (
            O => \N__8291\,
            I => \N__8288\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__8288\,
            I => \UMBE_0_o2_i\
        );

    \I__1783\ : IoInMux
    port map (
            O => \N__8285\,
            I => \N__8282\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8282\,
            I => \N__8279\
        );

    \I__1781\ : Span4Mux_s2_v
    port map (
            O => \N__8279\,
            I => \N__8276\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__8276\,
            I => \N__8273\
        );

    \I__1779\ : Odrv4
    port map (
            O => \N__8273\,
            I => \U712_BYTE_ENABLE_UUBE_i\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8270\,
            I => \N__8266\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8269\,
            I => \N__8263\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__8266\,
            I => \N__8257\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__8263\,
            I => \N__8254\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8262\,
            I => \N__8251\
        );

    \I__1773\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8248\
        );

    \I__1772\ : InMux
    port map (
            O => \N__8260\,
            I => \N__8244\
        );

    \I__1771\ : Span4Mux_v
    port map (
            O => \N__8257\,
            I => \N__8235\
        );

    \I__1770\ : Span4Mux_h
    port map (
            O => \N__8254\,
            I => \N__8235\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__8251\,
            I => \N__8235\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8248\,
            I => \N__8235\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8247\,
            I => \N__8232\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__8244\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__8235\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8232\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1763\ : CascadeMux
    port map (
            O => \N__8225\,
            I => \N__8220\
        );

    \I__1762\ : CascadeMux
    port map (
            O => \N__8224\,
            I => \N__8216\
        );

    \I__1761\ : InMux
    port map (
            O => \N__8223\,
            I => \N__8213\
        );

    \I__1760\ : InMux
    port map (
            O => \N__8220\,
            I => \N__8210\
        );

    \I__1759\ : InMux
    port map (
            O => \N__8219\,
            I => \N__8205\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8216\,
            I => \N__8205\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__8213\,
            I => \N__8201\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8210\,
            I => \N__8195\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__8205\,
            I => \N__8195\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8204\,
            I => \N__8192\
        );

    \I__1753\ : Span4Mux_h
    port map (
            O => \N__8201\,
            I => \N__8189\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8186\
        );

    \I__1751\ : Span4Mux_h
    port map (
            O => \N__8195\,
            I => \N__8181\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__8192\,
            I => \N__8181\
        );

    \I__1749\ : Odrv4
    port map (
            O => \N__8189\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8186\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__8181\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8174\,
            I => \N__8170\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8173\,
            I => \N__8167\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__8170\,
            I => \N__8162\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8167\,
            I => \N__8159\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8166\,
            I => \N__8156\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__8165\,
            I => \N__8153\
        );

    \I__1740\ : Span4Mux_v
    port map (
            O => \N__8162\,
            I => \N__8146\
        );

    \I__1739\ : Span4Mux_h
    port map (
            O => \N__8159\,
            I => \N__8146\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8156\,
            I => \N__8146\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8153\,
            I => \N__8143\
        );

    \I__1736\ : Odrv4
    port map (
            O => \N__8146\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8143\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1734\ : IoInMux
    port map (
            O => \N__8138\,
            I => \N__8135\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8135\,
            I => \N__8132\
        );

    \I__1732\ : Span4Mux_s3_v
    port map (
            O => \N__8132\,
            I => \N__8129\
        );

    \I__1731\ : Sp12to4
    port map (
            O => \N__8129\,
            I => \N__8126\
        );

    \I__1730\ : Span12Mux_h
    port map (
            O => \N__8126\,
            I => \N__8123\
        );

    \I__1729\ : Odrv12
    port map (
            O => \N__8123\,
            I => \CMA_c_10\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8120\,
            I => \N__8117\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__8117\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8114\,
            I => \N__8111\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8111\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8105\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8105\,
            I => \N__8102\
        );

    \I__1722\ : Odrv4
    port map (
            O => \N__8102\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8096\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8096\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1719\ : IoInMux
    port map (
            O => \N__8093\,
            I => \N__8090\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__8090\,
            I => \N__8087\
        );

    \I__1717\ : Span12Mux_s11_v
    port map (
            O => \N__8087\,
            I => \N__8084\
        );

    \I__1716\ : Odrv12
    port map (
            O => \N__8084\,
            I => \CMA_c_2\
        );

    \I__1715\ : IoInMux
    port map (
            O => \N__8081\,
            I => \N__8078\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8078\,
            I => \N__8075\
        );

    \I__1713\ : Span4Mux_s3_h
    port map (
            O => \N__8075\,
            I => \N__8072\
        );

    \I__1712\ : Sp12to4
    port map (
            O => \N__8072\,
            I => \N__8069\
        );

    \I__1711\ : Span12Mux_s6_v
    port map (
            O => \N__8069\,
            I => \N__8066\
        );

    \I__1710\ : Span12Mux_h
    port map (
            O => \N__8066\,
            I => \N__8063\
        );

    \I__1709\ : Odrv12
    port map (
            O => \N__8063\,
            I => \CMA_c_3\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8060\,
            I => \N__8057\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__8057\,
            I => \N__8054\
        );

    \I__1706\ : Odrv4
    port map (
            O => \N__8054\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8051\,
            I => \N__8048\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__8048\,
            I => \N__8045\
        );

    \I__1703\ : Span4Mux_h
    port map (
            O => \N__8045\,
            I => \N__8042\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__8042\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8039\,
            I => \N__8036\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8036\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8033\,
            I => \N__8027\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8032\,
            I => \N__8027\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__8027\,
            I => \N__8024\
        );

    \I__1696\ : Span4Mux_h
    port map (
            O => \N__8024\,
            I => \N__8021\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__8021\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__8012\,
            I => \N__8009\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__8009\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1690\ : InMux
    port map (
            O => \N__8006\,
            I => \N__8003\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__8003\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1688\ : InMux
    port map (
            O => \N__8000\,
            I => \N__7996\
        );

    \I__1687\ : InMux
    port map (
            O => \N__7999\,
            I => \N__7993\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__7996\,
            I => \N__7990\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__7993\,
            I => \N__7987\
        );

    \I__1684\ : Odrv12
    port map (
            O => \N__7990\,
            I => \DBRn_c_i\
        );

    \I__1683\ : Odrv12
    port map (
            O => \N__7987\,
            I => \DBRn_c_i\
        );

    \I__1682\ : InMux
    port map (
            O => \N__7982\,
            I => \N__7979\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__7979\,
            I => \N__7976\
        );

    \I__1680\ : Span4Mux_h
    port map (
            O => \N__7976\,
            I => \N__7972\
        );

    \I__1679\ : InMux
    port map (
            O => \N__7975\,
            I => \N__7969\
        );

    \I__1678\ : Span4Mux_h
    port map (
            O => \N__7972\,
            I => \N__7966\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__7969\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__7966\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__1675\ : InMux
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__7958\,
            I => \N__7954\
        );

    \I__1673\ : InMux
    port map (
            O => \N__7957\,
            I => \N__7951\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__7954\,
            I => \U712_BYTE_ENABLE.N_370\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__7951\,
            I => \U712_BYTE_ENABLE.N_370\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__7946\,
            I => \U712_BYTE_ENABLE.N_369_cascade_\
        );

    \I__1669\ : IoInMux
    port map (
            O => \N__7943\,
            I => \N__7940\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__7940\,
            I => \N__7937\
        );

    \I__1667\ : Span4Mux_s0_h
    port map (
            O => \N__7937\,
            I => \N__7934\
        );

    \I__1666\ : Span4Mux_h
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__1665\ : Sp12to4
    port map (
            O => \N__7931\,
            I => \N__7928\
        );

    \I__1664\ : Span12Mux_s11_v
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__1663\ : Span12Mux_h
    port map (
            O => \N__7925\,
            I => \N__7922\
        );

    \I__1662\ : Odrv12
    port map (
            O => \N__7922\,
            I => \N_55_i\
        );

    \I__1661\ : IoInMux
    port map (
            O => \N__7919\,
            I => \N__7916\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7916\,
            I => \N__7913\
        );

    \I__1659\ : Span4Mux_s3_h
    port map (
            O => \N__7913\,
            I => \N__7910\
        );

    \I__1658\ : Sp12to4
    port map (
            O => \N__7910\,
            I => \N__7907\
        );

    \I__1657\ : Span12Mux_s6_v
    port map (
            O => \N__7907\,
            I => \N__7904\
        );

    \I__1656\ : Odrv12
    port map (
            O => \N__7904\,
            I => \WEn_c\
        );

    \I__1655\ : IoInMux
    port map (
            O => \N__7901\,
            I => \N__7898\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__7898\,
            I => \N__7895\
        );

    \I__1653\ : Span4Mux_s3_v
    port map (
            O => \N__7895\,
            I => \N__7892\
        );

    \I__1652\ : Span4Mux_v
    port map (
            O => \N__7892\,
            I => \N__7889\
        );

    \I__1651\ : Span4Mux_h
    port map (
            O => \N__7889\,
            I => \N__7886\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__7886\,
            I => \CRCSn_c\
        );

    \I__1649\ : IoInMux
    port map (
            O => \N__7883\,
            I => \N__7880\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__7880\,
            I => \N__7877\
        );

    \I__1647\ : Span4Mux_s2_v
    port map (
            O => \N__7877\,
            I => \N__7874\
        );

    \I__1646\ : Sp12to4
    port map (
            O => \N__7874\,
            I => \N__7871\
        );

    \I__1645\ : Span12Mux_h
    port map (
            O => \N__7871\,
            I => \N__7868\
        );

    \I__1644\ : Odrv12
    port map (
            O => \N__7868\,
            I => \RASn_c\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__7865\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\
        );

    \I__1642\ : InMux
    port map (
            O => \N__7862\,
            I => \N__7859\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7859\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1640\ : InMux
    port map (
            O => \N__7856\,
            I => \N__7853\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__7853\,
            I => \N__7850\
        );

    \I__1638\ : Span4Mux_h
    port map (
            O => \N__7850\,
            I => \N__7847\
        );

    \I__1637\ : Odrv4
    port map (
            O => \N__7847\,
            I => \U712_CHIP_RAM.N_392\
        );

    \I__1636\ : InMux
    port map (
            O => \N__7844\,
            I => \N__7841\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__7841\,
            I => \N__7838\
        );

    \I__1634\ : Span12Mux_h
    port map (
            O => \N__7838\,
            I => \N__7835\
        );

    \I__1633\ : Odrv12
    port map (
            O => \N__7835\,
            I => \A_c_13\
        );

    \I__1632\ : InMux
    port map (
            O => \N__7832\,
            I => \N__7829\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__1630\ : Span4Mux_v
    port map (
            O => \N__7826\,
            I => \N__7823\
        );

    \I__1629\ : Span4Mux_v
    port map (
            O => \N__7823\,
            I => \N__7820\
        );

    \I__1628\ : Sp12to4
    port map (
            O => \N__7820\,
            I => \N__7817\
        );

    \I__1627\ : Span12Mux_h
    port map (
            O => \N__7817\,
            I => \N__7814\
        );

    \I__1626\ : Odrv12
    port map (
            O => \N__7814\,
            I => \A_c_6\
        );

    \I__1625\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7805\
        );

    \I__1624\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7805\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7805\,
            I => \N__7802\
        );

    \I__1622\ : Span4Mux_v
    port map (
            O => \N__7802\,
            I => \N__7799\
        );

    \I__1621\ : Span4Mux_v
    port map (
            O => \N__7799\,
            I => \N__7796\
        );

    \I__1620\ : Sp12to4
    port map (
            O => \N__7796\,
            I => \N__7793\
        );

    \I__1619\ : Span12Mux_h
    port map (
            O => \N__7793\,
            I => \N__7790\
        );

    \I__1618\ : Odrv12
    port map (
            O => \N__7790\,
            I => \A_c_14\
        );

    \I__1617\ : InMux
    port map (
            O => \N__7787\,
            I => \N__7784\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__7784\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1615\ : InMux
    port map (
            O => \N__7781\,
            I => \N__7778\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__7778\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1613\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7772\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__7772\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__1611\ : IoInMux
    port map (
            O => \N__7769\,
            I => \N__7766\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__7766\,
            I => \N__7763\
        );

    \I__1609\ : IoSpan4Mux
    port map (
            O => \N__7763\,
            I => \N__7760\
        );

    \I__1608\ : Span4Mux_s2_h
    port map (
            O => \N__7760\,
            I => \N__7757\
        );

    \I__1607\ : Sp12to4
    port map (
            O => \N__7757\,
            I => \N__7754\
        );

    \I__1606\ : Span12Mux_h
    port map (
            O => \N__7754\,
            I => \N__7751\
        );

    \I__1605\ : Odrv12
    port map (
            O => \N__7751\,
            I => \CMA_c_5\
        );

    \I__1604\ : InMux
    port map (
            O => \N__7748\,
            I => \N__7745\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__7745\,
            I => \N__7742\
        );

    \I__1602\ : Span12Mux_v
    port map (
            O => \N__7742\,
            I => \N__7739\
        );

    \I__1601\ : Span12Mux_h
    port map (
            O => \N__7739\,
            I => \N__7736\
        );

    \I__1600\ : Odrv12
    port map (
            O => \N__7736\,
            I => \A_c_11\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7730\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__7730\,
            I => \N__7727\
        );

    \I__1597\ : Span4Mux_v
    port map (
            O => \N__7727\,
            I => \N__7724\
        );

    \I__1596\ : Span4Mux_v
    port map (
            O => \N__7724\,
            I => \N__7721\
        );

    \I__1595\ : Sp12to4
    port map (
            O => \N__7721\,
            I => \N__7718\
        );

    \I__1594\ : Span12Mux_h
    port map (
            O => \N__7718\,
            I => \N__7715\
        );

    \I__1593\ : Odrv12
    port map (
            O => \N__7715\,
            I => \A_c_4\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__7712\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7709\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7706\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__1589\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7699\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7702\,
            I => \N__7696\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__7699\,
            I => \N__7684\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__7696\,
            I => \N__7681\
        );

    \I__1585\ : ClkMux
    port map (
            O => \N__7695\,
            I => \N__7658\
        );

    \I__1584\ : ClkMux
    port map (
            O => \N__7694\,
            I => \N__7658\
        );

    \I__1583\ : ClkMux
    port map (
            O => \N__7693\,
            I => \N__7658\
        );

    \I__1582\ : ClkMux
    port map (
            O => \N__7692\,
            I => \N__7658\
        );

    \I__1581\ : ClkMux
    port map (
            O => \N__7691\,
            I => \N__7658\
        );

    \I__1580\ : ClkMux
    port map (
            O => \N__7690\,
            I => \N__7658\
        );

    \I__1579\ : ClkMux
    port map (
            O => \N__7689\,
            I => \N__7658\
        );

    \I__1578\ : ClkMux
    port map (
            O => \N__7688\,
            I => \N__7658\
        );

    \I__1577\ : ClkMux
    port map (
            O => \N__7687\,
            I => \N__7658\
        );

    \I__1576\ : Glb2LocalMux
    port map (
            O => \N__7684\,
            I => \N__7658\
        );

    \I__1575\ : Glb2LocalMux
    port map (
            O => \N__7681\,
            I => \N__7658\
        );

    \I__1574\ : GlobalMux
    port map (
            O => \N__7658\,
            I => \N__7655\
        );

    \I__1573\ : gio2CtrlBuf
    port map (
            O => \N__7655\,
            I => \C1_c_g\
        );

    \I__1572\ : SRMux
    port map (
            O => \N__7652\,
            I => \N__7649\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__7649\,
            I => \N__7646\
        );

    \I__1570\ : Span4Mux_v
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__1569\ : Odrv4
    port map (
            O => \N__7643\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7636\
        );

    \I__1567\ : InMux
    port map (
            O => \N__7639\,
            I => \N__7633\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7636\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__7633\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7628\,
            I => \N__7624\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7627\,
            I => \N__7621\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__7624\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7621\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7616\,
            I => \N__7612\
        );

    \I__1559\ : InMux
    port map (
            O => \N__7615\,
            I => \N__7609\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7612\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7609\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7604\,
            I => \N__7601\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7601\,
            I => \N__7598\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__7598\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7595\,
            I => \N__7591\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7594\,
            I => \N__7588\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7591\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7588\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7583\,
            I => \N__7579\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7582\,
            I => \N__7576\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7579\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__7576\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__1545\ : CascadeMux
    port map (
            O => \N__7571\,
            I => \N__7567\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7564\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7567\,
            I => \N__7561\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__7564\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__7561\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7556\,
            I => \N__7552\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7555\,
            I => \N__7549\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7552\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__7549\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__1536\ : InMux
    port map (
            O => \N__7544\,
            I => \N__7541\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__7541\,
            I => \N__7538\
        );

    \I__1534\ : Odrv4
    port map (
            O => \N__7538\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__7535\,
            I => \N__7523\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__7534\,
            I => \N__7512\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7533\,
            I => \N__7509\
        );

    \I__1530\ : InMux
    port map (
            O => \N__7532\,
            I => \N__7506\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7531\,
            I => \N__7499\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7530\,
            I => \N__7499\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7529\,
            I => \N__7499\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7528\,
            I => \N__7496\
        );

    \I__1525\ : InMux
    port map (
            O => \N__7527\,
            I => \N__7492\
        );

    \I__1524\ : InMux
    port map (
            O => \N__7526\,
            I => \N__7485\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7485\
        );

    \I__1522\ : InMux
    port map (
            O => \N__7522\,
            I => \N__7485\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7521\,
            I => \N__7482\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__7520\,
            I => \N__7478\
        );

    \I__1519\ : InMux
    port map (
            O => \N__7519\,
            I => \N__7471\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7518\,
            I => \N__7471\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7517\,
            I => \N__7468\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7463\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7515\,
            I => \N__7463\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7460\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7509\,
            I => \N__7457\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__7506\,
            I => \N__7450\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7499\,
            I => \N__7450\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7496\,
            I => \N__7450\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7495\,
            I => \N__7447\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7492\,
            I => \N__7442\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7485\,
            I => \N__7437\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7482\,
            I => \N__7437\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7481\,
            I => \N__7432\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7478\,
            I => \N__7432\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7477\,
            I => \N__7429\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7476\,
            I => \N__7426\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7471\,
            I => \N__7421\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7468\,
            I => \N__7421\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__7463\,
            I => \N__7416\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7460\,
            I => \N__7416\
        );

    \I__1497\ : Span4Mux_v
    port map (
            O => \N__7457\,
            I => \N__7409\
        );

    \I__1496\ : Span4Mux_v
    port map (
            O => \N__7450\,
            I => \N__7409\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7447\,
            I => \N__7409\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7446\,
            I => \N__7404\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7445\,
            I => \N__7404\
        );

    \I__1492\ : Span4Mux_v
    port map (
            O => \N__7442\,
            I => \N__7393\
        );

    \I__1491\ : Span4Mux_v
    port map (
            O => \N__7437\,
            I => \N__7393\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__7432\,
            I => \N__7393\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7429\,
            I => \N__7393\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7426\,
            I => \N__7393\
        );

    \I__1487\ : Span4Mux_v
    port map (
            O => \N__7421\,
            I => \N__7384\
        );

    \I__1486\ : Span4Mux_h
    port map (
            O => \N__7416\,
            I => \N__7384\
        );

    \I__1485\ : Span4Mux_h
    port map (
            O => \N__7409\,
            I => \N__7384\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7404\,
            I => \N__7384\
        );

    \I__1483\ : Span4Mux_v
    port map (
            O => \N__7393\,
            I => \N__7378\
        );

    \I__1482\ : Span4Mux_v
    port map (
            O => \N__7384\,
            I => \N__7375\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7383\,
            I => \N__7372\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7382\,
            I => \N__7369\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7381\,
            I => \N__7366\
        );

    \I__1478\ : Sp12to4
    port map (
            O => \N__7378\,
            I => \N__7355\
        );

    \I__1477\ : Sp12to4
    port map (
            O => \N__7375\,
            I => \N__7355\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7372\,
            I => \N__7355\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__7369\,
            I => \N__7355\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7366\,
            I => \N__7355\
        );

    \I__1473\ : Span12Mux_h
    port map (
            O => \N__7355\,
            I => \N__7352\
        );

    \I__1472\ : Odrv12
    port map (
            O => \N__7352\,
            I => \RESETn_c\
        );

    \I__1471\ : IoInMux
    port map (
            O => \N__7349\,
            I => \N__7346\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7346\,
            I => \N__7343\
        );

    \I__1469\ : IoSpan4Mux
    port map (
            O => \N__7343\,
            I => \N__7340\
        );

    \I__1468\ : Span4Mux_s3_v
    port map (
            O => \N__7340\,
            I => \N__7336\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7339\,
            I => \N__7333\
        );

    \I__1466\ : Span4Mux_v
    port map (
            O => \N__7336\,
            I => \N__7330\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7333\,
            I => \N__7327\
        );

    \I__1464\ : Span4Mux_v
    port map (
            O => \N__7330\,
            I => \N__7324\
        );

    \I__1463\ : Span4Mux_h
    port map (
            O => \N__7327\,
            I => \N__7321\
        );

    \I__1462\ : Span4Mux_v
    port map (
            O => \N__7324\,
            I => \N__7316\
        );

    \I__1461\ : Span4Mux_v
    port map (
            O => \N__7321\,
            I => \N__7316\
        );

    \I__1460\ : Odrv4
    port map (
            O => \N__7316\,
            I => \RESETn_c_i\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7313\,
            I => \N__7310\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7310\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__1457\ : IoInMux
    port map (
            O => \N__7307\,
            I => \N__7304\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7304\,
            I => \N__7301\
        );

    \I__1455\ : Odrv12
    port map (
            O => \N__7301\,
            I => \CMA_c_1\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7298\,
            I => \N__7295\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7295\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7292\,
            I => \N__7289\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7289\,
            I => \N__7286\
        );

    \I__1450\ : Span4Mux_v
    port map (
            O => \N__7286\,
            I => \N__7283\
        );

    \I__1449\ : Span4Mux_v
    port map (
            O => \N__7283\,
            I => \N__7280\
        );

    \I__1448\ : Sp12to4
    port map (
            O => \N__7280\,
            I => \N__7277\
        );

    \I__1447\ : Span12Mux_h
    port map (
            O => \N__7277\,
            I => \N__7274\
        );

    \I__1446\ : Odrv12
    port map (
            O => \N__7274\,
            I => \A_c_16\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7268\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__7268\,
            I => \N__7265\
        );

    \I__1443\ : Span4Mux_v
    port map (
            O => \N__7265\,
            I => \N__7262\
        );

    \I__1442\ : Span4Mux_v
    port map (
            O => \N__7262\,
            I => \N__7259\
        );

    \I__1441\ : Sp12to4
    port map (
            O => \N__7259\,
            I => \N__7256\
        );

    \I__1440\ : Span12Mux_h
    port map (
            O => \N__7256\,
            I => \N__7253\
        );

    \I__1439\ : Odrv12
    port map (
            O => \N__7253\,
            I => \A_c_18\
        );

    \I__1438\ : CascadeMux
    port map (
            O => \N__7250\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7247\,
            I => \N__7244\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7244\,
            I => \U712_CHIP_RAM.CLK_EN_5_0_a2_0\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__7241\,
            I => \N__7238\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7235\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7235\,
            I => \U712_CHIP_RAM.N_112\
        );

    \I__1432\ : IoInMux
    port map (
            O => \N__7232\,
            I => \N__7229\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__7229\,
            I => \N__7226\
        );

    \I__1430\ : IoSpan4Mux
    port map (
            O => \N__7226\,
            I => \N__7223\
        );

    \I__1429\ : IoSpan4Mux
    port map (
            O => \N__7223\,
            I => \N__7220\
        );

    \I__1428\ : Span4Mux_s2_h
    port map (
            O => \N__7220\,
            I => \N__7217\
        );

    \I__1427\ : Sp12to4
    port map (
            O => \N__7217\,
            I => \N__7214\
        );

    \I__1426\ : Span12Mux_s9_h
    port map (
            O => \N__7214\,
            I => \N__7210\
        );

    \I__1425\ : InMux
    port map (
            O => \N__7213\,
            I => \N__7207\
        );

    \I__1424\ : Odrv12
    port map (
            O => \N__7210\,
            I => \CLK_EN_c\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__7207\,
            I => \CLK_EN_c\
        );

    \I__1422\ : InMux
    port map (
            O => \N__7202\,
            I => \bfn_11_7_0_\
        );

    \I__1421\ : InMux
    port map (
            O => \N__7199\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7196\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7190\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__7190\,
            I => \N__7186\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7183\
        );

    \I__1416\ : Span4Mux_h
    port map (
            O => \N__7186\,
            I => \N__7180\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__7183\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__7180\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7175\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7172\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7169\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__7166\,
            I => \N__7161\
        );

    \I__1409\ : CascadeMux
    port map (
            O => \N__7165\,
            I => \N__7156\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7164\,
            I => \N__7148\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7161\,
            I => \N__7148\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7160\,
            I => \N__7148\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7159\,
            I => \N__7141\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7141\
        );

    \I__1403\ : InMux
    port map (
            O => \N__7155\,
            I => \N__7141\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__7148\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7141\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7133\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7133\,
            I => \U712_REG_SM.m17_i_0_o2_1\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__7130\,
            I => \N__7127\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7127\,
            I => \N__7124\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7124\,
            I => \U712_REG_SM.N_435\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__7121\,
            I => \U712_REG_SM.N_435_cascade_\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7115\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7115\,
            I => \U712_REG_SM.N_363\
        );

    \I__1392\ : IoInMux
    port map (
            O => \N__7112\,
            I => \N__7108\
        );

    \I__1391\ : IoInMux
    port map (
            O => \N__7111\,
            I => \N__7105\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7108\,
            I => \N__7102\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__7105\,
            I => \N__7099\
        );

    \I__1388\ : Span4Mux_s0_v
    port map (
            O => \N__7102\,
            I => \N__7096\
        );

    \I__1387\ : Span4Mux_s0_v
    port map (
            O => \N__7099\,
            I => \N__7093\
        );

    \I__1386\ : Span4Mux_v
    port map (
            O => \N__7096\,
            I => \N__7090\
        );

    \I__1385\ : Span4Mux_v
    port map (
            O => \N__7093\,
            I => \N__7087\
        );

    \I__1384\ : Sp12to4
    port map (
            O => \N__7090\,
            I => \N__7084\
        );

    \I__1383\ : Sp12to4
    port map (
            O => \N__7087\,
            I => \N__7081\
        );

    \I__1382\ : Span12Mux_s10_h
    port map (
            O => \N__7084\,
            I => \N__7078\
        );

    \I__1381\ : Span12Mux_s9_h
    port map (
            O => \N__7081\,
            I => \N__7075\
        );

    \I__1380\ : Span12Mux_v
    port map (
            O => \N__7078\,
            I => \N__7069\
        );

    \I__1379\ : Span12Mux_v
    port map (
            O => \N__7075\,
            I => \N__7069\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7074\,
            I => \N__7066\
        );

    \I__1377\ : Odrv12
    port map (
            O => \N__7069\,
            I => \ASn_c\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__7066\,
            I => \ASn_c\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7061\,
            I => \N__7055\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7060\,
            I => \N__7055\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__7055\,
            I => \U712_REG_SM.ASn_0_sqmuxa\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__7052\,
            I => \N__7048\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__7051\,
            I => \N__7045\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7048\,
            I => \N__7031\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7045\,
            I => \N__7031\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7044\,
            I => \N__7022\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7043\,
            I => \N__7022\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7042\,
            I => \N__7022\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7022\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7040\,
            I => \N__7013\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7039\,
            I => \N__7013\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7038\,
            I => \N__7013\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7037\,
            I => \N__7013\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7036\,
            I => \N__7010\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7031\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__7022\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7013\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7010\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7001\,
            I => \N__6993\
        );

    \I__1354\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6993\
        );

    \I__1353\ : InMux
    port map (
            O => \N__6999\,
            I => \N__6990\
        );

    \I__1352\ : InMux
    port map (
            O => \N__6998\,
            I => \N__6987\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6993\,
            I => \U712_REG_SM.m17_i_0_o2\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6990\,
            I => \U712_REG_SM.m17_i_0_o2\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6987\,
            I => \U712_REG_SM.m17_i_0_o2\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6980\,
            I => \N__6973\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6979\,
            I => \N__6968\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6978\,
            I => \N__6968\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6963\
        );

    \I__1344\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6963\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__6973\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6968\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__6963\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__6956\,
            I => \N__6953\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6953\,
            I => \N__6945\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6952\,
            I => \N__6945\
        );

    \I__1337\ : InMux
    port map (
            O => \N__6951\,
            I => \N__6940\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6950\,
            I => \N__6940\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__6945\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__6940\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1333\ : InMux
    port map (
            O => \N__6935\,
            I => \N__6931\
        );

    \I__1332\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6927\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__6931\,
            I => \N__6924\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6930\,
            I => \N__6921\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6927\,
            I => \N__6916\
        );

    \I__1328\ : Span4Mux_v
    port map (
            O => \N__6924\,
            I => \N__6916\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__6921\,
            I => \N__6913\
        );

    \I__1326\ : Sp12to4
    port map (
            O => \N__6916\,
            I => \N__6910\
        );

    \I__1325\ : Span4Mux_v
    port map (
            O => \N__6913\,
            I => \N__6907\
        );

    \I__1324\ : Span12Mux_h
    port map (
            O => \N__6910\,
            I => \N__6904\
        );

    \I__1323\ : Sp12to4
    port map (
            O => \N__6907\,
            I => \N__6901\
        );

    \I__1322\ : Span12Mux_v
    port map (
            O => \N__6904\,
            I => \N__6896\
        );

    \I__1321\ : Span12Mux_h
    port map (
            O => \N__6901\,
            I => \N__6896\
        );

    \I__1320\ : Odrv12
    port map (
            O => \N__6896\,
            I => \RnW_c\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6888\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6892\,
            I => \N__6885\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__6891\,
            I => \N__6879\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6888\,
            I => \N__6874\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__6885\,
            I => \N__6874\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6884\,
            I => \N__6871\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6883\,
            I => \N__6868\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__6882\,
            I => \N__6864\
        );

    \I__1311\ : InMux
    port map (
            O => \N__6879\,
            I => \N__6861\
        );

    \I__1310\ : Span12Mux_h
    port map (
            O => \N__6874\,
            I => \N__6858\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6871\,
            I => \N__6852\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__6868\,
            I => \N__6852\
        );

    \I__1307\ : InMux
    port map (
            O => \N__6867\,
            I => \N__6849\
        );

    \I__1306\ : InMux
    port map (
            O => \N__6864\,
            I => \N__6843\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6861\,
            I => \N__6840\
        );

    \I__1304\ : Span12Mux_v
    port map (
            O => \N__6858\,
            I => \N__6837\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6857\,
            I => \N__6834\
        );

    \I__1302\ : Span4Mux_v
    port map (
            O => \N__6852\,
            I => \N__6829\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__6849\,
            I => \N__6829\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6826\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6847\,
            I => \N__6821\
        );

    \I__1298\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6821\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6843\,
            I => \N__6816\
        );

    \I__1296\ : Span4Mux_v
    port map (
            O => \N__6840\,
            I => \N__6816\
        );

    \I__1295\ : Odrv12
    port map (
            O => \N__6837\,
            I => \WRITE_CYCLEm\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6834\,
            I => \WRITE_CYCLEm\
        );

    \I__1293\ : Odrv4
    port map (
            O => \N__6829\,
            I => \WRITE_CYCLEm\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__6826\,
            I => \WRITE_CYCLEm\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__6821\,
            I => \WRITE_CYCLEm\
        );

    \I__1290\ : Odrv4
    port map (
            O => \N__6816\,
            I => \WRITE_CYCLEm\
        );

    \I__1289\ : IoInMux
    port map (
            O => \N__6803\,
            I => \N__6800\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6800\,
            I => \N__6797\
        );

    \I__1287\ : IoSpan4Mux
    port map (
            O => \N__6797\,
            I => \N__6794\
        );

    \I__1286\ : IoSpan4Mux
    port map (
            O => \N__6794\,
            I => \N__6791\
        );

    \I__1285\ : Sp12to4
    port map (
            O => \N__6791\,
            I => \N__6788\
        );

    \I__1284\ : Span12Mux_s7_h
    port map (
            O => \N__6788\,
            I => \N__6785\
        );

    \I__1283\ : Odrv12
    port map (
            O => \N__6785\,
            I => \N_276\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6779\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6779\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6770\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6767\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6758\
        );

    \I__1277\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6755\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__6770\,
            I => \N__6749\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6767\,
            I => \N__6746\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6766\,
            I => \N__6743\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6738\
        );

    \I__1272\ : InMux
    port map (
            O => \N__6764\,
            I => \N__6738\
        );

    \I__1271\ : InMux
    port map (
            O => \N__6763\,
            I => \N__6731\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6762\,
            I => \N__6731\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6761\,
            I => \N__6728\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6758\,
            I => \N__6725\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__6755\,
            I => \N__6715\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6754\,
            I => \N__6712\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6753\,
            I => \N__6709\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6752\,
            I => \N__6706\
        );

    \I__1263\ : Span4Mux_v
    port map (
            O => \N__6749\,
            I => \N__6699\
        );

    \I__1262\ : Span4Mux_v
    port map (
            O => \N__6746\,
            I => \N__6699\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__6743\,
            I => \N__6699\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6738\,
            I => \N__6696\
        );

    \I__1259\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6691\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6691\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6731\,
            I => \N__6684\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__6728\,
            I => \N__6684\
        );

    \I__1255\ : Span4Mux_h
    port map (
            O => \N__6725\,
            I => \N__6684\
        );

    \I__1254\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6681\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6678\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6722\,
            I => \N__6673\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6721\,
            I => \N__6673\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6666\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6666\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6718\,
            I => \N__6666\
        );

    \I__1247\ : Odrv4
    port map (
            O => \N__6715\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6712\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6709\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6706\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1243\ : Odrv4
    port map (
            O => \N__6699\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1242\ : Odrv4
    port map (
            O => \N__6696\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6691\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__6684\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__6681\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6678\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6673\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6666\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6641\,
            I => \N__6638\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6638\,
            I => \N__6635\
        );

    \I__1233\ : Span4Mux_h
    port map (
            O => \N__6635\,
            I => \N__6632\
        );

    \I__1232\ : Odrv4
    port map (
            O => \N__6632\,
            I => \U712_CHIP_RAM.N_300\
        );

    \I__1231\ : CascadeMux
    port map (
            O => \N__6629\,
            I => \N__6625\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__6628\,
            I => \N__6622\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6625\,
            I => \N__6615\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6622\,
            I => \N__6610\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6621\,
            I => \N__6610\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__6620\,
            I => \N__6605\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__6619\,
            I => \N__6597\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6618\,
            I => \N__6593\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6615\,
            I => \N__6589\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__6610\,
            I => \N__6586\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6609\,
            I => \N__6581\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6608\,
            I => \N__6576\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6605\,
            I => \N__6576\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6604\,
            I => \N__6571\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6603\,
            I => \N__6571\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__6602\,
            I => \N__6568\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__6601\,
            I => \N__6564\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6600\,
            I => \N__6561\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6597\,
            I => \N__6558\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6555\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6593\,
            I => \N__6552\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__6592\,
            I => \N__6545\
        );

    \I__1209\ : Span4Mux_v
    port map (
            O => \N__6589\,
            I => \N__6539\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__6586\,
            I => \N__6539\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6585\,
            I => \N__6536\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6584\,
            I => \N__6533\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6581\,
            I => \N__6528\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__6576\,
            I => \N__6528\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6571\,
            I => \N__6525\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6568\,
            I => \N__6522\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6567\,
            I => \N__6517\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6564\,
            I => \N__6517\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6561\,
            I => \N__6508\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6558\,
            I => \N__6508\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6555\,
            I => \N__6508\
        );

    \I__1196\ : Span4Mux_h
    port map (
            O => \N__6552\,
            I => \N__6508\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6551\,
            I => \N__6505\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6500\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6549\,
            I => \N__6500\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6548\,
            I => \N__6493\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6545\,
            I => \N__6493\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6544\,
            I => \N__6493\
        );

    \I__1189\ : Odrv4
    port map (
            O => \N__6539\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6536\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__6533\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1186\ : Odrv4
    port map (
            O => \N__6528\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1185\ : Odrv12
    port map (
            O => \N__6525\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6522\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6517\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1182\ : Odrv4
    port map (
            O => \N__6508\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6505\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6500\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6493\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6470\,
            I => \N__6461\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6469\,
            I => \N__6457\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__6468\,
            I => \N__6454\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__6467\,
            I => \N__6450\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6466\,
            I => \N__6447\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6465\,
            I => \N__6444\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6464\,
            I => \N__6439\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6461\,
            I => \N__6436\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6460\,
            I => \N__6432\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6457\,
            I => \N__6429\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6454\,
            I => \N__6426\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6453\,
            I => \N__6422\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6450\,
            I => \N__6419\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6447\,
            I => \N__6414\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__6444\,
            I => \N__6414\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6443\,
            I => \N__6411\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6442\,
            I => \N__6408\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__6439\,
            I => \N__6403\
        );

    \I__1160\ : Span4Mux_v
    port map (
            O => \N__6436\,
            I => \N__6403\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6435\,
            I => \N__6400\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6432\,
            I => \N__6393\
        );

    \I__1157\ : Span4Mux_h
    port map (
            O => \N__6429\,
            I => \N__6393\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6426\,
            I => \N__6393\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6425\,
            I => \N__6390\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6422\,
            I => \U712_CHIP_RAM.N_241\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6419\,
            I => \U712_CHIP_RAM.N_241\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__6414\,
            I => \U712_CHIP_RAM.N_241\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__6411\,
            I => \U712_CHIP_RAM.N_241\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6408\,
            I => \U712_CHIP_RAM.N_241\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__6403\,
            I => \U712_CHIP_RAM.N_241\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6400\,
            I => \U712_CHIP_RAM.N_241\
        );

    \I__1147\ : Odrv4
    port map (
            O => \N__6393\,
            I => \U712_CHIP_RAM.N_241\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6390\,
            I => \U712_CHIP_RAM.N_241\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__6371\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6356\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6353\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6366\,
            I => \N__6350\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6365\,
            I => \N__6345\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6364\,
            I => \N__6342\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6363\,
            I => \N__6339\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6362\,
            I => \N__6334\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6361\,
            I => \N__6334\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6360\,
            I => \N__6331\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6328\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6356\,
            I => \N__6323\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6353\,
            I => \N__6318\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6350\,
            I => \N__6318\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6315\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6312\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6345\,
            I => \N__6305\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6342\,
            I => \N__6305\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__6339\,
            I => \N__6300\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6334\,
            I => \N__6300\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6331\,
            I => \N__6295\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6328\,
            I => \N__6295\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6290\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6287\
        );

    \I__1121\ : Span4Mux_v
    port map (
            O => \N__6323\,
            I => \N__6284\
        );

    \I__1120\ : Span4Mux_h
    port map (
            O => \N__6318\,
            I => \N__6281\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6315\,
            I => \N__6276\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6312\,
            I => \N__6276\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6271\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6271\
        );

    \I__1115\ : Span4Mux_v
    port map (
            O => \N__6305\,
            I => \N__6264\
        );

    \I__1114\ : Span4Mux_h
    port map (
            O => \N__6300\,
            I => \N__6264\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__6295\,
            I => \N__6264\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6294\,
            I => \N__6259\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6259\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6290\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6287\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1108\ : Odrv4
    port map (
            O => \N__6284\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1107\ : Odrv4
    port map (
            O => \N__6281\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1106\ : Odrv4
    port map (
            O => \N__6276\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6271\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1104\ : Odrv4
    port map (
            O => \N__6264\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__6259\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6242\,
            I => \N__6239\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__6239\,
            I => \N__6236\
        );

    \I__1100\ : Span4Mux_v
    port map (
            O => \N__6236\,
            I => \N__6233\
        );

    \I__1099\ : Sp12to4
    port map (
            O => \N__6233\,
            I => \N__6230\
        );

    \I__1098\ : Span12Mux_h
    port map (
            O => \N__6230\,
            I => \N__6227\
        );

    \I__1097\ : Odrv12
    port map (
            O => \N__6227\,
            I => \A_c_9\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6224\,
            I => \N__6221\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__6221\,
            I => \N__6218\
        );

    \I__1094\ : Span4Mux_h
    port map (
            O => \N__6218\,
            I => \N__6215\
        );

    \I__1093\ : Sp12to4
    port map (
            O => \N__6215\,
            I => \N__6212\
        );

    \I__1092\ : Span12Mux_v
    port map (
            O => \N__6212\,
            I => \N__6209\
        );

    \I__1091\ : Odrv12
    port map (
            O => \N__6209\,
            I => \A_c_2\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6206\,
            I => \N__6202\
        );

    \I__1089\ : InMux
    port map (
            O => \N__6205\,
            I => \N__6198\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__6202\,
            I => \N__6195\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6192\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__6198\,
            I => \N__6189\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__6195\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__6192\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1083\ : Odrv4
    port map (
            O => \N__6189\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__6182\,
            I => \U712_REG_SM.N_360_1_cascade_\
        );

    \I__1081\ : CascadeMux
    port map (
            O => \N__6179\,
            I => \N__6175\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6178\,
            I => \N__6170\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6175\,
            I => \N__6170\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6170\,
            I => \U712_REG_SM.C3_SYNC_RNI7UAPZ0Z_1\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__6167\,
            I => \U712_REG_SM.m17_i_0_o2_cascade_\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__6164\,
            I => \U712_REG_SM.REG_CYCLE_RNOZ0Z_0_cascade_\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6158\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__6158\,
            I => \N__6152\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6149\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6156\,
            I => \N__6146\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6155\,
            I => \N__6143\
        );

    \I__1070\ : Odrv12
    port map (
            O => \N__6152\,
            I => \U712_CHIP_RAM.N_388\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6149\,
            I => \U712_CHIP_RAM.N_388\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6146\,
            I => \U712_CHIP_RAM.N_388\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__6143\,
            I => \U712_CHIP_RAM.N_388\
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__6134\,
            I => \N__6129\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6125\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6132\,
            I => \N__6122\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6129\,
            I => \N__6119\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__6128\,
            I => \N__6116\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__6125\,
            I => \N__6112\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6122\,
            I => \N__6107\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6119\,
            I => \N__6107\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6116\,
            I => \N__6102\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6115\,
            I => \N__6102\
        );

    \I__1056\ : Odrv4
    port map (
            O => \N__6112\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1055\ : Odrv4
    port map (
            O => \N__6107\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__6102\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6095\,
            I => \N__6089\
        );

    \I__1052\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6086\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6083\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__6092\,
            I => \N__6080\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6089\,
            I => \N__6073\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__6086\,
            I => \N__6073\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__6083\,
            I => \N__6070\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6080\,
            I => \N__6063\
        );

    \I__1045\ : InMux
    port map (
            O => \N__6079\,
            I => \N__6063\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6060\
        );

    \I__1043\ : Span4Mux_h
    port map (
            O => \N__6073\,
            I => \N__6055\
        );

    \I__1042\ : Span4Mux_h
    port map (
            O => \N__6070\,
            I => \N__6055\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6069\,
            I => \N__6050\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6068\,
            I => \N__6050\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__6063\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6060\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1037\ : Odrv4
    port map (
            O => \N__6055\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6050\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__6041\,
            I => \U712_CHIP_RAM.N_271_cascade_\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6035\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6035\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__6032\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1_1_cascade_\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6029\,
            I => \N__6026\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6026\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_2_1\
        );

    \I__1029\ : InMux
    port map (
            O => \N__6023\,
            I => \N__6020\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__6020\,
            I => \U712_CHIP_RAM.N_317\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__6017\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_0_cascade_\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6014\,
            I => \N__6010\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6013\,
            I => \N__6007\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__6010\,
            I => \U712_CHIP_RAM.N_434\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__6007\,
            I => \U712_CHIP_RAM.N_434\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6002\,
            I => \N__5999\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__5999\,
            I => \U712_CHIP_RAM.N_13\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5996\,
            I => \N__5993\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5993\,
            I => \N__5990\
        );

    \I__1018\ : Span4Mux_v
    port map (
            O => \N__5990\,
            I => \N__5987\
        );

    \I__1017\ : Span4Mux_v
    port map (
            O => \N__5987\,
            I => \N__5984\
        );

    \I__1016\ : Sp12to4
    port map (
            O => \N__5984\,
            I => \N__5981\
        );

    \I__1015\ : Span12Mux_h
    port map (
            O => \N__5981\,
            I => \N__5978\
        );

    \I__1014\ : Odrv12
    port map (
            O => \N__5978\,
            I => \A_c_15\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5975\,
            I => \N__5972\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5972\,
            I => \N__5969\
        );

    \I__1011\ : Span12Mux_v
    port map (
            O => \N__5969\,
            I => \N__5966\
        );

    \I__1010\ : Span12Mux_h
    port map (
            O => \N__5966\,
            I => \N__5963\
        );

    \I__1009\ : Odrv12
    port map (
            O => \N__5963\,
            I => \A_c_8\
        );

    \I__1008\ : InMux
    port map (
            O => \N__5960\,
            I => \N__5949\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5946\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5943\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5957\,
            I => \N__5940\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5956\,
            I => \N__5934\
        );

    \I__1003\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5931\
        );

    \I__1002\ : CascadeMux
    port map (
            O => \N__5954\,
            I => \N__5927\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5922\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5952\,
            I => \N__5922\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5949\,
            I => \N__5917\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__5946\,
            I => \N__5917\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5943\,
            I => \N__5914\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5940\,
            I => \N__5911\
        );

    \I__995\ : InMux
    port map (
            O => \N__5939\,
            I => \N__5904\
        );

    \I__994\ : InMux
    port map (
            O => \N__5938\,
            I => \N__5904\
        );

    \I__993\ : InMux
    port map (
            O => \N__5937\,
            I => \N__5904\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5934\,
            I => \N__5897\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5931\,
            I => \N__5897\
        );

    \I__990\ : InMux
    port map (
            O => \N__5930\,
            I => \N__5891\
        );

    \I__989\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5888\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5922\,
            I => \N__5885\
        );

    \I__987\ : Span4Mux_v
    port map (
            O => \N__5917\,
            I => \N__5876\
        );

    \I__986\ : Span4Mux_v
    port map (
            O => \N__5914\,
            I => \N__5876\
        );

    \I__985\ : Span4Mux_h
    port map (
            O => \N__5911\,
            I => \N__5876\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5904\,
            I => \N__5876\
        );

    \I__983\ : InMux
    port map (
            O => \N__5903\,
            I => \N__5873\
        );

    \I__982\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5870\
        );

    \I__981\ : Span4Mux_h
    port map (
            O => \N__5897\,
            I => \N__5867\
        );

    \I__980\ : InMux
    port map (
            O => \N__5896\,
            I => \N__5860\
        );

    \I__979\ : InMux
    port map (
            O => \N__5895\,
            I => \N__5860\
        );

    \I__978\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5860\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5891\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5888\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__975\ : Odrv4
    port map (
            O => \N__5885\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__974\ : Odrv4
    port map (
            O => \N__5876\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__5873\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5870\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__971\ : Odrv4
    port map (
            O => \N__5867\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5860\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__969\ : InMux
    port map (
            O => \N__5843\,
            I => \N__5835\
        );

    \I__968\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5830\
        );

    \I__967\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5830\
        );

    \I__966\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5827\
        );

    \I__965\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5824\
        );

    \I__964\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5819\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__5835\,
            I => \N__5814\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5830\,
            I => \N__5811\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__5827\,
            I => \N__5808\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__5824\,
            I => \N__5805\
        );

    \I__959\ : InMux
    port map (
            O => \N__5823\,
            I => \N__5800\
        );

    \I__958\ : InMux
    port map (
            O => \N__5822\,
            I => \N__5800\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__5819\,
            I => \N__5793\
        );

    \I__956\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5788\
        );

    \I__955\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5788\
        );

    \I__954\ : Span4Mux_v
    port map (
            O => \N__5814\,
            I => \N__5777\
        );

    \I__953\ : Span4Mux_v
    port map (
            O => \N__5811\,
            I => \N__5777\
        );

    \I__952\ : Span4Mux_v
    port map (
            O => \N__5808\,
            I => \N__5777\
        );

    \I__951\ : Span4Mux_h
    port map (
            O => \N__5805\,
            I => \N__5777\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5800\,
            I => \N__5777\
        );

    \I__949\ : InMux
    port map (
            O => \N__5799\,
            I => \N__5774\
        );

    \I__948\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5767\
        );

    \I__947\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5767\
        );

    \I__946\ : InMux
    port map (
            O => \N__5796\,
            I => \N__5767\
        );

    \I__945\ : Odrv4
    port map (
            O => \N__5793\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5788\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__943\ : Odrv4
    port map (
            O => \N__5777\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5774\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5767\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__5756\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_i_0_cascade_\
        );

    \I__939\ : CascadeMux
    port map (
            O => \N__5753\,
            I => \U712_BYTE_ENABLE.N_374_cascade_\
        );

    \I__938\ : IoInMux
    port map (
            O => \N__5750\,
            I => \N__5747\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__5747\,
            I => \N__5744\
        );

    \I__936\ : Span4Mux_s0_v
    port map (
            O => \N__5744\,
            I => \N__5741\
        );

    \I__935\ : Sp12to4
    port map (
            O => \N__5741\,
            I => \N__5738\
        );

    \I__934\ : Span12Mux_h
    port map (
            O => \N__5738\,
            I => \N__5735\
        );

    \I__933\ : Span12Mux_v
    port map (
            O => \N__5735\,
            I => \N__5732\
        );

    \I__932\ : Odrv12
    port map (
            O => \N__5732\,
            I => \N_51_i\
        );

    \I__931\ : IoInMux
    port map (
            O => \N__5729\,
            I => \N__5726\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__5726\,
            I => \N__5723\
        );

    \I__929\ : IoSpan4Mux
    port map (
            O => \N__5723\,
            I => \N__5719\
        );

    \I__928\ : InMux
    port map (
            O => \N__5722\,
            I => \N__5716\
        );

    \I__927\ : Span4Mux_s2_v
    port map (
            O => \N__5719\,
            I => \N__5713\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5716\,
            I => \N__5710\
        );

    \I__925\ : Span4Mux_v
    port map (
            O => \N__5713\,
            I => \N__5705\
        );

    \I__924\ : Span4Mux_v
    port map (
            O => \N__5710\,
            I => \N__5705\
        );

    \I__923\ : Odrv4
    port map (
            O => \N__5705\,
            I => \CONSTANT_ONE_NET\
        );

    \I__922\ : InMux
    port map (
            O => \N__5702\,
            I => \N__5699\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__5699\,
            I => \N__5696\
        );

    \I__920\ : Span12Mux_s11_v
    port map (
            O => \N__5696\,
            I => \N__5693\
        );

    \I__919\ : Span12Mux_h
    port map (
            O => \N__5693\,
            I => \N__5690\
        );

    \I__918\ : Odrv12
    port map (
            O => \N__5690\,
            I => \A_c_10\
        );

    \I__917\ : InMux
    port map (
            O => \N__5687\,
            I => \N__5684\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5684\,
            I => \N__5681\
        );

    \I__915\ : Span12Mux_v
    port map (
            O => \N__5681\,
            I => \N__5678\
        );

    \I__914\ : Span12Mux_h
    port map (
            O => \N__5678\,
            I => \N__5675\
        );

    \I__913\ : Span12Mux_v
    port map (
            O => \N__5675\,
            I => \N__5672\
        );

    \I__912\ : Odrv12
    port map (
            O => \N__5672\,
            I => \A_c_3\
        );

    \I__911\ : CascadeMux
    port map (
            O => \N__5669\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_1_cascade_\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__5666\,
            I => \U712_CHIP_RAM.N_322_cascade_\
        );

    \I__909\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5660\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__5660\,
            I => \N__5657\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__5657\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0\
        );

    \I__906\ : CEMux
    port map (
            O => \N__5654\,
            I => \N__5651\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__5651\,
            I => \N__5647\
        );

    \I__904\ : CEMux
    port map (
            O => \N__5650\,
            I => \N__5644\
        );

    \I__903\ : Span4Mux_v
    port map (
            O => \N__5647\,
            I => \N__5641\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5644\,
            I => \N__5638\
        );

    \I__901\ : Span4Mux_h
    port map (
            O => \N__5641\,
            I => \N__5635\
        );

    \I__900\ : Span4Mux_v
    port map (
            O => \N__5638\,
            I => \N__5632\
        );

    \I__899\ : Odrv4
    port map (
            O => \N__5635\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\
        );

    \I__898\ : Odrv4
    port map (
            O => \N__5632\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\
        );

    \I__897\ : InMux
    port map (
            O => \N__5627\,
            I => \N__5624\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5624\,
            I => \U712_REG_SM.N_289\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__5621\,
            I => \U712_REG_SM.N_358_cascade_\
        );

    \I__894\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5615\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5615\,
            I => \U712_REG_SM.N_360\
        );

    \I__892\ : InMux
    port map (
            O => \N__5612\,
            I => \N__5608\
        );

    \I__891\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5605\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5608\,
            I => \U712_REG_SM.N_359\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__5605\,
            I => \U712_REG_SM.N_359\
        );

    \I__888\ : InMux
    port map (
            O => \N__5600\,
            I => \N__5597\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5597\,
            I => \U712_REG_SM.N_270_i\
        );

    \I__886\ : InMux
    port map (
            O => \N__5594\,
            I => \N__5591\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5591\,
            I => \U712_REG_SM.REG_TACK_7\
        );

    \I__884\ : CascadeMux
    port map (
            O => \N__5588\,
            I => \N__5584\
        );

    \I__883\ : InMux
    port map (
            O => \N__5587\,
            I => \N__5581\
        );

    \I__882\ : InMux
    port map (
            O => \N__5584\,
            I => \N__5577\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5581\,
            I => \N__5574\
        );

    \I__880\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5571\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5577\,
            I => \REG_TACK\
        );

    \I__878\ : Odrv4
    port map (
            O => \N__5574\,
            I => \REG_TACK\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5571\,
            I => \REG_TACK\
        );

    \I__876\ : InMux
    port map (
            O => \N__5564\,
            I => \N__5561\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5561\,
            I => \N__5557\
        );

    \I__874\ : IoInMux
    port map (
            O => \N__5560\,
            I => \N__5554\
        );

    \I__873\ : Span4Mux_v
    port map (
            O => \N__5557\,
            I => \N__5551\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5554\,
            I => \N__5548\
        );

    \I__871\ : Sp12to4
    port map (
            O => \N__5551\,
            I => \N__5545\
        );

    \I__870\ : IoSpan4Mux
    port map (
            O => \N__5548\,
            I => \N__5542\
        );

    \I__869\ : Span12Mux_h
    port map (
            O => \N__5545\,
            I => \N__5539\
        );

    \I__868\ : IoSpan4Mux
    port map (
            O => \N__5542\,
            I => \N__5536\
        );

    \I__867\ : Span12Mux_v
    port map (
            O => \N__5539\,
            I => \N__5533\
        );

    \I__866\ : IoSpan4Mux
    port map (
            O => \N__5536\,
            I => \N__5530\
        );

    \I__865\ : Odrv12
    port map (
            O => \N__5533\,
            I => \C1_c\
        );

    \I__864\ : Odrv4
    port map (
            O => \N__5530\,
            I => \C1_c\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__5525\,
            I => \U712_REG_SM.N_340_cascade_\
        );

    \I__862\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5519\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5519\,
            I => \N__5516\
        );

    \I__860\ : Span4Mux_h
    port map (
            O => \N__5516\,
            I => \N__5513\
        );

    \I__859\ : Span4Mux_h
    port map (
            O => \N__5513\,
            I => \N__5510\
        );

    \I__858\ : Sp12to4
    port map (
            O => \N__5510\,
            I => \N__5507\
        );

    \I__857\ : Span12Mux_v
    port map (
            O => \N__5507\,
            I => \N__5504\
        );

    \I__856\ : Odrv12
    port map (
            O => \N__5504\,
            I => \REGSPACEn_c\
        );

    \I__855\ : IoInMux
    port map (
            O => \N__5501\,
            I => \N__5498\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__5498\,
            I => \N__5493\
        );

    \I__853\ : InMux
    port map (
            O => \N__5497\,
            I => \N__5490\
        );

    \I__852\ : InMux
    port map (
            O => \N__5496\,
            I => \N__5487\
        );

    \I__851\ : Span4Mux_s3_v
    port map (
            O => \N__5493\,
            I => \N__5484\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5490\,
            I => \N__5479\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5487\,
            I => \N__5479\
        );

    \I__848\ : Span4Mux_v
    port map (
            O => \N__5484\,
            I => \N__5476\
        );

    \I__847\ : Span4Mux_v
    port map (
            O => \N__5479\,
            I => \N__5473\
        );

    \I__846\ : Span4Mux_v
    port map (
            O => \N__5476\,
            I => \N__5469\
        );

    \I__845\ : Span4Mux_v
    port map (
            O => \N__5473\,
            I => \N__5466\
        );

    \I__844\ : InMux
    port map (
            O => \N__5472\,
            I => \N__5463\
        );

    \I__843\ : Odrv4
    port map (
            O => \N__5469\,
            I => \DBENn_c\
        );

    \I__842\ : Odrv4
    port map (
            O => \N__5466\,
            I => \DBENn_c\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5463\,
            I => \DBENn_c\
        );

    \I__840\ : InMux
    port map (
            O => \N__5456\,
            I => \N__5452\
        );

    \I__839\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5449\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5452\,
            I => \N__5443\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5449\,
            I => \N__5443\
        );

    \I__836\ : InMux
    port map (
            O => \N__5448\,
            I => \N__5439\
        );

    \I__835\ : Span4Mux_v
    port map (
            O => \N__5443\,
            I => \N__5436\
        );

    \I__834\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5432\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__5439\,
            I => \N__5428\
        );

    \I__832\ : Span4Mux_v
    port map (
            O => \N__5436\,
            I => \N__5425\
        );

    \I__831\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5422\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5432\,
            I => \N__5419\
        );

    \I__829\ : InMux
    port map (
            O => \N__5431\,
            I => \N__5416\
        );

    \I__828\ : Span4Mux_h
    port map (
            O => \N__5428\,
            I => \N__5413\
        );

    \I__827\ : Odrv4
    port map (
            O => \N__5425\,
            I => \DMA_CYCLEm\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5422\,
            I => \DMA_CYCLEm\
        );

    \I__825\ : Odrv12
    port map (
            O => \N__5419\,
            I => \DMA_CYCLEm\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5416\,
            I => \DMA_CYCLEm\
        );

    \I__823\ : Odrv4
    port map (
            O => \N__5413\,
            I => \DMA_CYCLEm\
        );

    \I__822\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5398\
        );

    \I__821\ : InMux
    port map (
            O => \N__5401\,
            I => \N__5395\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5398\,
            I => \N__5390\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__5395\,
            I => \N__5390\
        );

    \I__818\ : Span4Mux_v
    port map (
            O => \N__5390\,
            I => \N__5387\
        );

    \I__817\ : Sp12to4
    port map (
            O => \N__5387\,
            I => \N__5384\
        );

    \I__816\ : Span12Mux_h
    port map (
            O => \N__5384\,
            I => \N__5381\
        );

    \I__815\ : Span12Mux_v
    port map (
            O => \N__5381\,
            I => \N__5378\
        );

    \I__814\ : Odrv12
    port map (
            O => \N__5378\,
            I => \TSn_c\
        );

    \I__813\ : InMux
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5372\,
            I => \N__5369\
        );

    \I__811\ : Span4Mux_h
    port map (
            O => \N__5369\,
            I => \N__5366\
        );

    \I__810\ : Span4Mux_v
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__809\ : Span4Mux_v
    port map (
            O => \N__5363\,
            I => \N__5360\
        );

    \I__808\ : Span4Mux_v
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__807\ : Odrv4
    port map (
            O => \N__5357\,
            I => \RAMSPACEn_c\
        );

    \I__806\ : InMux
    port map (
            O => \N__5354\,
            I => \N__5351\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5351\,
            I => \N__5348\
        );

    \I__804\ : Odrv12
    port map (
            O => \N__5348\,
            I => \U712_CHIP_RAM.N_345\
        );

    \I__803\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5341\
        );

    \I__802\ : InMux
    port map (
            O => \N__5344\,
            I => \N__5338\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5341\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__5338\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__5333\,
            I => \N__5329\
        );

    \I__798\ : InMux
    port map (
            O => \N__5332\,
            I => \N__5326\
        );

    \I__797\ : InMux
    port map (
            O => \N__5329\,
            I => \N__5322\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5326\,
            I => \N__5319\
        );

    \I__795\ : InMux
    port map (
            O => \N__5325\,
            I => \N__5316\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__5322\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__793\ : Odrv4
    port map (
            O => \N__5319\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5316\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__5309\,
            I => \U712_REG_SM.m17_i_0_o2_1_cascade_\
        );

    \I__790\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5303\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5303\,
            I => \N__5300\
        );

    \I__788\ : Span4Mux_h
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__787\ : Span4Mux_v
    port map (
            O => \N__5297\,
            I => \N__5294\
        );

    \I__786\ : Sp12to4
    port map (
            O => \N__5294\,
            I => \N__5291\
        );

    \I__785\ : Odrv12
    port map (
            O => \N__5291\,
            I => \A_c_7\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__5288\,
            I => \U712_REG_SM.C3_SYNC_RNI7UAPZ0Z_1_cascade_\
        );

    \I__783\ : InMux
    port map (
            O => \N__5285\,
            I => \N__5279\
        );

    \I__782\ : InMux
    port map (
            O => \N__5284\,
            I => \N__5274\
        );

    \I__781\ : InMux
    port map (
            O => \N__5283\,
            I => \N__5274\
        );

    \I__780\ : InMux
    port map (
            O => \N__5282\,
            I => \N__5271\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5279\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5274\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5271\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__776\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5257\
        );

    \I__775\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5252\
        );

    \I__774\ : InMux
    port map (
            O => \N__5262\,
            I => \N__5252\
        );

    \I__773\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5247\
        );

    \I__772\ : InMux
    port map (
            O => \N__5260\,
            I => \N__5247\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5257\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5252\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5247\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__5240\,
            I => \U712_REG_SM.m15_i_0_a2_0_0_cascade_\
        );

    \I__767\ : InMux
    port map (
            O => \N__5237\,
            I => \N__5234\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5234\,
            I => \U712_CHIP_RAM.N_386\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__5231\,
            I => \U712_CHIP_RAM.N_434_cascade_\
        );

    \I__764\ : InMux
    port map (
            O => \N__5228\,
            I => \N__5225\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__5225\,
            I => \N__5222\
        );

    \I__762\ : Span4Mux_h
    port map (
            O => \N__5222\,
            I => \N__5217\
        );

    \I__761\ : InMux
    port map (
            O => \N__5221\,
            I => \N__5212\
        );

    \I__760\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5212\
        );

    \I__759\ : Odrv4
    port map (
            O => \N__5217\,
            I => \U712_CHIP_RAM.N_439\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5212\,
            I => \U712_CHIP_RAM.N_439\
        );

    \I__757\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5204\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__5204\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_a2_0\
        );

    \I__755\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5198\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5198\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__753\ : InMux
    port map (
            O => \N__5195\,
            I => \N__5192\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__5192\,
            I => \N__5189\
        );

    \I__751\ : Span4Mux_v
    port map (
            O => \N__5189\,
            I => \N__5186\
        );

    \I__750\ : Span4Mux_h
    port map (
            O => \N__5186\,
            I => \N__5183\
        );

    \I__749\ : Sp12to4
    port map (
            O => \N__5183\,
            I => \N__5180\
        );

    \I__748\ : Odrv12
    port map (
            O => \N__5180\,
            I => \A_c_12\
        );

    \I__747\ : InMux
    port map (
            O => \N__5177\,
            I => \N__5174\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__5174\,
            I => \N__5171\
        );

    \I__745\ : Span4Mux_h
    port map (
            O => \N__5171\,
            I => \N__5168\
        );

    \I__744\ : Sp12to4
    port map (
            O => \N__5168\,
            I => \N__5165\
        );

    \I__743\ : Span12Mux_v
    port map (
            O => \N__5165\,
            I => \N__5162\
        );

    \I__742\ : Odrv12
    port map (
            O => \N__5162\,
            I => \A_c_5\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__5159\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_cascade_\
        );

    \I__740\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5153\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5153\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_1\
        );

    \I__738\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5146\
        );

    \I__737\ : InMux
    port map (
            O => \N__5149\,
            I => \N__5142\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__5146\,
            I => \N__5139\
        );

    \I__735\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5136\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__5142\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__733\ : Odrv4
    port map (
            O => \N__5139\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__5136\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__731\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5124\
        );

    \I__730\ : InMux
    port map (
            O => \N__5128\,
            I => \N__5121\
        );

    \I__729\ : InMux
    port map (
            O => \N__5127\,
            I => \N__5118\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__5124\,
            I => \N__5115\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__5121\,
            I => \CPU_TACKm\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5118\,
            I => \CPU_TACKm\
        );

    \I__725\ : Odrv12
    port map (
            O => \N__5115\,
            I => \CPU_TACKm\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__5108\,
            I => \N__5103\
        );

    \I__723\ : InMux
    port map (
            O => \N__5107\,
            I => \N__5099\
        );

    \I__722\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5096\
        );

    \I__721\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5093\
        );

    \I__720\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5090\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__5099\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5096\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5093\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5090\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__5081\,
            I => \U712_CYCLE_TERM.N_351_cascade_\
        );

    \I__714\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5073\
        );

    \I__713\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5069\
        );

    \I__712\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5066\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__5073\,
            I => \N__5063\
        );

    \I__710\ : InMux
    port map (
            O => \N__5072\,
            I => \N__5060\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__5069\,
            I => \N__5055\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__5066\,
            I => \N__5055\
        );

    \I__707\ : Span4Mux_v
    port map (
            O => \N__5063\,
            I => \N__5050\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5060\,
            I => \N__5050\
        );

    \I__705\ : Span4Mux_v
    port map (
            O => \N__5055\,
            I => \N__5047\
        );

    \I__704\ : Span4Mux_h
    port map (
            O => \N__5050\,
            I => \N__5044\
        );

    \I__703\ : Sp12to4
    port map (
            O => \N__5047\,
            I => \N__5041\
        );

    \I__702\ : Span4Mux_h
    port map (
            O => \N__5044\,
            I => \N__5038\
        );

    \I__701\ : Span12Mux_h
    port map (
            O => \N__5041\,
            I => \N__5033\
        );

    \I__700\ : Sp12to4
    port map (
            O => \N__5038\,
            I => \N__5033\
        );

    \I__699\ : Span12Mux_v
    port map (
            O => \N__5033\,
            I => \N__5030\
        );

    \I__698\ : Odrv12
    port map (
            O => \N__5030\,
            I => \CLK40_PLL_i\
        );

    \I__697\ : InMux
    port map (
            O => \N__5027\,
            I => \N__5024\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5024\,
            I => \N__5020\
        );

    \I__695\ : InMux
    port map (
            O => \N__5023\,
            I => \N__5017\
        );

    \I__694\ : Span4Mux_v
    port map (
            O => \N__5020\,
            I => \N__5012\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__5017\,
            I => \N__5009\
        );

    \I__692\ : InMux
    port map (
            O => \N__5016\,
            I => \N__5006\
        );

    \I__691\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5003\
        );

    \I__690\ : Odrv4
    port map (
            O => \N__5012\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__689\ : Odrv4
    port map (
            O => \N__5009\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__5006\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__5003\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__686\ : InMux
    port map (
            O => \N__4994\,
            I => \N__4990\
        );

    \I__685\ : InMux
    port map (
            O => \N__4993\,
            I => \N__4987\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__4990\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4987\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0\
        );

    \I__682\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4979\,
            I => \N__4976\
        );

    \I__680\ : Odrv4
    port map (
            O => \N__4976\,
            I => \U712_CHIP_RAM.N_325\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__4973\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\
        );

    \I__678\ : InMux
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4967\,
            I => \N__4964\
        );

    \I__676\ : Odrv4
    port map (
            O => \N__4964\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__675\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4957\
        );

    \I__674\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4954\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4957\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4954\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__671\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4945\
        );

    \I__670\ : InMux
    port map (
            O => \N__4948\,
            I => \N__4942\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__4945\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4942\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__4937\,
            I => \N__4933\
        );

    \I__666\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4930\
        );

    \I__665\ : InMux
    port map (
            O => \N__4933\,
            I => \N__4927\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4930\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4927\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__662\ : InMux
    port map (
            O => \N__4922\,
            I => \N__4918\
        );

    \I__661\ : InMux
    port map (
            O => \N__4921\,
            I => \N__4915\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4918\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__4915\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__4910\,
            I => \U712_CHIP_RAM.N_241_cascade_\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__4907\,
            I => \U712_CHIP_RAM.N_388_cascade_\
        );

    \I__656\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4900\
        );

    \I__655\ : InMux
    port map (
            O => \N__4903\,
            I => \N__4897\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4900\,
            I => \U712_CHIP_RAM.N_325_1\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4897\,
            I => \U712_CHIP_RAM.N_325_1\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__4892\,
            I => \N__4888\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__4891\,
            I => \N__4884\
        );

    \I__650\ : InMux
    port map (
            O => \N__4888\,
            I => \N__4879\
        );

    \I__649\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4875\
        );

    \I__648\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4872\
        );

    \I__647\ : InMux
    port map (
            O => \N__4883\,
            I => \N__4867\
        );

    \I__646\ : InMux
    port map (
            O => \N__4882\,
            I => \N__4867\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4879\,
            I => \N__4864\
        );

    \I__644\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4861\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4875\,
            I => \U712_CHIP_RAM.N_381\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__4872\,
            I => \U712_CHIP_RAM.N_381\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__4867\,
            I => \U712_CHIP_RAM.N_381\
        );

    \I__640\ : Odrv4
    port map (
            O => \N__4864\,
            I => \U712_CHIP_RAM.N_381\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4861\,
            I => \U712_CHIP_RAM.N_381\
        );

    \I__638\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4844\
        );

    \I__637\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4844\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__4844\,
            I => \N__4841\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__4841\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__634\ : IoInMux
    port map (
            O => \N__4838\,
            I => \N__4835\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4835\,
            I => \N__4832\
        );

    \I__632\ : IoSpan4Mux
    port map (
            O => \N__4832\,
            I => \N__4829\
        );

    \I__631\ : Span4Mux_s3_v
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__630\ : Span4Mux_v
    port map (
            O => \N__4826\,
            I => \N__4823\
        );

    \I__629\ : Odrv4
    port map (
            O => \N__4823\,
            I => \N_249_i\
        );

    \I__628\ : InMux
    port map (
            O => \N__4820\,
            I => \N__4817\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__4817\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1_0\
        );

    \I__626\ : CascadeMux
    port map (
            O => \N__4814\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1_tz_cascade_\
        );

    \I__625\ : CascadeMux
    port map (
            O => \N__4811\,
            I => \U712_CHIP_RAM.N_325_cascade_\
        );

    \I__624\ : IoInMux
    port map (
            O => \N__4808\,
            I => \N__4805\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__4805\,
            I => \N__4802\
        );

    \I__622\ : IoSpan4Mux
    port map (
            O => \N__4802\,
            I => \N__4799\
        );

    \I__621\ : Span4Mux_s3_h
    port map (
            O => \N__4799\,
            I => \N__4795\
        );

    \I__620\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4792\
        );

    \I__619\ : Span4Mux_h
    port map (
            O => \N__4795\,
            I => \N__4789\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__4792\,
            I => \N__4786\
        );

    \I__617\ : Sp12to4
    port map (
            O => \N__4789\,
            I => \N__4783\
        );

    \I__616\ : Span4Mux_v
    port map (
            O => \N__4786\,
            I => \N__4780\
        );

    \I__615\ : Span12Mux_h
    port map (
            O => \N__4783\,
            I => \N__4775\
        );

    \I__614\ : Sp12to4
    port map (
            O => \N__4780\,
            I => \N__4775\
        );

    \I__613\ : Span12Mux_h
    port map (
            O => \N__4775\,
            I => \N__4772\
        );

    \I__612\ : Span12Mux_v
    port map (
            O => \N__4772\,
            I => \N__4769\
        );

    \I__611\ : Odrv12
    port map (
            O => \N__4769\,
            I => \C3_c\
        );

    \I__610\ : InMux
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__4763\,
            I => \N__4759\
        );

    \I__608\ : InMux
    port map (
            O => \N__4762\,
            I => \N__4756\
        );

    \I__607\ : Span4Mux_h
    port map (
            O => \N__4759\,
            I => \N__4751\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__4756\,
            I => \N__4751\
        );

    \I__605\ : Span4Mux_v
    port map (
            O => \N__4751\,
            I => \N__4748\
        );

    \I__604\ : Span4Mux_h
    port map (
            O => \N__4748\,
            I => \N__4745\
        );

    \I__603\ : Sp12to4
    port map (
            O => \N__4745\,
            I => \N__4742\
        );

    \I__602\ : Span12Mux_v
    port map (
            O => \N__4742\,
            I => \N__4739\
        );

    \I__601\ : Odrv12
    port map (
            O => \N__4739\,
            I => \DBRn_c\
        );

    \I__600\ : InMux
    port map (
            O => \N__4736\,
            I => \N__4733\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4733\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__598\ : InMux
    port map (
            O => \N__4730\,
            I => \N__4727\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4727\,
            I => \N__4724\
        );

    \I__596\ : Span4Mux_h
    port map (
            O => \N__4724\,
            I => \N__4721\
        );

    \I__595\ : Sp12to4
    port map (
            O => \N__4721\,
            I => \N__4718\
        );

    \I__594\ : Span12Mux_v
    port map (
            O => \N__4718\,
            I => \N__4715\
        );

    \I__593\ : Odrv12
    port map (
            O => \N__4715\,
            I => \A_c_20\
        );

    \I__592\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4709\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4709\,
            I => \N__4706\
        );

    \I__590\ : Span4Mux_v
    port map (
            O => \N__4706\,
            I => \N__4703\
        );

    \I__589\ : Odrv4
    port map (
            O => \N__4703\,
            I => \U712_CHIP_RAM.BANK0_9_u_0_0_a2_0_0\
        );

    \I__588\ : InMux
    port map (
            O => \N__4700\,
            I => \N__4696\
        );

    \I__587\ : InMux
    port map (
            O => \N__4699\,
            I => \N__4693\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4696\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__4693\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__584\ : CascadeMux
    port map (
            O => \N__4688\,
            I => \N__4685\
        );

    \I__583\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4681\
        );

    \I__582\ : InMux
    port map (
            O => \N__4684\,
            I => \N__4678\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__4681\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4678\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__4673\,
            I => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\
        );

    \I__578\ : CascadeMux
    port map (
            O => \N__4670\,
            I => \U712_CYCLE_TERM.N_269_i_0_en_cascade_\
        );

    \I__577\ : CEMux
    port map (
            O => \N__4667\,
            I => \N__4664\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__4664\,
            I => \N__4661\
        );

    \I__575\ : Odrv4
    port map (
            O => \N__4661\,
            I => \U712_CYCLE_TERM.N_269_i_0_en_0\
        );

    \I__574\ : CascadeMux
    port map (
            O => \N__4658\,
            I => \U712_CHIP_RAM.N_76_cascade_\
        );

    \I__573\ : InMux
    port map (
            O => \N__4655\,
            I => \N__4651\
        );

    \I__572\ : InMux
    port map (
            O => \N__4654\,
            I => \N__4648\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4651\,
            I => \U712_CHIP_RAM.N_328\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4648\,
            I => \U712_CHIP_RAM.N_328\
        );

    \I__569\ : IoInMux
    port map (
            O => \N__4643\,
            I => \N__4640\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4640\,
            I => \N__4637\
        );

    \I__567\ : Span4Mux_s3_v
    port map (
            O => \N__4637\,
            I => \N__4634\
        );

    \I__566\ : Sp12to4
    port map (
            O => \N__4634\,
            I => \N__4631\
        );

    \I__565\ : Span12Mux_s11_h
    port map (
            O => \N__4631\,
            I => \N__4628\
        );

    \I__564\ : Span12Mux_v
    port map (
            O => \N__4628\,
            I => \N__4624\
        );

    \I__563\ : InMux
    port map (
            O => \N__4627\,
            I => \N__4621\
        );

    \I__562\ : Odrv12
    port map (
            O => \N__4624\,
            I => \LATCH_CLK_c\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__4621\,
            I => \LATCH_CLK_c\
        );

    \I__560\ : CascadeMux
    port map (
            O => \N__4616\,
            I => \U712_CHIP_RAM.N_438_cascade_\
        );

    \I__559\ : InMux
    port map (
            O => \N__4613\,
            I => \N__4607\
        );

    \I__558\ : InMux
    port map (
            O => \N__4612\,
            I => \N__4607\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__4607\,
            I => \U712_CHIP_RAM.N_336\
        );

    \I__556\ : CascadeMux
    port map (
            O => \N__4604\,
            I => \N__4600\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__4603\,
            I => \N__4595\
        );

    \I__554\ : InMux
    port map (
            O => \N__4600\,
            I => \N__4592\
        );

    \I__553\ : InMux
    port map (
            O => \N__4599\,
            I => \N__4589\
        );

    \I__552\ : InMux
    port map (
            O => \N__4598\,
            I => \N__4585\
        );

    \I__551\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4582\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4592\,
            I => \N__4577\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4589\,
            I => \N__4577\
        );

    \I__548\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4574\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4585\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__4582\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__4577\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4574\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__543\ : InMux
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4562\,
            I => \N__4559\
        );

    \I__541\ : Span4Mux_h
    port map (
            O => \N__4559\,
            I => \N__4556\
        );

    \I__540\ : Odrv4
    port map (
            O => \N__4556\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__4553\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\
        );

    \I__538\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4546\
        );

    \I__537\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4543\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4546\,
            I => \U712_CHIP_RAM.N_438\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4543\,
            I => \U712_CHIP_RAM.N_438\
        );

    \I__534\ : InMux
    port map (
            O => \N__4538\,
            I => \N__4535\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__4535\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0_a2_0\
        );

    \I__532\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4529\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__4529\,
            I => \U712_CHIP_RAM.N_247\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__4526\,
            I => \U712_CHIP_RAM.N_247_cascade_\
        );

    \I__529\ : InMux
    port map (
            O => \N__4523\,
            I => \N__4520\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__4520\,
            I => \N__4517\
        );

    \I__527\ : Span4Mux_h
    port map (
            O => \N__4517\,
            I => \N__4513\
        );

    \I__526\ : InMux
    port map (
            O => \N__4516\,
            I => \N__4510\
        );

    \I__525\ : Odrv4
    port map (
            O => \N__4513\,
            I => \U712_CHIP_RAM.N_244\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4510\,
            I => \U712_CHIP_RAM.N_244\
        );

    \I__523\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4502\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4502\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_0\
        );

    \I__521\ : InMux
    port map (
            O => \N__4499\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__520\ : InMux
    port map (
            O => \N__4496\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__519\ : InMux
    port map (
            O => \N__4493\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__518\ : InMux
    port map (
            O => \N__4490\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__517\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4474\
        );

    \I__516\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4474\
        );

    \I__515\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4474\
        );

    \I__514\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4471\
        );

    \I__513\ : InMux
    port map (
            O => \N__4483\,
            I => \N__4464\
        );

    \I__512\ : InMux
    port map (
            O => \N__4482\,
            I => \N__4464\
        );

    \I__511\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4464\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__4474\,
            I => \U712_CHIP_RAM.N_236\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4471\,
            I => \U712_CHIP_RAM.N_236\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4464\,
            I => \U712_CHIP_RAM.N_236\
        );

    \I__507\ : InMux
    port map (
            O => \N__4457\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__506\ : CEMux
    port map (
            O => \N__4454\,
            I => \N__4451\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4451\,
            I => \N__4447\
        );

    \I__504\ : CEMux
    port map (
            O => \N__4450\,
            I => \N__4444\
        );

    \I__503\ : Span4Mux_v
    port map (
            O => \N__4447\,
            I => \N__4441\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4444\,
            I => \N__4438\
        );

    \I__501\ : Span4Mux_h
    port map (
            O => \N__4441\,
            I => \N__4435\
        );

    \I__500\ : Span4Mux_h
    port map (
            O => \N__4438\,
            I => \N__4432\
        );

    \I__499\ : Odrv4
    port map (
            O => \N__4435\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__498\ : Odrv4
    port map (
            O => \N__4432\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__4427\,
            I => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0_cascade_\
        );

    \I__496\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4421\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_1\
        );

    \I__494\ : InMux
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__4415\,
            I => \U712_CHIP_RAM.N_348\
        );

    \I__492\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4409\,
            I => \N__4405\
        );

    \I__490\ : InMux
    port map (
            O => \N__4408\,
            I => \N__4402\
        );

    \I__489\ : Odrv4
    port map (
            O => \N__4405\,
            I => \U712_CHIP_RAM.N_437\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4402\,
            I => \U712_CHIP_RAM.N_437\
        );

    \I__487\ : CascadeMux
    port map (
            O => \N__4397\,
            I => \N__4393\
        );

    \I__486\ : InMux
    port map (
            O => \N__4396\,
            I => \N__4388\
        );

    \I__485\ : InMux
    port map (
            O => \N__4393\,
            I => \N__4385\
        );

    \I__484\ : InMux
    port map (
            O => \N__4392\,
            I => \N__4382\
        );

    \I__483\ : InMux
    port map (
            O => \N__4391\,
            I => \N__4379\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4388\,
            I => \U712_CHIP_RAM.N_426\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4385\,
            I => \U712_CHIP_RAM.N_426\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__4382\,
            I => \U712_CHIP_RAM.N_426\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4379\,
            I => \U712_CHIP_RAM.N_426\
        );

    \I__478\ : CascadeMux
    port map (
            O => \N__4370\,
            I => \U712_CHIP_RAM.N_300_cascade_\
        );

    \I__477\ : InMux
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4364\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__475\ : InMux
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4358\,
            I => \U712_CHIP_RAM.DMA_CYCLE_esr_RNIULZ0Z431\
        );

    \I__473\ : InMux
    port map (
            O => \N__4355\,
            I => \N__4352\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4352\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_1\
        );

    \I__471\ : InMux
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4346\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_1\
        );

    \I__469\ : InMux
    port map (
            O => \N__4343\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__468\ : InMux
    port map (
            O => \N__4340\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__4337\,
            I => \N__4334\
        );

    \I__466\ : InMux
    port map (
            O => \N__4334\,
            I => \N__4329\
        );

    \I__465\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4324\
        );

    \I__464\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4324\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4329\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4324\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__461\ : CascadeMux
    port map (
            O => \N__4319\,
            I => \N__4316\
        );

    \I__460\ : InMux
    port map (
            O => \N__4316\,
            I => \N__4310\
        );

    \I__459\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4310\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4310\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__457\ : InMux
    port map (
            O => \N__4307\,
            I => \N__4304\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__4304\,
            I => \N__4301\
        );

    \I__455\ : Span4Mux_v
    port map (
            O => \N__4301\,
            I => \N__4298\
        );

    \I__454\ : Odrv4
    port map (
            O => \N__4298\,
            I => \TACK_EN_i_ess\
        );

    \I__453\ : IoInMux
    port map (
            O => \N__4295\,
            I => \N__4292\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__451\ : Odrv12
    port map (
            O => \N__4289\,
            I => \VBENn_c\
        );

    \I__450\ : CascadeMux
    port map (
            O => \N__4286\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_0_cascade_\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__4283\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_cascade_\
        );

    \I__448\ : CEMux
    port map (
            O => \N__4280\,
            I => \N__4277\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__4277\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0\
        );

    \I__446\ : InMux
    port map (
            O => \N__4274\,
            I => \N__4271\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4271\,
            I => \N__4268\
        );

    \I__444\ : Odrv4
    port map (
            O => \N__4268\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_a2_0\
        );

    \I__443\ : CascadeMux
    port map (
            O => \N__4265\,
            I => \U712_CHIP_RAM.N_350_cascade_\
        );

    \I__442\ : CascadeMux
    port map (
            O => \N__4262\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_\
        );

    \I__441\ : CEMux
    port map (
            O => \N__4259\,
            I => \N__4256\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4256\,
            I => \N__4253\
        );

    \I__439\ : Span4Mux_h
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__438\ : Odrv4
    port map (
            O => \N__4250\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0\
        );

    \I__437\ : InMux
    port map (
            O => \N__4247\,
            I => \N__4244\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4244\,
            I => \U712_CHIP_RAM.N_350\
        );

    \I__435\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4237\
        );

    \I__434\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4234\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__4237\,
            I => \N__4231\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__4234\,
            I => \N__4228\
        );

    \I__431\ : Span4Mux_h
    port map (
            O => \N__4231\,
            I => \N__4223\
        );

    \I__430\ : Span4Mux_v
    port map (
            O => \N__4228\,
            I => \N__4223\
        );

    \I__429\ : Sp12to4
    port map (
            O => \N__4223\,
            I => \N__4220\
        );

    \I__428\ : Span12Mux_h
    port map (
            O => \N__4220\,
            I => \N__4217\
        );

    \I__427\ : Span12Mux_v
    port map (
            O => \N__4217\,
            I => \N__4214\
        );

    \I__426\ : Odrv12
    port map (
            O => \N__4214\,
            I => \AWEn_c\
        );

    \I__425\ : InMux
    port map (
            O => \N__4211\,
            I => \N__4208\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__4208\,
            I => \U712_CHIP_RAM.N_287\
        );

    \I__423\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4202\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4202\,
            I => \U712_CHIP_RAM.un3_DMA_CYCLE_START\
        );

    \I__421\ : InMux
    port map (
            O => \N__4199\,
            I => \N__4196\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__4196\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__4193\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_a2_0_cascade_\
        );

    \I__418\ : CascadeMux
    port map (
            O => \N__4190\,
            I => \U712_CHIP_RAM.N_265_cascade_\
        );

    \I__417\ : InMux
    port map (
            O => \N__4187\,
            I => \N__4184\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__4184\,
            I => \U712_CHIP_RAM.N_265\
        );

    \I__415\ : CascadeMux
    port map (
            O => \N__4181\,
            I => \U712_CHIP_RAM.N_236_cascade_\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__4178\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__4175\,
            I => \U712_CHIP_RAM.N_426_cascade_\
        );

    \I__412\ : IoInMux
    port map (
            O => \N__4172\,
            I => \N__4169\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__4169\,
            I => \N__4166\
        );

    \I__410\ : IoSpan4Mux
    port map (
            O => \N__4166\,
            I => \N__4163\
        );

    \I__409\ : Span4Mux_s3_v
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__408\ : Span4Mux_v
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__407\ : Span4Mux_v
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__406\ : Odrv4
    port map (
            O => \N__4154\,
            I => \BANK0_c\
        );

    \I__405\ : InMux
    port map (
            O => \N__4151\,
            I => \N__4148\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4148\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\
        );

    \I__403\ : CascadeMux
    port map (
            O => \N__4145\,
            I => \U712_CHIP_RAM.N_186_cascade_\
        );

    \I__402\ : IoInMux
    port map (
            O => \N__4142\,
            I => \N__4139\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__4139\,
            I => \N__4136\
        );

    \I__400\ : Span4Mux_s3_v
    port map (
            O => \N__4136\,
            I => \N__4133\
        );

    \I__399\ : Span4Mux_v
    port map (
            O => \N__4133\,
            I => \N__4129\
        );

    \I__398\ : InMux
    port map (
            O => \N__4132\,
            I => \N__4126\
        );

    \I__397\ : Odrv4
    port map (
            O => \N__4129\,
            I => \DBDIR_c\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__4126\,
            I => \DBDIR_c\
        );

    \I__395\ : IoInMux
    port map (
            O => \N__4121\,
            I => \N__4118\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__4118\,
            I => \N__4115\
        );

    \I__393\ : Span4Mux_s2_h
    port map (
            O => \N__4115\,
            I => \N__4112\
        );

    \I__392\ : Sp12to4
    port map (
            O => \N__4112\,
            I => \N__4109\
        );

    \I__391\ : Span12Mux_v
    port map (
            O => \N__4109\,
            I => \N__4105\
        );

    \I__390\ : InMux
    port map (
            O => \N__4108\,
            I => \N__4102\
        );

    \I__389\ : Odrv12
    port map (
            O => \N__4105\,
            I => \TACK_OUTn\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__4102\,
            I => \TACK_OUTn\
        );

    \I__387\ : IoInMux
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__4094\,
            I => \N__4090\
        );

    \I__385\ : IoInMux
    port map (
            O => \N__4093\,
            I => \N__4087\
        );

    \I__384\ : IoSpan4Mux
    port map (
            O => \N__4090\,
            I => \N__4082\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__4087\,
            I => \N__4082\
        );

    \I__382\ : IoSpan4Mux
    port map (
            O => \N__4082\,
            I => \N__4078\
        );

    \I__381\ : IoInMux
    port map (
            O => \N__4081\,
            I => \N__4075\
        );

    \I__380\ : IoSpan4Mux
    port map (
            O => \N__4078\,
            I => \N__4072\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__4075\,
            I => \N__4069\
        );

    \I__378\ : Sp12to4
    port map (
            O => \N__4072\,
            I => \N__4066\
        );

    \I__377\ : IoSpan4Mux
    port map (
            O => \N__4069\,
            I => \N__4063\
        );

    \I__376\ : Span12Mux_s6_v
    port map (
            O => \N__4066\,
            I => \N__4060\
        );

    \I__375\ : Span4Mux_s2_h
    port map (
            O => \N__4063\,
            I => \N__4057\
        );

    \I__374\ : Span12Mux_h
    port map (
            O => \N__4060\,
            I => \N__4054\
        );

    \I__373\ : Span4Mux_h
    port map (
            O => \N__4057\,
            I => \N__4051\
        );

    \I__372\ : Odrv12
    port map (
            O => \N__4054\,
            I => \CLK40_PLL_i_i\
        );

    \I__371\ : Odrv4
    port map (
            O => \N__4051\,
            I => \CLK40_PLL_i_i\
        );

    \I__370\ : CascadeMux
    port map (
            O => \N__4046\,
            I => \N__4043\
        );

    \I__369\ : InMux
    port map (
            O => \N__4043\,
            I => \N__4040\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__4040\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_i_i_a2_0\
        );

    \I__367\ : IoInMux
    port map (
            O => \N__4037\,
            I => \N__4034\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__4034\,
            I => \N__4031\
        );

    \I__365\ : IoSpan4Mux
    port map (
            O => \N__4031\,
            I => \N__4028\
        );

    \I__364\ : Span4Mux_s3_h
    port map (
            O => \N__4028\,
            I => \N__4025\
        );

    \I__363\ : Odrv4
    port map (
            O => \N__4025\,
            I => \DBRn_c_i_0\
        );

    \I__362\ : IoInMux
    port map (
            O => \N__4022\,
            I => \N__4019\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__4019\,
            I => \N__4016\
        );

    \I__360\ : Span4Mux_s2_h
    port map (
            O => \N__4016\,
            I => \N__4013\
        );

    \I__359\ : Span4Mux_h
    port map (
            O => \N__4013\,
            I => \N__4010\
        );

    \I__358\ : Span4Mux_v
    port map (
            O => \N__4010\,
            I => \N__4007\
        );

    \I__357\ : Odrv4
    port map (
            O => \N__4007\,
            I => \N_996_i\
        );

    \I__356\ : IoInMux
    port map (
            O => \N__4004\,
            I => \N__4001\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__4001\,
            I => \N__3998\
        );

    \I__354\ : Span4Mux_s2_v
    port map (
            O => \N__3998\,
            I => \N__3995\
        );

    \I__353\ : Span4Mux_v
    port map (
            O => \N__3995\,
            I => \N__3992\
        );

    \I__352\ : Span4Mux_h
    port map (
            O => \N__3992\,
            I => \N__3989\
        );

    \I__351\ : Odrv4
    port map (
            O => \N__3989\,
            I => \CLK80_PLL_i_i\
        );

    \I__350\ : IoInMux
    port map (
            O => \N__3986\,
            I => \N__3983\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__3983\,
            I => \N__3980\
        );

    \I__348\ : Span4Mux_s0_v
    port map (
            O => \N__3980\,
            I => \N__3977\
        );

    \I__347\ : Span4Mux_v
    port map (
            O => \N__3977\,
            I => \N__3974\
        );

    \I__346\ : Sp12to4
    port map (
            O => \N__3974\,
            I => \N__3971\
        );

    \I__345\ : Span12Mux_h
    port map (
            O => \N__3971\,
            I => \N__3968\
        );

    \I__344\ : Span12Mux_v
    port map (
            O => \N__3968\,
            I => \N__3965\
        );

    \I__343\ : Odrv12
    port map (
            O => \N__3965\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__7693\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__7695\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__7690\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__7692\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__7687\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__7688\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__7689\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__7691\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7349\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5560\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4037\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4808\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10997\,
            in2 => \_gnd_net_\,
            in3 => \N__7999\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4307\,
            lcout => \N_996_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4762\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8696\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011101110"
        )
    port map (
            in0 => \N__5472\,
            in1 => \N__4151\,
            in2 => \N__4603\,
            in3 => \N__10316\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8679\,
            ce => 'H',
            sr => \N__10976\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNICLGI4_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__4391\,
            in1 => \N__6367\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_186_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBDIR_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101111101010000"
        )
    port map (
            in0 => \N__4240\,
            in1 => \_gnd_net_\,
            in2 => \N__4145\,
            in3 => \N__4132\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8679\,
            ce => 'H',
            sr => \N__10976\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6161\,
            in2 => \_gnd_net_\,
            in3 => \N__4523\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_i_i_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4396\,
            in2 => \_gnd_net_\,
            in3 => \N__6363\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8684\,
            ce => \N__4280\,
            sr => \N__10972\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111100011111010"
        )
    port map (
            in0 => \N__4108\,
            in1 => \N__5076\,
            in2 => \N__4337\,
            in3 => \N__5023\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8688\,
            ce => 'H',
            sr => \N__10967\
        );

    \pll_RNI8MQ3_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5077\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__4349\,
            in1 => \N__4484\,
            in2 => \N__4046\,
            in3 => \N__4598\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8672\,
            ce => \N__4450\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIS5012_1_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4361\,
            in1 => \N__6723\,
            in2 => \_gnd_net_\,
            in3 => \N__5902\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_a2_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINE0O4_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111010101"
        )
    port map (
            in0 => \N__7533\,
            in1 => \N__6368\,
            in2 => \N__4193\,
            in3 => \N__6470\,
            lcout => \U712_CHIP_RAM.N_265\,
            ltout => \U712_CHIP_RAM.N_265_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIMBRQ8_3_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__4367\,
            in1 => \_gnd_net_\,
            in2 => \N__4190\,
            in3 => \N__4887\,
            lcout => \U712_CHIP_RAM.N_236\,
            ltout => \U712_CHIP_RAM.N_236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__4970\,
            in1 => \N__4187\,
            in2 => \N__4181\,
            in3 => \N__5228\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8672\,
            ce => \N__4450\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6551\,
            in1 => \N__5903\,
            in2 => \N__4892\,
            in3 => \N__6724\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER15\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIH4474_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6078\,
            in2 => \N__4178\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_426\,
            ltout => \U712_CHIP_RAM.N_426_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNIQ2RS7_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__5431\,
            in1 => \N__6366\,
            in2 => \N__4175\,
            in3 => \N__4408\,
            lcout => \U712_CHIP_RAM.N_328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__4565\,
            in1 => \N__4712\,
            in2 => \N__4397\,
            in3 => \N__7982\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8675\,
            ce => \N__4259\,
            sr => \N__10973\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011111000"
        )
    port map (
            in0 => \N__4205\,
            in1 => \N__7515\,
            in2 => \N__6092\,
            in3 => \N__5435\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIIE53C_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__4505\,
            in1 => \N__4549\,
            in2 => \_gnd_net_\,
            in3 => \N__4654\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__7339\,
            in1 => \_gnd_net_\,
            in2 => \N__4283\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ6QH5_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6361\,
            in1 => \N__4588\,
            in2 => \_gnd_net_\,
            in3 => \N__4516\,
            lcout => \U712_CHIP_RAM.N_350\,
            ltout => \U712_CHIP_RAM.N_350_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__4274\,
            in1 => \N__6362\,
            in2 => \N__4265\,
            in3 => \N__6469\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10996\,
            in1 => \_gnd_net_\,
            in2 => \N__4262\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__4211\,
            in1 => \N__7516\,
            in2 => \N__6882\,
            in3 => \N__4247\,
            lcout => \WRITE_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__4241\,
            in1 => \N__6935\,
            in2 => \_gnd_net_\,
            in3 => \N__6079\,
            lcout => \U712_CHIP_RAM.N_287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_5_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6761\,
            in1 => \N__9321\,
            in2 => \N__6619\,
            in3 => \N__6848\,
            lcout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4199\,
            in2 => \_gnd_net_\,
            in3 => \N__4849\,
            lcout => \U712_CHIP_RAM.un3_DMA_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4850\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7532\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7531\,
            in2 => \_gnd_net_\,
            in3 => \N__4333\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7529\,
            in1 => \N__5072\,
            in2 => \_gnd_net_\,
            in3 => \N__5027\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__7530\,
            in1 => \_gnd_net_\,
            in2 => \N__4319\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4332\,
            in2 => \_gnd_net_\,
            in3 => \N__4315\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__7528\,
            in1 => \N__4700\,
            in2 => \_gnd_net_\,
            in3 => \N__5107\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8691\,
            ce => \N__4667\,
            sr => \N__10949\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__10843\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9385\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111110"
        )
    port map (
            in0 => \N__6764\,
            in1 => \N__5817\,
            in2 => \N__6620\,
            in3 => \N__6364\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111111"
        )
    port map (
            in0 => \N__6460\,
            in1 => \_gnd_net_\,
            in2 => \N__4286\,
            in3 => \N__7527\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011101010"
        )
    port map (
            in0 => \N__5818\,
            in1 => \N__6765\,
            in2 => \N__5954\,
            in3 => \N__6608\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_129_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6435\,
            in1 => \N__4355\,
            in2 => \_gnd_net_\,
            in3 => \N__6155\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__6359\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5896\,
            lcout => \U712_CHIP_RAM.N_300\,
            ltout => \U712_CHIP_RAM.N_300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100101"
        )
    port map (
            in0 => \N__6720\,
            in1 => \_gnd_net_\,
            in2 => \N__4370\,
            in3 => \N__6548\,
            lcout => \U712_CHIP_RAM.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIGGM16_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__6095\,
            in1 => \N__6132\,
            in2 => \N__4604\,
            in3 => \N__4904\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_0_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5798\,
            in1 => \N__5895\,
            in2 => \N__6468\,
            in3 => \N__6719\,
            lcout => \U712_CHIP_RAM.N_437\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNIUL431_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111100"
        )
    port map (
            in0 => \N__5448\,
            in1 => \N__6544\,
            in2 => \N__6891\,
            in3 => \N__5796\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_esr_RNIULZ0Z431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100011001100"
        )
    port map (
            in0 => \N__5797\,
            in1 => \N__6718\,
            in2 => \N__6592\,
            in3 => \N__5894\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5799\,
            in2 => \_gnd_net_\,
            in3 => \N__6425\,
            lcout => \U712_CHIP_RAM.N_381\,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5930\,
            in2 => \_gnd_net_\,
            in3 => \N__4343\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4485\,
            in1 => \N__6585\,
            in2 => \_gnd_net_\,
            in3 => \N__4340\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \N__8673\,
            ce => \N__4454\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4481\,
            in1 => \N__6754\,
            in2 => \_gnd_net_\,
            in3 => \N__4499\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__8673\,
            ce => \N__4454\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4486\,
            in1 => \N__4922\,
            in2 => \_gnd_net_\,
            in3 => \N__4496\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__8673\,
            ce => \N__4454\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4482\,
            in1 => \N__4949\,
            in2 => \_gnd_net_\,
            in3 => \N__4493\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__8673\,
            ce => \N__4454\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4487\,
            in1 => \N__4961\,
            in2 => \_gnd_net_\,
            in3 => \N__4490\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__8673\,
            ce => \N__4454\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4483\,
            in1 => \N__4936\,
            in2 => \_gnd_net_\,
            in3 => \N__4457\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8673\,
            ce => \N__4454\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__5156\,
            in1 => \N__4418\,
            in2 => \N__6467\,
            in3 => \N__5838\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__5201\,
            in1 => \N__5128\,
            in2 => \N__4427\,
            in3 => \N__4612\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8676\,
            ce => 'H',
            sr => \N__10963\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__5953\,
            in1 => \N__4424\,
            in2 => \_gnd_net_\,
            in3 => \N__4883\,
            lcout => \U712_CHIP_RAM.N_348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__5442\,
            in1 => \N__4412\,
            in2 => \_gnd_net_\,
            in3 => \N__4392\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_76_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111101001110"
        )
    port map (
            in0 => \N__4613\,
            in1 => \N__4627\,
            in2 => \N__4658\,
            in3 => \N__4655\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8676\,
            ce => 'H',
            sr => \N__10963\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__5952\,
            in1 => \N__6360\,
            in2 => \_gnd_net_\,
            in3 => \N__4882\,
            lcout => \U712_CHIP_RAM.N_438\,
            ltout => \U712_CHIP_RAM.N_438_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6609\,
            in1 => \N__6857\,
            in2 => \N__4616\,
            in3 => \N__6753\,
            lcout => \U712_CHIP_RAM.N_336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIVLD65_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6069\,
            in1 => \N__4599\,
            in2 => \N__6128\,
            in3 => \N__4532\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011001100"
        )
    port map (
            in0 => \N__4538\,
            in1 => \N__9341\,
            in2 => \N__4553\,
            in3 => \N__4550\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8681\,
            ce => 'H',
            sr => \N__10955\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__6763\,
            in1 => \N__6600\,
            in2 => \_gnd_net_\,
            in3 => \N__6847\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5145\,
            in2 => \_gnd_net_\,
            in3 => \N__5325\,
            lcout => \U712_CHIP_RAM.N_247\,
            ltout => \U712_CHIP_RAM.N_247_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIR9VE1_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6115\,
            in2 => \N__4526\,
            in3 => \N__6068\,
            lcout => \U712_CHIP_RAM.N_244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIOVA11_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6846\,
            in1 => \N__6762\,
            in2 => \_gnd_net_\,
            in3 => \N__6596\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_1_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5345\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8681\,
            ce => 'H',
            sr => \N__10955\
        );

    \U712_REG_SM.C3_SYNC_1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5264\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8686\,
            ce => 'H',
            sr => \N__10950\
        );

    \U712_REG_SM.C3_SYNC_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8686\,
            ce => 'H',
            sr => \N__10950\
        );

    \DBR_SYNC_0_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4766\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8686\,
            ce => 'H',
            sr => \N__10950\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010001010000"
        )
    port map (
            in0 => \N__5016\,
            in1 => \N__4699\,
            in2 => \N__4688\,
            in3 => \N__4736\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8686\,
            ce => 'H',
            sr => \N__10950\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9965\,
            in2 => \_gnd_net_\,
            in3 => \N__4730\,
            lcout => \U712_CHIP_RAM.BANK0_9_u_0_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5580\,
            in2 => \_gnd_net_\,
            in3 => \N__5129\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__7476\,
            in1 => \N__4684\,
            in2 => \N__4673\,
            in3 => \N__5102\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_269_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10994\,
            in1 => \_gnd_net_\,
            in2 => \N__4670\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.N_269_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__10776\,
            in1 => \N__7383\,
            in2 => \_gnd_net_\,
            in3 => \N__10715\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8692\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0_0_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5496\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5455\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.N_249_i_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__10787\,
            in1 => \N__10701\,
            in2 => \_gnd_net_\,
            in3 => \N__6892\,
            lcout => \N_249_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__6365\,
            in1 => \N__6773\,
            in2 => \_gnd_net_\,
            in3 => \N__5843\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_0_1_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101010111010"
        )
    port map (
            in0 => \N__4820\,
            in1 => \N__6884\,
            in2 => \N__4814\,
            in3 => \N__5960\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8665\,
            ce => \N__5650\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIIPOI5_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6093\,
            in1 => \N__4903\,
            in2 => \N__6134\,
            in3 => \N__6013\,
            lcout => \U712_CHIP_RAM.N_325\,
            ltout => \U712_CHIP_RAM.N_325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNI0N6TH_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__7522\,
            in1 => \N__4993\,
            in2 => \N__4811\,
            in3 => \N__5221\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_5_1_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__6736\,
            in1 => \N__7526\,
            in2 => \N__6601\,
            in3 => \N__5937\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011010000"
        )
    port map (
            in0 => \N__5938\,
            in1 => \N__5822\,
            in2 => \N__6602\,
            in3 => \N__6737\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6567\,
            in1 => \N__5939\,
            in2 => \N__4891\,
            in3 => \N__6157\,
            lcout => \U712_CHIP_RAM.N_317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__4994\,
            in1 => \N__5220\,
            in2 => \N__7535\,
            in3 => \N__4982\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__6002\,
            in1 => \_gnd_net_\,
            in2 => \N__4973\,
            in3 => \N__9034\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8669\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__5722\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5823\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4960\,
            in1 => \N__4948\,
            in2 => \N__4937\,
            in3 => \N__4921\,
            lcout => \U712_CHIP_RAM.N_241\,
            ltout => \U712_CHIP_RAM.N_241_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4GV43_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__6721\,
            in1 => \N__6549\,
            in2 => \N__4910\,
            in3 => \N__6310\,
            lcout => \U712_CHIP_RAM.N_386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7521\,
            in2 => \_gnd_net_\,
            in3 => \N__6293\,
            lcout => \U712_CHIP_RAM.N_388\,
            ltout => \U712_CHIP_RAM.N_388_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIHHIB1_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5150\,
            in2 => \N__4907\,
            in3 => \N__5332\,
            lcout => \U712_CHIP_RAM.N_325_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6550\,
            in1 => \N__6722\,
            in2 => \_gnd_net_\,
            in3 => \N__4878\,
            lcout => \U712_CHIP_RAM.N_434\,
            ltout => \U712_CHIP_RAM.N_434_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3DQ77_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__5955\,
            in1 => \N__5237\,
            in2 => \N__5231\,
            in3 => \N__6311\,
            lcout => \U712_CHIP_RAM.N_439\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__5207\,
            in1 => \N__6294\,
            in2 => \_gnd_net_\,
            in3 => \N__6443\,
            lcout => \U712_CHIP_RAM.N_335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5195\,
            in1 => \N__5177\,
            in2 => \_gnd_net_\,
            in3 => \N__9054\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_6_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9339\,
            in2 => \_gnd_net_\,
            in3 => \N__6867\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6752\,
            in1 => \N__6584\,
            in2 => \N__5159\,
            in3 => \N__5958\,
            lcout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__5354\,
            in1 => \N__9340\,
            in2 => \N__7534\,
            in3 => \N__5149\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8674\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010110000"
        )
    port map (
            in0 => \N__7193\,
            in1 => \N__7604\,
            in2 => \N__7520\,
            in3 => \N__7544\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8677\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011111"
        )
    port map (
            in0 => \N__5587\,
            in1 => \N__5127\,
            in2 => \N__5108\,
            in3 => \N__5015\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_351_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__5106\,
            in1 => \N__7481\,
            in2 => \N__5081\,
            in3 => \N__5078\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8677\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_o2_1_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__5262\,
            in1 => \N__5344\,
            in2 => \N__5333\,
            in3 => \N__5283\,
            lcout => \U712_REG_SM.m17_i_0_o2_1\,
            ltout => \U712_REG_SM.m17_i_0_o2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_m2_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__5284\,
            in1 => \N__7036\,
            in2 => \N__5309\,
            in3 => \N__5263\,
            lcout => \U712_REG_SM.N_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5306\,
            in1 => \N__9320\,
            in2 => \_gnd_net_\,
            in3 => \N__9512\,
            lcout => \U712_CHIP_RAM.N_392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI7UAP_1_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5260\,
            in2 => \_gnd_net_\,
            in3 => \N__5282\,
            lcout => \U712_REG_SM.C3_SYNC_RNI7UAPZ0Z_1\,
            ltout => \U712_REG_SM.C3_SYNC_RNI7UAPZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__7043\,
            in1 => \N__6206\,
            in2 => \N__5288\,
            in3 => \N__7703\,
            lcout => \U712_REG_SM.N_360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7160\,
            in2 => \_gnd_net_\,
            in3 => \N__7041\,
            lcout => \U712_REG_SM.N_270_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_0_0_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6952\,
            in2 => \_gnd_net_\,
            in3 => \N__6978\,
            lcout => OPEN,
            ltout => \U712_REG_SM.m15_i_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_0_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5285\,
            in1 => \N__5261\,
            in2 => \N__5240\,
            in3 => \N__7042\,
            lcout => \U712_REG_SM.N_359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000101010"
        )
    port map (
            in0 => \N__7044\,
            in1 => \N__6934\,
            in2 => \N__7166\,
            in3 => \N__6998\,
            lcout => \U712_REG_SM.REG_TACK_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_ns_1_0__m15_i_0_a2_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001001100"
        )
    port map (
            in0 => \N__6979\,
            in1 => \N__7164\,
            in2 => \N__6956\,
            in3 => \N__5627\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__7477\,
            in1 => \N__5611\,
            in2 => \N__5621\,
            in3 => \N__5618\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__5612\,
            in1 => \N__5600\,
            in2 => \N__5588\,
            in3 => \N__5594\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8687\,
            ce => 'H',
            sr => \N__10940\
        );

    \U712_REG_SM.C1_SYNC_0_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5564\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8687\,
            ce => 'H',
            sr => \N__10940\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10826\,
            in2 => \_gnd_net_\,
            in3 => \N__6201\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_340_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__7382\,
            in1 => \N__5402\,
            in2 => \N__5525\,
            in3 => \N__5522\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8690\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5497\,
            in2 => \_gnd_net_\,
            in3 => \N__5456\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5401\,
            in2 => \_gnd_net_\,
            in3 => \N__5375\,
            lcout => \U712_CHIP_RAM.N_345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__9441\,
            in1 => \N__10540\,
            in2 => \_gnd_net_\,
            in3 => \N__10460\,
            lcout => \U712_BYTE_ENABLE.N_370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__10632\,
            in1 => \N__10459\,
            in2 => \N__10170\,
            in3 => \N__9440\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_374_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_51_i_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__8341\,
            in1 => \N__7957\,
            in2 => \N__5753\,
            in3 => \N__10714\,
            lcout => \N_51_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_10_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5702\,
            in1 => \N__5687\,
            in2 => \_gnd_net_\,
            in3 => \N__9069\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011011010"
        )
    port map (
            in0 => \N__5841\,
            in1 => \N__6776\,
            in2 => \N__6628\,
            in3 => \N__5959\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_i_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6465\,
            in2 => \N__5669\,
            in3 => \N__7518\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8660\,
            ce => \N__5654\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6349\,
            in1 => \N__6621\,
            in2 => \_gnd_net_\,
            in3 => \N__5842\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__7519\,
            in1 => \N__6466\,
            in2 => \N__5666\,
            in3 => \N__5663\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8660\,
            ce => \N__5654\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8260\,
            in1 => \N__9008\,
            in2 => \_gnd_net_\,
            in3 => \N__8200\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_4_1_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6156\,
            in1 => \N__6133\,
            in2 => \_gnd_net_\,
            in3 => \N__6094\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_7_1_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__6774\,
            in1 => \N__6618\,
            in2 => \_gnd_net_\,
            in3 => \N__5957\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_271_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_6_1_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7517\,
            in2 => \N__6041\,
            in3 => \N__6348\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_a2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__6038\,
            in1 => \N__5839\,
            in2 => \N__6032\,
            in3 => \N__6442\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_59_i_a2_i_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__6029\,
            in1 => \N__6023\,
            in2 => \N__6017\,
            in3 => \N__6014\,
            lcout => \U712_CHIP_RAM.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9009\,
            in1 => \N__5996\,
            in2 => \_gnd_net_\,
            in3 => \N__5975\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6883\,
            in2 => \_gnd_net_\,
            in3 => \N__6604\,
            lcout => \U712_CHIP_RAM.CLK_EN_5_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_2_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111111111"
        )
    port map (
            in0 => \N__6766\,
            in1 => \N__6603\,
            in2 => \_gnd_net_\,
            in3 => \N__5956\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__6326\,
            in1 => \N__5840\,
            in2 => \N__5756\,
            in3 => \N__6464\,
            lcout => \U712_CHIP_RAM.N_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__6775\,
            in1 => \N__6641\,
            in2 => \N__6629\,
            in3 => \N__6453\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__7495\,
            in1 => \_gnd_net_\,
            in2 => \N__6371\,
            in3 => \N__6327\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8671\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6242\,
            in1 => \N__6224\,
            in2 => \_gnd_net_\,
            in3 => \N__9053\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNIC74N_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6205\,
            in2 => \_gnd_net_\,
            in3 => \N__7702\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_360_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI8VBS1_0_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6178\,
            in1 => \N__7159\,
            in2 => \N__6182\,
            in3 => \N__7037\,
            lcout => \U712_REG_SM.ASn_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__7040\,
            in1 => \N__7446\,
            in2 => \N__7130\,
            in3 => \N__6999\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_o2_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__6950\,
            in1 => \N__7155\,
            in2 => \N__6179\,
            in3 => \N__6977\,
            lcout => \U712_REG_SM.m17_i_0_o2\,
            ltout => \U712_REG_SM.m17_i_0_o2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__7039\,
            in1 => \_gnd_net_\,
            in2 => \N__6167\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U712_REG_SM.REG_CYCLE_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011000100"
        )
    port map (
            in0 => \N__7445\,
            in1 => \N__10816\,
            in2 => \N__6164\,
            in3 => \N__7118\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_ns_1_0__m17_i_0_a2_0_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6976\,
            in1 => \N__6951\,
            in2 => \N__7165\,
            in3 => \N__7136\,
            lcout => \U712_REG_SM.N_435\,
            ltout => \U712_REG_SM.N_435_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7121\,
            in3 => \N__7038\,
            lcout => \U712_REG_SM.N_363\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__7074\,
            in1 => \N__7060\,
            in2 => \N__7051\,
            in3 => \N__7000\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8683\,
            ce => 'H',
            sr => \N__10938\
        );

    \U712_REG_SM.DS_EN_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001110"
        )
    port map (
            in0 => \N__10192\,
            in1 => \N__7061\,
            in2 => \N__7052\,
            in3 => \N__7001\,
            lcout => \DS_ENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8683\,
            ce => 'H',
            sr => \N__10938\
        );

    \U712_REG_SM.C1_SYNC_1_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6980\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8683\,
            ce => 'H',
            sr => \N__10938\
        );

    \U712_BUFFERS.DRDDIR_0_m2_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__6930\,
            in1 => \N__10839\,
            in2 => \_gnd_net_\,
            in3 => \N__6893\,
            lcout => \N_276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9454\,
            in1 => \N__6782\,
            in2 => \N__9114\,
            in3 => \N__8018\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8247\,
            in1 => \N__8204\,
            in2 => \N__8165\,
            in3 => \N__9073\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7292\,
            in1 => \N__7271\,
            in2 => \_gnd_net_\,
            in3 => \N__9060\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9061\,
            in1 => \N__9413\,
            in2 => \N__7250\,
            in3 => \N__10328\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111011100000111"
        )
    port map (
            in0 => \N__7247\,
            in1 => \N__9456\,
            in2 => \N__7241\,
            in3 => \N__7213\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8666\,
            ce => 'H',
            sr => \N__10951\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7583\,
            in2 => \_gnd_net_\,
            in3 => \N__7202\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__7694\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7556\,
            in2 => \_gnd_net_\,
            in3 => \N__7199\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__7694\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7595\,
            in2 => \_gnd_net_\,
            in3 => \N__7196\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__7694\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7189\,
            in2 => \_gnd_net_\,
            in3 => \N__7175\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__7694\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7570\,
            in2 => \_gnd_net_\,
            in3 => \N__7172\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__7694\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7616\,
            in2 => \_gnd_net_\,
            in3 => \N__7169\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__7694\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7628\,
            in2 => \_gnd_net_\,
            in3 => \N__7709\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__7694\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7640\,
            in2 => \_gnd_net_\,
            in3 => \N__7706\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7694\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7639\,
            in1 => \N__7627\,
            in2 => \_gnd_net_\,
            in3 => \N__7615\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__7594\,
            in1 => \N__7582\,
            in2 => \N__7571\,
            in3 => \N__7555\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7381\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7298\,
            in1 => \N__7862\,
            in2 => \_gnd_net_\,
            in3 => \N__7313\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8655\,
            ce => \N__8546\,
            sr => \N__10962\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100101111"
        )
    port map (
            in0 => \N__8033\,
            in1 => \N__8825\,
            in2 => \N__9102\,
            in3 => \N__9443\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000101"
        )
    port map (
            in0 => \N__8166\,
            in1 => \N__8262\,
            in2 => \N__8224\,
            in3 => \N__9074\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8261\,
            in2 => \_gnd_net_\,
            in3 => \N__8219\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011110000"
        )
    port map (
            in0 => \N__9442\,
            in1 => \N__8032\,
            in2 => \N__7865\,
            in3 => \N__9078\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__9059\,
            in1 => \N__8826\,
            in2 => \_gnd_net_\,
            in3 => \N__7856\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7844\,
            in1 => \N__7832\,
            in2 => \_gnd_net_\,
            in3 => \N__9058\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__8762\,
            in1 => \N__7810\,
            in2 => \N__8501\,
            in3 => \N__9452\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011111111"
        )
    port map (
            in0 => \N__7811\,
            in1 => \N__8497\,
            in2 => \N__9470\,
            in3 => \N__8763\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7787\,
            in1 => \N__7781\,
            in2 => \_gnd_net_\,
            in3 => \N__7775\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8659\,
            ce => \N__8576\,
            sr => \N__10943\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7748\,
            in1 => \N__7733\,
            in2 => \_gnd_net_\,
            in3 => \N__9103\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9104\,
            in1 => \N__9455\,
            in2 => \N__7712\,
            in3 => \N__8006\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9958\,
            in1 => \N__8414\,
            in2 => \_gnd_net_\,
            in3 => \N__8482\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__9675\,
            sr => \N__10937\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8483\,
            in1 => \N__9959\,
            in2 => \_gnd_net_\,
            in3 => \N__9584\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__9675\,
            sr => \N__10937\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8480\,
            in1 => \N__9957\,
            in2 => \_gnd_net_\,
            in3 => \N__8413\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9711\,
            ce => \N__9673\,
            sr => \N__10935\
        );

    \U712_CHIP_RAM.DMA_A20_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__8000\,
            in1 => \N__9947\,
            in2 => \N__9783\,
            in3 => \N__7975\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__10934\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__10619\,
            in1 => \N__10161\,
            in2 => \N__9476\,
            in3 => \N__10468\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_369_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_55_i_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__9496\,
            in1 => \N__7961\,
            in2 => \N__7946\,
            in3 => \N__10700\,
            lcout => \N_55_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_13_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8223\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8654\,
            ce => 'H',
            sr => \N__10977\
        );

    \U712_CHIP_RAM.CRCSn_LC_13_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8174\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8656\,
            ce => 'H',
            sr => \N__10974\
        );

    \U712_CHIP_RAM.RASn_LC_13_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8270\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8656\,
            ce => 'H',
            sr => \N__10974\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8269\,
            in1 => \N__9111\,
            in2 => \N__8225\,
            in3 => \N__8173\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8658\,
            ce => \N__8547\,
            sr => \N__10964\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10995\,
            in2 => \_gnd_net_\,
            in3 => \N__8120\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9448\,
            in1 => \N__8114\,
            in2 => \N__9095\,
            in3 => \N__8435\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9447\,
            in2 => \_gnd_net_\,
            in3 => \N__9062\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8895\,
            in1 => \N__8108\,
            in2 => \N__8867\,
            in3 => \N__8099\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8667\,
            ce => \N__8563\,
            sr => \N__10952\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__8856\,
            in1 => \N__8896\,
            in2 => \N__8447\,
            in3 => \N__8039\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8667\,
            ce => \N__8563\,
            sr => \N__10952\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9460\,
            in1 => \N__8060\,
            in2 => \N__9115\,
            in3 => \N__8357\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9461\,
            in1 => \N__8051\,
            in2 => \N__9116\,
            in3 => \N__8423\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9950\,
            in1 => \N__8412\,
            in2 => \_gnd_net_\,
            in3 => \N__10304\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9712\,
            ce => \N__9677\,
            sr => \N__10941\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9620\,
            in1 => \_gnd_net_\,
            in2 => \N__9964\,
            in3 => \N__10064\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9712\,
            ce => \N__9677\,
            sr => \N__10941\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__9583\,
            in1 => \_gnd_net_\,
            in2 => \N__9963\,
            in3 => \N__8481\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9712\,
            ce => \N__9677\,
            sr => \N__10941\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9949\,
            in1 => \N__10057\,
            in2 => \_gnd_net_\,
            in3 => \N__9616\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__9676\,
            sr => \N__10939\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9615\,
            in1 => \N__9948\,
            in2 => \_gnd_net_\,
            in3 => \N__9581\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__9676\,
            sr => \N__10939\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8402\,
            in1 => \N__10300\,
            in2 => \_gnd_net_\,
            in3 => \N__9946\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9674\,
            sr => \N__10936\
        );

    \U712_BYTE_ENABLE.N_53_i_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000111111"
        )
    port map (
            in0 => \N__10780\,
            in1 => \N__8309\,
            in2 => \N__9475\,
            in3 => \N__8348\,
            lcout => \N_53_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LMBE_0_o2_i_o2_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000101111"
        )
    port map (
            in0 => \N__10633\,
            in1 => \N__10178\,
            in2 => \N__10472\,
            in3 => \N__10544\,
            lcout => \U712_BYTE_ENABLE.N_303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_0_o2_i_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110100000"
        )
    port map (
            in0 => \N__10620\,
            in1 => \N__10179\,
            in2 => \N__10461\,
            in3 => \N__10524\,
            lcout => \UMBE_0_o2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_i_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10621\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10180\,
            lcout => \U712_BYTE_ENABLE_UUBE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_14_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9112\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8657\,
            ce => 'H',
            sr => \N__10978\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8900\,
            in1 => \N__9521\,
            in2 => \N__8868\,
            in3 => \N__9188\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8661\,
            ce => \N__8570\,
            sr => \N__10968\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8770\,
            in1 => \N__9161\,
            in2 => \N__9469\,
            in3 => \N__10373\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8661\,
            ce => \N__8570\,
            sr => \N__10968\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9453\,
            in1 => \N__9125\,
            in2 => \N__9113\,
            in3 => \N__9638\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__8863\,
            in1 => \N__8897\,
            in2 => \N__8942\,
            in3 => \N__9977\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8668\,
            ce => \N__8572\,
            sr => \N__10965\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8898\,
            in1 => \N__9629\,
            in2 => \N__8869\,
            in3 => \N__8924\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8668\,
            ce => \N__8572\,
            sr => \N__10965\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__10223\,
            in1 => \N__8899\,
            in2 => \N__8870\,
            in3 => \N__8795\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8670\,
            ce => \N__8571\,
            sr => \N__10956\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8771\,
            in1 => \N__8738\,
            in2 => \N__9474\,
            in3 => \N__9722\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8670\,
            ce => \N__8571\,
            sr => \N__10956\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__9863\,
            in1 => \_gnd_net_\,
            in2 => \N__10019\,
            in3 => \N__10363\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__9681\,
            sr => \N__10953\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10362\,
            in1 => \N__10015\,
            in2 => \_gnd_net_\,
            in3 => \N__9907\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9710\,
            ce => \N__9679\,
            sr => \N__10944\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9614\,
            in1 => \N__9906\,
            in2 => \_gnd_net_\,
            in3 => \N__9582\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9710\,
            ce => \N__9679\,
            sr => \N__10944\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10014\,
            in1 => \N__9905\,
            in2 => \_gnd_net_\,
            in3 => \N__10056\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__9678\,
            sr => \N__10942\
        );

    \U712_BYTE_ENABLE.N_57_i_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__10772\,
            in1 => \N__9497\,
            in2 => \N__9251\,
            in3 => \N__9468\,
            lcout => \N_57_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_0_a2_0_a2_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__10177\,
            in1 => \N__10634\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_BYTE_ENABLE.UUBE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_0_o2_i_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100101010"
        )
    port map (
            in0 => \N__10539\,
            in1 => \N__10583\,
            in2 => \N__10181\,
            in3 => \N__10453\,
            lcout => \N_185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100001111"
        )
    port map (
            in0 => \N__10452\,
            in1 => \N__10175\,
            in2 => \N__10210\,
            in3 => \N__10528\,
            lcout => \N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_303_i_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110110000"
        )
    port map (
            in0 => \N__10174\,
            in1 => \N__10628\,
            in2 => \N__10538\,
            in3 => \N__10451\,
            lcout => \N_303_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9785\,
            in1 => \N__9944\,
            in2 => \_gnd_net_\,
            in3 => \N__10364\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9713\,
            ce => \N__9685\,
            sr => \N__10966\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9862\,
            in1 => \N__9784\,
            in2 => \_gnd_net_\,
            in3 => \N__10361\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__9683\,
            sr => \N__10957\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10250\,
            in1 => \N__9904\,
            in2 => \_gnd_net_\,
            in3 => \N__10299\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__9682\,
            sr => \N__10954\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9903\,
            in1 => \N__10281\,
            in2 => \_gnd_net_\,
            in3 => \N__10246\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9707\,
            ce => \N__9680\,
            sr => \N__10945\
        );

    \U712_BYTE_ENABLE.N_337_i_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__10214\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10176\,
            lcout => \N_337_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10055\,
            in1 => \N__9911\,
            in2 => \_gnd_net_\,
            in3 => \N__10004\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9708\,
            ce => \N__9684\,
            sr => \N__10958\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9945\,
            in1 => \N__9800\,
            in2 => \_gnd_net_\,
            in3 => \N__9765\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9709\,
            ce => \N__9686\,
            sr => \N__10975\
        );

    \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__10847\,
            in1 => \N__10768\,
            in2 => \_gnd_net_\,
            in3 => \N__10688\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

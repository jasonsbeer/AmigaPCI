// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 13 2025 12:13:37

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U400_TOP" view "INTERFACE"

module U400_TOP (
    SIZ,
    MA,
    A,
    LBENn,
    CS0n,
    UUBEn,
    TAn,
    CLK40,
    RnW,
    BANK1,
    UMBEn,
    WEn,
    LLBEn,
    TSn,
    LMBEn,
    RASn,
    CS1n,
    RESETn,
    CLK_EN,
    CASn,
    BANK0);

    input [1:0] SIZ;
    output [12:0] MA;
    input [31:0] A;
    output LBENn;
    output CS0n;
    output UUBEn;
    output TAn;
    input CLK40;
    input RnW;
    output BANK1;
    output UMBEn;
    output WEn;
    output LLBEn;
    input TSn;
    output LMBEn;
    output RASn;
    output CS1n;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;

    wire N__7451;
    wire N__7450;
    wire N__7449;
    wire N__7442;
    wire N__7441;
    wire N__7440;
    wire N__7433;
    wire N__7432;
    wire N__7431;
    wire N__7424;
    wire N__7423;
    wire N__7422;
    wire N__7415;
    wire N__7414;
    wire N__7413;
    wire N__7406;
    wire N__7405;
    wire N__7404;
    wire N__7397;
    wire N__7396;
    wire N__7395;
    wire N__7388;
    wire N__7387;
    wire N__7386;
    wire N__7379;
    wire N__7378;
    wire N__7377;
    wire N__7370;
    wire N__7369;
    wire N__7368;
    wire N__7361;
    wire N__7360;
    wire N__7359;
    wire N__7352;
    wire N__7351;
    wire N__7350;
    wire N__7343;
    wire N__7342;
    wire N__7341;
    wire N__7334;
    wire N__7333;
    wire N__7332;
    wire N__7325;
    wire N__7324;
    wire N__7323;
    wire N__7316;
    wire N__7315;
    wire N__7314;
    wire N__7307;
    wire N__7306;
    wire N__7305;
    wire N__7298;
    wire N__7297;
    wire N__7296;
    wire N__7289;
    wire N__7288;
    wire N__7287;
    wire N__7280;
    wire N__7279;
    wire N__7278;
    wire N__7271;
    wire N__7270;
    wire N__7269;
    wire N__7262;
    wire N__7261;
    wire N__7260;
    wire N__7253;
    wire N__7252;
    wire N__7251;
    wire N__7244;
    wire N__7243;
    wire N__7242;
    wire N__7235;
    wire N__7234;
    wire N__7233;
    wire N__7226;
    wire N__7225;
    wire N__7224;
    wire N__7217;
    wire N__7216;
    wire N__7215;
    wire N__7208;
    wire N__7207;
    wire N__7206;
    wire N__7199;
    wire N__7198;
    wire N__7197;
    wire N__7190;
    wire N__7189;
    wire N__7188;
    wire N__7181;
    wire N__7180;
    wire N__7179;
    wire N__7172;
    wire N__7171;
    wire N__7170;
    wire N__7163;
    wire N__7162;
    wire N__7161;
    wire N__7154;
    wire N__7153;
    wire N__7152;
    wire N__7145;
    wire N__7144;
    wire N__7143;
    wire N__7136;
    wire N__7135;
    wire N__7134;
    wire N__7127;
    wire N__7126;
    wire N__7125;
    wire N__7118;
    wire N__7117;
    wire N__7116;
    wire N__7109;
    wire N__7108;
    wire N__7107;
    wire N__7100;
    wire N__7099;
    wire N__7098;
    wire N__7091;
    wire N__7090;
    wire N__7089;
    wire N__7082;
    wire N__7081;
    wire N__7080;
    wire N__7073;
    wire N__7072;
    wire N__7071;
    wire N__7064;
    wire N__7063;
    wire N__7062;
    wire N__7055;
    wire N__7054;
    wire N__7053;
    wire N__7046;
    wire N__7045;
    wire N__7044;
    wire N__7037;
    wire N__7036;
    wire N__7035;
    wire N__7028;
    wire N__7027;
    wire N__7026;
    wire N__7019;
    wire N__7018;
    wire N__7017;
    wire N__7010;
    wire N__7009;
    wire N__7008;
    wire N__7001;
    wire N__7000;
    wire N__6999;
    wire N__6992;
    wire N__6991;
    wire N__6990;
    wire N__6983;
    wire N__6982;
    wire N__6981;
    wire N__6974;
    wire N__6973;
    wire N__6972;
    wire N__6965;
    wire N__6964;
    wire N__6963;
    wire N__6956;
    wire N__6955;
    wire N__6954;
    wire N__6947;
    wire N__6946;
    wire N__6945;
    wire N__6938;
    wire N__6937;
    wire N__6936;
    wire N__6929;
    wire N__6928;
    wire N__6927;
    wire N__6920;
    wire N__6919;
    wire N__6918;
    wire N__6911;
    wire N__6910;
    wire N__6909;
    wire N__6902;
    wire N__6901;
    wire N__6900;
    wire N__6893;
    wire N__6892;
    wire N__6891;
    wire N__6884;
    wire N__6883;
    wire N__6882;
    wire N__6875;
    wire N__6874;
    wire N__6873;
    wire N__6856;
    wire N__6853;
    wire N__6850;
    wire N__6847;
    wire N__6846;
    wire N__6845;
    wire N__6844;
    wire N__6843;
    wire N__6842;
    wire N__6841;
    wire N__6840;
    wire N__6839;
    wire N__6836;
    wire N__6835;
    wire N__6834;
    wire N__6827;
    wire N__6824;
    wire N__6823;
    wire N__6822;
    wire N__6821;
    wire N__6818;
    wire N__6813;
    wire N__6810;
    wire N__6807;
    wire N__6804;
    wire N__6801;
    wire N__6796;
    wire N__6793;
    wire N__6790;
    wire N__6787;
    wire N__6780;
    wire N__6777;
    wire N__6776;
    wire N__6773;
    wire N__6772;
    wire N__6771;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6757;
    wire N__6754;
    wire N__6753;
    wire N__6750;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6732;
    wire N__6727;
    wire N__6724;
    wire N__6721;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6691;
    wire N__6688;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6676;
    wire N__6673;
    wire N__6670;
    wire N__6667;
    wire N__6666;
    wire N__6665;
    wire N__6664;
    wire N__6663;
    wire N__6660;
    wire N__6659;
    wire N__6658;
    wire N__6649;
    wire N__6648;
    wire N__6645;
    wire N__6642;
    wire N__6639;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6616;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6597;
    wire N__6594;
    wire N__6593;
    wire N__6592;
    wire N__6589;
    wire N__6588;
    wire N__6585;
    wire N__6582;
    wire N__6581;
    wire N__6580;
    wire N__6579;
    wire N__6576;
    wire N__6573;
    wire N__6570;
    wire N__6569;
    wire N__6564;
    wire N__6561;
    wire N__6558;
    wire N__6555;
    wire N__6554;
    wire N__6547;
    wire N__6544;
    wire N__6535;
    wire N__6532;
    wire N__6527;
    wire N__6522;
    wire N__6517;
    wire N__6514;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6506;
    wire N__6505;
    wire N__6504;
    wire N__6503;
    wire N__6502;
    wire N__6501;
    wire N__6500;
    wire N__6497;
    wire N__6496;
    wire N__6495;
    wire N__6494;
    wire N__6493;
    wire N__6492;
    wire N__6491;
    wire N__6490;
    wire N__6489;
    wire N__6488;
    wire N__6487;
    wire N__6486;
    wire N__6483;
    wire N__6482;
    wire N__6481;
    wire N__6480;
    wire N__6479;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6402;
    wire N__6401;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6389;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6365;
    wire N__6362;
    wire N__6357;
    wire N__6352;
    wire N__6349;
    wire N__6348;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6309;
    wire N__6308;
    wire N__6307;
    wire N__6306;
    wire N__6305;
    wire N__6302;
    wire N__6301;
    wire N__6296;
    wire N__6293;
    wire N__6292;
    wire N__6289;
    wire N__6288;
    wire N__6287;
    wire N__6286;
    wire N__6283;
    wire N__6280;
    wire N__6277;
    wire N__6274;
    wire N__6271;
    wire N__6268;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6255;
    wire N__6244;
    wire N__6241;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6221;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6198;
    wire N__6197;
    wire N__6196;
    wire N__6195;
    wire N__6194;
    wire N__6189;
    wire N__6188;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6175;
    wire N__6172;
    wire N__6171;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6163;
    wire N__6160;
    wire N__6157;
    wire N__6154;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6140;
    wire N__6135;
    wire N__6132;
    wire N__6123;
    wire N__6122;
    wire N__6117;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6094;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__5998;
    wire N__5995;
    wire N__5992;
    wire N__5989;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5977;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5947;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5904;
    wire N__5903;
    wire N__5900;
    wire N__5897;
    wire N__5894;
    wire N__5887;
    wire N__5884;
    wire N__5881;
    wire N__5878;
    wire N__5875;
    wire N__5872;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5848;
    wire N__5845;
    wire N__5842;
    wire N__5841;
    wire N__5840;
    wire N__5839;
    wire N__5832;
    wire N__5829;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5815;
    wire N__5812;
    wire N__5811;
    wire N__5808;
    wire N__5805;
    wire N__5804;
    wire N__5803;
    wire N__5800;
    wire N__5795;
    wire N__5792;
    wire N__5789;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5773;
    wire N__5770;
    wire N__5767;
    wire N__5766;
    wire N__5765;
    wire N__5764;
    wire N__5761;
    wire N__5760;
    wire N__5759;
    wire N__5752;
    wire N__5749;
    wire N__5744;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5722;
    wire N__5721;
    wire N__5718;
    wire N__5713;
    wire N__5710;
    wire N__5709;
    wire N__5706;
    wire N__5705;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5676;
    wire N__5671;
    wire N__5670;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5632;
    wire N__5631;
    wire N__5628;
    wire N__5627;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5586;
    wire N__5585;
    wire N__5582;
    wire N__5581;
    wire N__5578;
    wire N__5577;
    wire N__5574;
    wire N__5569;
    wire N__5566;
    wire N__5565;
    wire N__5562;
    wire N__5561;
    wire N__5558;
    wire N__5553;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5535;
    wire N__5532;
    wire N__5529;
    wire N__5524;
    wire N__5523;
    wire N__5522;
    wire N__5521;
    wire N__5520;
    wire N__5519;
    wire N__5518;
    wire N__5517;
    wire N__5510;
    wire N__5503;
    wire N__5498;
    wire N__5491;
    wire N__5490;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5469;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5446;
    wire N__5445;
    wire N__5444;
    wire N__5441;
    wire N__5436;
    wire N__5431;
    wire N__5430;
    wire N__5427;
    wire N__5426;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5416;
    wire N__5413;
    wire N__5404;
    wire N__5403;
    wire N__5400;
    wire N__5397;
    wire N__5394;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5373;
    wire N__5372;
    wire N__5371;
    wire N__5370;
    wire N__5367;
    wire N__5360;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5338;
    wire N__5337;
    wire N__5336;
    wire N__5335;
    wire N__5334;
    wire N__5333;
    wire N__5332;
    wire N__5331;
    wire N__5330;
    wire N__5329;
    wire N__5326;
    wire N__5321;
    wire N__5316;
    wire N__5315;
    wire N__5314;
    wire N__5311;
    wire N__5310;
    wire N__5309;
    wire N__5308;
    wire N__5305;
    wire N__5304;
    wire N__5303;
    wire N__5300;
    wire N__5295;
    wire N__5292;
    wire N__5287;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5271;
    wire N__5268;
    wire N__5261;
    wire N__5258;
    wire N__5251;
    wire N__5236;
    wire N__5235;
    wire N__5234;
    wire N__5233;
    wire N__5230;
    wire N__5229;
    wire N__5228;
    wire N__5227;
    wire N__5224;
    wire N__5217;
    wire N__5214;
    wire N__5213;
    wire N__5212;
    wire N__5211;
    wire N__5210;
    wire N__5209;
    wire N__5208;
    wire N__5207;
    wire N__5204;
    wire N__5203;
    wire N__5200;
    wire N__5193;
    wire N__5190;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5182;
    wire N__5181;
    wire N__5176;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5164;
    wire N__5161;
    wire N__5156;
    wire N__5153;
    wire N__5148;
    wire N__5145;
    wire N__5142;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5113;
    wire N__5106;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5077;
    wire N__5076;
    wire N__5075;
    wire N__5074;
    wire N__5069;
    wire N__5068;
    wire N__5067;
    wire N__5066;
    wire N__5063;
    wire N__5062;
    wire N__5061;
    wire N__5060;
    wire N__5059;
    wire N__5058;
    wire N__5057;
    wire N__5056;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5040;
    wire N__5039;
    wire N__5036;
    wire N__5031;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4994;
    wire N__4991;
    wire N__4978;
    wire N__4977;
    wire N__4976;
    wire N__4975;
    wire N__4974;
    wire N__4973;
    wire N__4972;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4964;
    wire N__4963;
    wire N__4962;
    wire N__4961;
    wire N__4958;
    wire N__4953;
    wire N__4952;
    wire N__4947;
    wire N__4946;
    wire N__4945;
    wire N__4944;
    wire N__4941;
    wire N__4936;
    wire N__4929;
    wire N__4926;
    wire N__4925;
    wire N__4924;
    wire N__4919;
    wire N__4918;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4904;
    wire N__4897;
    wire N__4890;
    wire N__4887;
    wire N__4882;
    wire N__4867;
    wire N__4866;
    wire N__4865;
    wire N__4864;
    wire N__4861;
    wire N__4858;
    wire N__4857;
    wire N__4856;
    wire N__4853;
    wire N__4852;
    wire N__4849;
    wire N__4848;
    wire N__4847;
    wire N__4846;
    wire N__4845;
    wire N__4842;
    wire N__4839;
    wire N__4838;
    wire N__4837;
    wire N__4834;
    wire N__4833;
    wire N__4828;
    wire N__4825;
    wire N__4822;
    wire N__4819;
    wire N__4814;
    wire N__4811;
    wire N__4810;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4798;
    wire N__4793;
    wire N__4792;
    wire N__4791;
    wire N__4790;
    wire N__4785;
    wire N__4778;
    wire N__4775;
    wire N__4774;
    wire N__4771;
    wire N__4770;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4750;
    wire N__4743;
    wire N__4736;
    wire N__4733;
    wire N__4720;
    wire N__4719;
    wire N__4718;
    wire N__4717;
    wire N__4716;
    wire N__4715;
    wire N__4714;
    wire N__4713;
    wire N__4712;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4694;
    wire N__4693;
    wire N__4692;
    wire N__4691;
    wire N__4688;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4674;
    wire N__4673;
    wire N__4672;
    wire N__4665;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4647;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4639;
    wire N__4638;
    wire N__4637;
    wire N__4632;
    wire N__4627;
    wire N__4618;
    wire N__4613;
    wire N__4608;
    wire N__4603;
    wire N__4600;
    wire N__4585;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4573;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4558;
    wire N__4555;
    wire N__4554;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4546;
    wire N__4543;
    wire N__4536;
    wire N__4533;
    wire N__4530;
    wire N__4525;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4491;
    wire N__4490;
    wire N__4489;
    wire N__4488;
    wire N__4485;
    wire N__4484;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4474;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4453;
    wire N__4450;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4420;
    wire N__4417;
    wire N__4414;
    wire N__4411;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4399;
    wire N__4396;
    wire N__4393;
    wire N__4390;
    wire N__4387;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4375;
    wire N__4372;
    wire N__4371;
    wire N__4368;
    wire N__4367;
    wire N__4366;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4354;
    wire N__4351;
    wire N__4342;
    wire N__4339;
    wire N__4338;
    wire N__4337;
    wire N__4332;
    wire N__4331;
    wire N__4330;
    wire N__4329;
    wire N__4328;
    wire N__4327;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4315;
    wire N__4312;
    wire N__4307;
    wire N__4304;
    wire N__4291;
    wire N__4288;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4276;
    wire N__4273;
    wire N__4270;
    wire N__4267;
    wire N__4264;
    wire N__4261;
    wire N__4258;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4222;
    wire N__4219;
    wire N__4216;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4189;
    wire N__4186;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4174;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4161;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4144;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4134;
    wire N__4133;
    wire N__4130;
    wire N__4129;
    wire N__4128;
    wire N__4127;
    wire N__4122;
    wire N__4119;
    wire N__4116;
    wire N__4111;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4093;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4075;
    wire N__4074;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4057;
    wire N__4056;
    wire N__4055;
    wire N__4054;
    wire N__4053;
    wire N__4052;
    wire N__4051;
    wire N__4050;
    wire N__4049;
    wire N__4048;
    wire N__4047;
    wire N__4046;
    wire N__4045;
    wire N__4044;
    wire N__4043;
    wire N__4042;
    wire N__4041;
    wire N__4040;
    wire N__4039;
    wire N__4038;
    wire N__4037;
    wire N__4036;
    wire N__4035;
    wire N__4034;
    wire N__4033;
    wire N__4032;
    wire N__4031;
    wire N__4030;
    wire N__4029;
    wire N__4028;
    wire N__4027;
    wire N__4026;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3947;
    wire N__3944;
    wire N__3943;
    wire N__3942;
    wire N__3939;
    wire N__3938;
    wire N__3937;
    wire N__3934;
    wire N__3931;
    wire N__3926;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3904;
    wire N__3903;
    wire N__3900;
    wire N__3897;
    wire N__3896;
    wire N__3895;
    wire N__3892;
    wire N__3889;
    wire N__3886;
    wire N__3883;
    wire N__3874;
    wire N__3871;
    wire N__3868;
    wire N__3865;
    wire N__3864;
    wire N__3861;
    wire N__3858;
    wire N__3855;
    wire N__3852;
    wire N__3847;
    wire N__3844;
    wire N__3841;
    wire N__3838;
    wire N__3835;
    wire N__3832;
    wire N__3831;
    wire N__3828;
    wire N__3825;
    wire N__3820;
    wire N__3817;
    wire N__3816;
    wire N__3813;
    wire N__3810;
    wire N__3805;
    wire N__3802;
    wire N__3801;
    wire N__3798;
    wire N__3795;
    wire N__3790;
    wire N__3787;
    wire N__3784;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3772;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3760;
    wire N__3757;
    wire N__3754;
    wire N__3751;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3736;
    wire N__3733;
    wire N__3730;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3715;
    wire N__3712;
    wire N__3709;
    wire N__3706;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3696;
    wire N__3693;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3679;
    wire N__3676;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3664;
    wire N__3661;
    wire N__3658;
    wire N__3657;
    wire N__3652;
    wire N__3649;
    wire N__3648;
    wire N__3645;
    wire N__3642;
    wire N__3637;
    wire N__3634;
    wire N__3633;
    wire N__3632;
    wire N__3629;
    wire N__3624;
    wire N__3621;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3607;
    wire N__3606;
    wire N__3603;
    wire N__3600;
    wire N__3595;
    wire N__3592;
    wire N__3591;
    wire N__3588;
    wire N__3585;
    wire N__3580;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3568;
    wire N__3567;
    wire N__3562;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3550;
    wire N__3547;
    wire N__3544;
    wire N__3541;
    wire N__3540;
    wire N__3535;
    wire N__3532;
    wire N__3531;
    wire N__3530;
    wire N__3529;
    wire N__3528;
    wire N__3527;
    wire N__3526;
    wire N__3523;
    wire N__3520;
    wire N__3517;
    wire N__3508;
    wire N__3499;
    wire N__3498;
    wire N__3497;
    wire N__3494;
    wire N__3491;
    wire N__3488;
    wire N__3481;
    wire N__3480;
    wire N__3479;
    wire N__3476;
    wire N__3471;
    wire N__3466;
    wire N__3465;
    wire N__3464;
    wire N__3461;
    wire N__3458;
    wire N__3455;
    wire N__3452;
    wire N__3445;
    wire N__3444;
    wire N__3443;
    wire N__3440;
    wire N__3435;
    wire N__3430;
    wire N__3427;
    wire N__3424;
    wire N__3421;
    wire N__3418;
    wire N__3415;
    wire N__3412;
    wire N__3409;
    wire N__3406;
    wire N__3403;
    wire N__3400;
    wire N__3397;
    wire N__3394;
    wire N__3391;
    wire N__3388;
    wire N__3385;
    wire N__3382;
    wire N__3379;
    wire N__3376;
    wire N__3373;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3361;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3337;
    wire N__3334;
    wire N__3331;
    wire N__3330;
    wire N__3325;
    wire N__3322;
    wire N__3319;
    wire N__3316;
    wire N__3315;
    wire N__3312;
    wire N__3309;
    wire N__3308;
    wire N__3303;
    wire N__3300;
    wire N__3295;
    wire N__3292;
    wire N__3289;
    wire N__3288;
    wire N__3283;
    wire N__3280;
    wire N__3277;
    wire N__3276;
    wire N__3273;
    wire N__3270;
    wire N__3267;
    wire N__3262;
    wire N__3259;
    wire N__3256;
    wire N__3253;
    wire N__3250;
    wire N__3247;
    wire N__3244;
    wire N__3241;
    wire N__3238;
    wire N__3235;
    wire N__3232;
    wire N__3229;
    wire N__3226;
    wire N__3225;
    wire N__3222;
    wire N__3219;
    wire N__3216;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3190;
    wire N__3187;
    wire N__3186;
    wire N__3183;
    wire N__3180;
    wire N__3175;
    wire N__3172;
    wire N__3169;
    wire N__3166;
    wire N__3163;
    wire N__3160;
    wire N__3159;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3121;
    wire N__3118;
    wire N__3115;
    wire N__3112;
    wire N__3111;
    wire N__3110;
    wire N__3107;
    wire N__3102;
    wire N__3097;
    wire N__3096;
    wire N__3095;
    wire N__3094;
    wire N__3093;
    wire N__3088;
    wire N__3087;
    wire N__3084;
    wire N__3081;
    wire N__3078;
    wire N__3075;
    wire N__3072;
    wire N__3061;
    wire N__3058;
    wire N__3055;
    wire N__3052;
    wire N__3049;
    wire N__3046;
    wire N__3043;
    wire N__3040;
    wire N__3039;
    wire N__3036;
    wire N__3033;
    wire N__3028;
    wire N__3025;
    wire N__3022;
    wire N__3019;
    wire N__3016;
    wire N__3013;
    wire N__3010;
    wire N__3007;
    wire N__3006;
    wire N__3003;
    wire N__3000;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2980;
    wire N__2977;
    wire N__2974;
    wire N__2973;
    wire N__2972;
    wire N__2971;
    wire N__2970;
    wire N__2969;
    wire N__2966;
    wire N__2963;
    wire N__2960;
    wire N__2953;
    wire N__2944;
    wire N__2943;
    wire N__2942;
    wire N__2941;
    wire N__2940;
    wire N__2939;
    wire N__2938;
    wire N__2937;
    wire N__2932;
    wire N__2929;
    wire N__2918;
    wire N__2911;
    wire N__2910;
    wire N__2909;
    wire N__2908;
    wire N__2905;
    wire N__2904;
    wire N__2901;
    wire N__2898;
    wire N__2895;
    wire N__2892;
    wire N__2889;
    wire N__2886;
    wire N__2881;
    wire N__2878;
    wire N__2869;
    wire N__2868;
    wire N__2865;
    wire N__2862;
    wire N__2857;
    wire N__2856;
    wire N__2853;
    wire N__2850;
    wire N__2849;
    wire N__2848;
    wire N__2845;
    wire N__2842;
    wire N__2839;
    wire N__2836;
    wire N__2827;
    wire N__2826;
    wire N__2823;
    wire N__2820;
    wire N__2815;
    wire N__2812;
    wire N__2809;
    wire N__2806;
    wire N__2803;
    wire N__2800;
    wire N__2797;
    wire N__2796;
    wire N__2791;
    wire N__2788;
    wire N__2785;
    wire N__2782;
    wire N__2779;
    wire N__2776;
    wire N__2773;
    wire N__2770;
    wire N__2767;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2755;
    wire N__2752;
    wire N__2749;
    wire N__2746;
    wire N__2743;
    wire N__2740;
    wire N__2737;
    wire N__2734;
    wire N__2731;
    wire N__2728;
    wire N__2725;
    wire N__2722;
    wire N__2719;
    wire N__2716;
    wire N__2713;
    wire N__2710;
    wire N__2707;
    wire CLK40_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0 ;
    wire \U400_SDRAM.CO1 ;
    wire \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_ ;
    wire \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0 ;
    wire RESETn_c_i;
    wire CONSTANT_ONE_NET;
    wire A_c_31;
    wire A_c_30;
    wire A_c_27;
    wire \U400_SDRAM.un1_TA_COUNTER26_0_cascade_ ;
    wire \U400_SDRAM.TA_COUNTER23_cascade_ ;
    wire \U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_ ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_1 ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_0 ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_3 ;
    wire \U400_SDRAM.TA_COUNTER_0_sqmuxa ;
    wire \U400_SDRAM.TA_COUNTER23 ;
    wire \U400_SDRAM.TA_COUNTER27 ;
    wire \U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_ ;
    wire \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en ;
    wire \U400_SDRAM.BURSTZ0 ;
    wire \INVU400_SDRAM.BURSTC_net ;
    wire \U400_SDRAM.TACKZ0 ;
    wire \INVU400_SDRAM.TACKC_net ;
    wire A_c_22;
    wire BANK1_c;
    wire A_c_21;
    wire BANK0_c;
    wire \INVU400_SDRAM.BANK1C_net ;
    wire RASn_c;
    wire \INVU400_SDRAM.RASnC_net ;
    wire \U400_SDRAM.N_299_cascade_ ;
    wire \INVU400_SDRAM.SDRAM_CMD_2C_net ;
    wire \U400_SDRAM.N_52 ;
    wire \U400_SDRAM.N_295_0_cascade_ ;
    wire \U400_SDRAM.N_300_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_76_i_0 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_2_0_cascade_ ;
    wire \INVU400_SDRAM.SDRAM_CMD_0C_net ;
    wire \U400_SDRAM.N_110_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_a4_1_0_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_3_0_cascade_ ;
    wire \U400_SDRAM.N_55_cascade_ ;
    wire \U400_SDRAM.N_105_cascade_ ;
    wire \U400_SDRAM.N_68 ;
    wire \U400_SDRAM.N_62_cascade_ ;
    wire \U400_SDRAM.N_39_cascade_ ;
    wire \U400_SDRAM.N_62 ;
    wire A_c_23;
    wire \U400_SDRAM.N_41_cascade_ ;
    wire \INVU400_SDRAM.CS0_ENC_net ;
    wire \U400_SDRAM.N_57_cascade_ ;
    wire \U400_SDRAM.N_46 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_o5_0_cascade_ ;
    wire \U400_SDRAM.N_266_0_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD12 ;
    wire \U400_SDRAM.SDRAM_CMD12_cascade_ ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER52_0 ;
    wire \U400_SDRAM.CS0_ENZ0 ;
    wire CS0n_c;
    wire WEn_c;
    wire CASn_c;
    wire \INVU400_SDRAM.CS0nC_net ;
    wire \U400_SDRAM.CS1_ENZ0 ;
    wire CS1n_c;
    wire \INVU400_SDRAM.CS1nC_net ;
    wire A_c_9;
    wire A_c_17;
    wire MA_c_7;
    wire \INVU400_SDRAM.MA_nesr_7C_net ;
    wire A_c_8;
    wire A_c_16;
    wire MA_c_6;
    wire \INVU400_SDRAM.MA_nesr_6C_net ;
    wire bfn_5_4_0_;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_0 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_1 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_2 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_3 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_4 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_5 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_6 ;
    wire \INVU400_SDRAM.SDRAM_COUNTER_2C_net ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_76_i_a4_1_1 ;
    wire \U400_SDRAM.N_111 ;
    wire TSn_c;
    wire \U400_SDRAM.un3_RAM_CYCLE_START_cascade_ ;
    wire \U400_SDRAM.RAM_CYCLE_STARTZ0 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U400_SDRAM.N_54_cascade_ ;
    wire \U400_SDRAM.N_57 ;
    wire \U400_SDRAM.N_51 ;
    wire \INVU400_SDRAM.REFRESH_COUNTER_0C_net ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_0 ;
    wire bfn_5_7_0_;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_1 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_2 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_3 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_4 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_5 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_6 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_7 ;
    wire \INVU400_SDRAM.REFRESH_COUNTER_2C_net ;
    wire \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1 ;
    wire A_c_24;
    wire A_c_18;
    wire MA_c_8;
    wire \INVU400_SDRAM.MA_nesr_8C_net ;
    wire A_c_19;
    wire MA_c_9;
    wire \INVU400_SDRAM.MA_nesr_9C_net ;
    wire \U400_SDRAM.N_110 ;
    wire RnW_c;
    wire \INVU400_SDRAM.WRITE_CYCLEC_net ;
    wire \U400_SDRAM.TA_COUNTERZ0Z_2 ;
    wire \U400_SDRAM.TA_EN11_m ;
    wire \U400_SDRAM.un1_TA_COUNTER26_2_0 ;
    wire TA_OUT;
    wire CLK40_c_g;
    wire \U400_SDRAM.N_105 ;
    wire \U400_SDRAM.N_59 ;
    wire \U400_SDRAM.SDRAM_CMD_5_sqmuxa_cascade_ ;
    wire \U400_SDRAM.N_84 ;
    wire \U400_SDRAM.RAM_CYCLEZ0 ;
    wire \INVU400_SDRAM.RAM_CYCLEC_net ;
    wire \U400_SDRAM.N_30_2_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_1_0_cascade_ ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_3_0 ;
    wire \U400_SDRAM.N_30_2 ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER52_2_i_1 ;
    wire \U400_SDRAM.SDRAM_COUNTER44_5_cascade_ ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER44_0_cascade_ ;
    wire \U400_SDRAM.N_117 ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_1_cascade_ ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_4 ;
    wire \U400_SDRAM.SDRAM_COUNTER42 ;
    wire \U400_SDRAM.un1_SDRAM_COUNTER44_0 ;
    wire \U400_SDRAM.TACK_4_m ;
    wire \U400_SDRAM.TACK_7_0 ;
    wire \U400_SDRAM.N_56 ;
    wire \U400_SDRAM.N_56_cascade_ ;
    wire \U400_SDRAM.N_108 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_o2_0_0_cascade_ ;
    wire \U400_SDRAM.N_94_1 ;
    wire \U400_SDRAM.N_275_cascade_ ;
    wire \U400_SDRAM.N_54 ;
    wire \U400_SDRAM.N_276 ;
    wire A_c_26;
    wire MA_c_12;
    wire \INVU400_SDRAM.MA_nesr_12C_net ;
    wire A_c_20;
    wire MA_c_10;
    wire \INVU400_SDRAM.MA_nesr_10C_net ;
    wire \U400_BYTE_ENABLE.un2_LLBEn_0_0_cascade_ ;
    wire U400_BYTE_ENABLE_un1_LLBEn_i;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_76_i_a4_0 ;
    wire \U400_SDRAM.N_321_0_cascade_ ;
    wire \U400_SDRAM.N_322_0 ;
    wire \U400_SDRAM.WRITE_CYCLEZ0 ;
    wire \U400_SDRAM.N_320_0 ;
    wire \U400_SDRAM.SDRAM_COUNTER_s_0 ;
    wire \U400_SDRAM.N_88 ;
    wire \U400_SDRAM.SDRAM_COUNTER_s_3 ;
    wire \U400_SDRAM.N_303_0_i ;
    wire \U400_SDRAM.SDRAM_CMD_5_sqmuxa ;
    wire \U400_SDRAM.SDRAM_COUNTER_s_1 ;
    wire \INVU400_SDRAM.SDRAM_COUNTER_0C_net ;
    wire \U400_SDRAM.SDRAM_COUNTERe_0_i ;
    wire \INVU400_SDRAM.SDRAM_CONFIGUREDC_net ;
    wire \U400_SDRAM.N_66 ;
    wire \U400_SDRAM.N_55 ;
    wire \U400_SDRAM.SDRAM_CMD_3_sqmuxa ;
    wire \U400_SDRAM.SDRAM_CMD_3_sqmuxa_cascade_ ;
    wire \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_1_0 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_0 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_8 ;
    wire \U400_SDRAM.SDRAM_CONFIGUREDZ0 ;
    wire RESETn_c;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_a5_0_0 ;
    wire \U400_SDRAM.N_299_2 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_0_tz_cascade_ ;
    wire \U400_SDRAM.N_266_0 ;
    wire \U400_SDRAM.N_270 ;
    wire \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_0_0_cascade_ ;
    wire \U400_SDRAM.N_43 ;
    wire \INVU400_SDRAM.SDRAM_CMD_1C_net ;
    wire A_c_25;
    wire MA_c_11;
    wire \INVU400_SDRAM.MA_nesr_11C_net ;
    wire U400_BYTE_ENABLE_un1_UMBEn_i;
    wire U400_BYTE_ENABLE_un1_LMBEn_i;
    wire RAM_SPACEm;
    wire U400_BYTE_ENABLE_un1_UUBEn_i;
    wire A_c_0;
    wire A_c_1;
    wire \U400_BYTE_ENABLE.un2_UMBEn_0_0 ;
    wire \U400_BYTE_ENABLE.LW_TRANS_0 ;
    wire U400_ADDRESS_DECODE_RAM_SPACE_3;
    wire A_c_29;
    wire A_c_28;
    wire RAM_SPACEm_i;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire \U400_SDRAM.BURSTZ0Z8 ;
    wire A_c_7;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_1 ;
    wire A_c_3;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_0 ;
    wire A_c_15;
    wire \U400_SDRAM.MA_5_iv_0_5 ;
    wire MA_c_5;
    wire \INVU400_SDRAM.MA_nesr_5C_net ;
    wire A_c_5;
    wire A_c_13;
    wire MA_c_3;
    wire \INVU400_SDRAM.MA_nesr_3C_net ;
    wire A_c_6;
    wire A_c_14;
    wire MA_c_4;
    wire A_c_2;
    wire A_c_10;
    wire MA_c_0;
    wire A_c_11;
    wire \U400_SDRAM.MA_5_iv_0_1 ;
    wire MA_c_1;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_2 ;
    wire A_c_4;
    wire A_c_12;
    wire \U400_SDRAM.MA19 ;
    wire MA_c_2;
    wire \INVU400_SDRAM.MA_nesr_4C_net ;
    wire \U400_SDRAM.un1_MA20_0_i_0 ;
    wire RESETn_c_i_g;
    wire TA_EN_i_ess;
    wire N_474_i;
    wire _gnd_net_;

    IO_PAD MA_obuf_7_iopad (
            .OE(N__7451),
            .DIN(N__7450),
            .DOUT(N__7449),
            .PACKAGEPIN(MA[7]));
    defparam MA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_7_preio (
            .PADOEN(N__7451),
            .PADOUT(N__7450),
            .PADIN(N__7449),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3400),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__7442),
            .DIN(N__7441),
            .DOUT(N__7440),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__7442),
            .PADOUT(N__7441),
            .PADIN(N__7440),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__7433),
            .DIN(N__7432),
            .DOUT(N__7431),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__7433),
            .PADOUT(N__7432),
            .PADIN(N__7431),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3238),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__7424),
            .DIN(N__7423),
            .DOUT(N__7422),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__7424),
            .PADOUT(N__7423),
            .PADIN(N__7422),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3049),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_8_iopad (
            .OE(N__7415),
            .DIN(N__7414),
            .DOUT(N__7413),
            .PACKAGEPIN(MA[8]));
    defparam MA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_8_preio (
            .PADOEN(N__7415),
            .PADOUT(N__7414),
            .PADIN(N__7413),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3736),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_10_iopad (
            .OE(N__7406),
            .DIN(N__7405),
            .DOUT(N__7404),
            .PACKAGEPIN(MA[10]));
    defparam MA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_10_preio (
            .PADOEN(N__7406),
            .PADOUT(N__7405),
            .PADIN(N__7404),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4243),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__7397),
            .DIN(N__7396),
            .DOUT(N__7395),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__7397),
            .PADOUT(N__7396),
            .PADIN(N__7395),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_2_iopad (
            .OE(N__7388),
            .DIN(N__7387),
            .DOUT(N__7386),
            .PACKAGEPIN(MA[2]));
    defparam MA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_2_preio (
            .PADOEN(N__7388),
            .PADOUT(N__7387),
            .PADIN(N__7386),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6607),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__7379),
            .DIN(N__7378),
            .DOUT(N__7377),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__7379),
            .PADOUT(N__7378),
            .PADIN(N__7377),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__7370),
            .DIN(N__7369),
            .DOUT(N__7368),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__7370),
            .PADOUT(N__7369),
            .PADIN(N__7368),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__7361),
            .DIN(N__7360),
            .DOUT(N__7359),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__7361),
            .PADOUT(N__7360),
            .PADIN(N__7359),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5824),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__7352),
            .DIN(N__7351),
            .DOUT(N__7350),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__7352),
            .PADOUT(N__7351),
            .PADIN(N__7350),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__7343),
            .DIN(N__7342),
            .DOUT(N__7341),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__7343),
            .PADOUT(N__7342),
            .PADIN(N__7341),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__7334),
            .DIN(N__7333),
            .DOUT(N__7332),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__7334),
            .PADOUT(N__7333),
            .PADIN(N__7332),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_12_iopad (
            .OE(N__7325),
            .DIN(N__7324),
            .DOUT(N__7323),
            .PACKAGEPIN(MA[12]));
    defparam MA_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_12_preio (
            .PADOEN(N__7325),
            .PADOUT(N__7324),
            .PADIN(N__7323),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4267),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_1_iopad (
            .OE(N__7316),
            .DIN(N__7315),
            .DOUT(N__7314),
            .PACKAGEPIN(MA[1]));
    defparam MA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_1_preio (
            .PADOEN(N__7316),
            .PADOUT(N__7315),
            .PADIN(N__7314),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6856),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__7307),
            .DIN(N__7306),
            .DOUT(N__7305),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__7307),
            .PADOUT(N__7306),
            .PADIN(N__7305),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__7298),
            .DIN(N__7297),
            .DOUT(N__7296),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__7298),
            .PADOUT(N__7297),
            .PADIN(N__7296),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__7289),
            .DIN(N__7288),
            .DOUT(N__7287),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__7289),
            .PADOUT(N__7288),
            .PADIN(N__7287),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_4_iopad (
            .OE(N__7280),
            .DIN(N__7279),
            .DOUT(N__7278),
            .PACKAGEPIN(MA[4]));
    defparam MA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_4_preio (
            .PADOEN(N__7280),
            .PADOUT(N__7279),
            .PADIN(N__7278),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5992),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__7271),
            .DIN(N__7270),
            .DOUT(N__7269),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__7271),
            .PADOUT(N__7270),
            .PADIN(N__7269),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__7262),
            .DIN(N__7261),
            .DOUT(N__7260),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__7262),
            .PADOUT(N__7261),
            .PADIN(N__7260),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__7253),
            .DIN(N__7252),
            .DOUT(N__7251),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__7253),
            .PADOUT(N__7252),
            .PADIN(N__7251),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4522),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__7244),
            .DIN(N__7243),
            .DOUT(N__7242),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__7244),
            .PADOUT(N__7243),
            .PADIN(N__7242),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_9_iopad (
            .OE(N__7235),
            .DIN(N__7234),
            .DOUT(N__7233),
            .PACKAGEPIN(MA[9]));
    defparam MA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_9_preio (
            .PADOEN(N__7235),
            .PADOUT(N__7234),
            .PADIN(N__7233),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3709),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__7226),
            .DIN(N__7225),
            .DOUT(N__7224),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__7226),
            .PADOUT(N__7225),
            .PADIN(N__7224),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5863),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__7217),
            .DIN(N__7216),
            .DOUT(N__7215),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__7217),
            .PADOUT(N__7216),
            .PADIN(N__7215),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__7208),
            .DIN(N__7207),
            .DOUT(N__7206),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__7208),
            .PADOUT(N__7207),
            .PADIN(N__7206),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__7199),
            .DIN(N__7198),
            .DOUT(N__7197),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__7199),
            .PADOUT(N__7198),
            .PADIN(N__7197),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2767),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__7190),
            .DIN(N__7189),
            .DOUT(N__7188),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__7190),
            .PADOUT(N__7189),
            .PADIN(N__7188),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__7181),
            .DIN(N__7180),
            .DOUT(N__7179),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__7181),
            .PADOUT(N__7180),
            .PADIN(N__7179),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_3_iopad (
            .OE(N__7172),
            .DIN(N__7171),
            .DOUT(N__7170),
            .PACKAGEPIN(MA[3]));
    defparam MA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_3_preio (
            .PADOEN(N__7172),
            .PADOUT(N__7171),
            .PADIN(N__7170),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6037),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__7163),
            .DIN(N__7162),
            .DOUT(N__7161),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__7163),
            .PADOUT(N__7162),
            .PADIN(N__7161),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__7154),
            .DIN(N__7153),
            .DOUT(N__7152),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__7154),
            .PADOUT(N__7153),
            .PADIN(N__7152),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__7145),
            .DIN(N__7144),
            .DOUT(N__7143),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__7145),
            .PADOUT(N__7144),
            .PADIN(N__7143),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_6_iopad (
            .OE(N__7136),
            .DIN(N__7135),
            .DOUT(N__7134),
            .PACKAGEPIN(MA[6]));
    defparam MA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_6_preio (
            .PADOEN(N__7136),
            .PADOUT(N__7135),
            .PADIN(N__7134),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3364),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__7127),
            .DIN(N__7126),
            .DOUT(N__7125),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__7127),
            .PADOUT(N__7126),
            .PADIN(N__7125),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__7118),
            .DIN(N__7117),
            .DOUT(N__7116),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__7118),
            .PADOUT(N__7117),
            .PADIN(N__7116),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__7109),
            .DIN(N__7108),
            .DOUT(N__7107),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__7109),
            .PADOUT(N__7108),
            .PADIN(N__7107),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__7100),
            .DIN(N__7099),
            .DOUT(N__7098),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__7100),
            .PADOUT(N__7099),
            .PADIN(N__7098),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2995),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__7091),
            .DIN(N__7090),
            .DOUT(N__7089),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__7091),
            .PADOUT(N__7090),
            .PADIN(N__7089),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__7082),
            .DIN(N__7081),
            .DOUT(N__7080),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__7082),
            .PADOUT(N__7081),
            .PADIN(N__7080),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3013),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_11_iopad (
            .OE(N__7073),
            .DIN(N__7072),
            .DOUT(N__7071),
            .PACKAGEPIN(MA[11]));
    defparam MA_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_11_preio (
            .PADOEN(N__7073),
            .PADOUT(N__7072),
            .PADIN(N__7071),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5872),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TAn_obuft_iopad (
            .OE(N__7064),
            .DIN(N__7063),
            .DOUT(N__7062),
            .PACKAGEPIN(TAn));
    defparam TAn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TAn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TAn_obuft_preio (
            .PADOEN(N__7064),
            .PADOUT(N__7063),
            .PADIN(N__7062),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6412),
            .DIN0(),
            .DOUT0(N__4084),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__7055),
            .DIN(N__7054),
            .DOUT(N__7053),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__7055),
            .PADOUT(N__7054),
            .PADIN(N__7053),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_5_iopad (
            .OE(N__7046),
            .DIN(N__7045),
            .DOUT(N__7044),
            .PACKAGEPIN(MA[5]));
    defparam MA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_5_preio (
            .PADOEN(N__7046),
            .PADOUT(N__7045),
            .PADIN(N__7044),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6076),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__7037),
            .DIN(N__7036),
            .DOUT(N__7035),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__7037),
            .PADOUT(N__7036),
            .PADIN(N__7035),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__7028),
            .DIN(N__7027),
            .DOUT(N__7026),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__7028),
            .PADOUT(N__7027),
            .PADIN(N__7026),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LBENn_obuf_iopad.PULLUP=1'b1;
    IO_PAD LBENn_obuf_iopad (
            .OE(N__7019),
            .DIN(N__7018),
            .DOUT(N__7017),
            .PACKAGEPIN(LBENn));
    defparam LBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LBENn_obuf_preio (
            .PADOEN(N__7019),
            .PADOUT(N__7018),
            .PADIN(N__7017),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5599),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__7010),
            .DIN(N__7009),
            .DOUT(N__7008),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__7010),
            .PADOUT(N__7009),
            .PADIN(N__7008),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CS1n_obuf_iopad (
            .OE(N__7001),
            .DIN(N__7000),
            .DOUT(N__6999),
            .PACKAGEPIN(CS1n));
    defparam CS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CS1n_obuf_preio (
            .PADOEN(N__7001),
            .PADOUT(N__7000),
            .PADIN(N__6999),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3211),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__6992),
            .DIN(N__6991),
            .DOUT(N__6990),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__6992),
            .PADOUT(N__6991),
            .PADIN(N__6990),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__6983),
            .DIN(N__6982),
            .DOUT(N__6981),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__6983),
            .PADOUT(N__6982),
            .PADIN(N__6981),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__6974),
            .DIN(N__6973),
            .DOUT(N__6972),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__6974),
            .PADOUT(N__6973),
            .PADIN(N__6972),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__6965),
            .DIN(N__6964),
            .DOUT(N__6963),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__6965),
            .PADOUT(N__6964),
            .PADIN(N__6963),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__6956),
            .DIN(N__6955),
            .DOUT(N__6954),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__6956),
            .PADOUT(N__6955),
            .PADIN(N__6954),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3247),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_0_iopad (
            .OE(N__6947),
            .DIN(N__6946),
            .DOUT(N__6945),
            .PACKAGEPIN(MA[0]));
    defparam MA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_0_preio (
            .PADOEN(N__6947),
            .PADOUT(N__6946),
            .PADIN(N__6945),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5950),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__6938),
            .DIN(N__6937),
            .DOUT(N__6936),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__6938),
            .PADOUT(N__6937),
            .PADIN(N__6936),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__6929),
            .DIN(N__6928),
            .DOUT(N__6927),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__6929),
            .PADOUT(N__6928),
            .PADIN(N__6927),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__6920),
            .DIN(N__6919),
            .DOUT(N__6918),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__6920),
            .PADOUT(N__6919),
            .PADIN(N__6918),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CS0n_obuf_iopad (
            .OE(N__6911),
            .DIN(N__6910),
            .DOUT(N__6909),
            .PACKAGEPIN(CS0n));
    defparam CS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CS0n_obuf_preio (
            .PADOEN(N__6911),
            .PADOUT(N__6910),
            .PADIN(N__6909),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3262),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__6902),
            .DIN(N__6901),
            .DOUT(N__6900),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__6902),
            .PADOUT(N__6901),
            .PADIN(N__6900),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__6893),
            .DIN(N__6892),
            .DOUT(N__6891),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__6893),
            .PADOUT(N__6892),
            .PADIN(N__6891),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5854),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__6884),
            .DIN(N__6883),
            .DOUT(N__6882),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__6884),
            .PADOUT(N__6883),
            .PADIN(N__6882),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_ibuf_gb_io_iopad (
            .OE(N__6875),
            .DIN(N__6874),
            .DOUT(N__6873),
            .PACKAGEPIN(CLK40));
    defparam CLK40_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_ibuf_gb_io_preio (
            .PADOEN(N__6875),
            .PADOUT(N__6874),
            .PADIN(N__6873),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__1634 (
            .O(N__6856),
            .I(N__6853));
    LocalMux I__1633 (
            .O(N__6853),
            .I(N__6850));
    Odrv4 I__1632 (
            .O(N__6850),
            .I(MA_c_1));
    InMux I__1631 (
            .O(N__6847),
            .I(N__6836));
    InMux I__1630 (
            .O(N__6846),
            .I(N__6827));
    InMux I__1629 (
            .O(N__6845),
            .I(N__6827));
    InMux I__1628 (
            .O(N__6844),
            .I(N__6827));
    InMux I__1627 (
            .O(N__6843),
            .I(N__6824));
    InMux I__1626 (
            .O(N__6842),
            .I(N__6818));
    InMux I__1625 (
            .O(N__6841),
            .I(N__6813));
    InMux I__1624 (
            .O(N__6840),
            .I(N__6813));
    InMux I__1623 (
            .O(N__6839),
            .I(N__6810));
    LocalMux I__1622 (
            .O(N__6836),
            .I(N__6807));
    InMux I__1621 (
            .O(N__6835),
            .I(N__6804));
    InMux I__1620 (
            .O(N__6834),
            .I(N__6801));
    LocalMux I__1619 (
            .O(N__6827),
            .I(N__6796));
    LocalMux I__1618 (
            .O(N__6824),
            .I(N__6796));
    InMux I__1617 (
            .O(N__6823),
            .I(N__6793));
    InMux I__1616 (
            .O(N__6822),
            .I(N__6790));
    InMux I__1615 (
            .O(N__6821),
            .I(N__6787));
    LocalMux I__1614 (
            .O(N__6818),
            .I(N__6780));
    LocalMux I__1613 (
            .O(N__6813),
            .I(N__6780));
    LocalMux I__1612 (
            .O(N__6810),
            .I(N__6780));
    Span4Mux_v I__1611 (
            .O(N__6807),
            .I(N__6777));
    LocalMux I__1610 (
            .O(N__6804),
            .I(N__6773));
    LocalMux I__1609 (
            .O(N__6801),
            .I(N__6767));
    Span4Mux_v I__1608 (
            .O(N__6796),
            .I(N__6764));
    LocalMux I__1607 (
            .O(N__6793),
            .I(N__6757));
    LocalMux I__1606 (
            .O(N__6790),
            .I(N__6757));
    LocalMux I__1605 (
            .O(N__6787),
            .I(N__6757));
    Span4Mux_v I__1604 (
            .O(N__6780),
            .I(N__6754));
    Sp12to4 I__1603 (
            .O(N__6777),
            .I(N__6750));
    InMux I__1602 (
            .O(N__6776),
            .I(N__6747));
    Span4Mux_s3_h I__1601 (
            .O(N__6773),
            .I(N__6744));
    InMux I__1600 (
            .O(N__6772),
            .I(N__6741));
    InMux I__1599 (
            .O(N__6771),
            .I(N__6738));
    InMux I__1598 (
            .O(N__6770),
            .I(N__6735));
    Span4Mux_h I__1597 (
            .O(N__6767),
            .I(N__6732));
    Span4Mux_h I__1596 (
            .O(N__6764),
            .I(N__6727));
    Span4Mux_v I__1595 (
            .O(N__6757),
            .I(N__6727));
    Span4Mux_h I__1594 (
            .O(N__6754),
            .I(N__6724));
    InMux I__1593 (
            .O(N__6753),
            .I(N__6721));
    Span12Mux_s8_h I__1592 (
            .O(N__6750),
            .I(N__6706));
    LocalMux I__1591 (
            .O(N__6747),
            .I(N__6706));
    Sp12to4 I__1590 (
            .O(N__6744),
            .I(N__6706));
    LocalMux I__1589 (
            .O(N__6741),
            .I(N__6706));
    LocalMux I__1588 (
            .O(N__6738),
            .I(N__6706));
    LocalMux I__1587 (
            .O(N__6735),
            .I(N__6706));
    Sp12to4 I__1586 (
            .O(N__6732),
            .I(N__6706));
    Span4Mux_v I__1585 (
            .O(N__6727),
            .I(N__6703));
    Span4Mux_v I__1584 (
            .O(N__6724),
            .I(N__6700));
    LocalMux I__1583 (
            .O(N__6721),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    Odrv12 I__1582 (
            .O(N__6706),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1581 (
            .O(N__6703),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1580 (
            .O(N__6700),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    InMux I__1579 (
            .O(N__6691),
            .I(N__6688));
    LocalMux I__1578 (
            .O(N__6688),
            .I(N__6685));
    Span4Mux_v I__1577 (
            .O(N__6685),
            .I(N__6682));
    Odrv4 I__1576 (
            .O(N__6682),
            .I(A_c_4));
    CascadeMux I__1575 (
            .O(N__6679),
            .I(N__6676));
    InMux I__1574 (
            .O(N__6676),
            .I(N__6673));
    LocalMux I__1573 (
            .O(N__6673),
            .I(N__6670));
    Odrv4 I__1572 (
            .O(N__6670),
            .I(A_c_12));
    InMux I__1571 (
            .O(N__6667),
            .I(N__6660));
    InMux I__1570 (
            .O(N__6666),
            .I(N__6649));
    InMux I__1569 (
            .O(N__6665),
            .I(N__6649));
    InMux I__1568 (
            .O(N__6664),
            .I(N__6649));
    InMux I__1567 (
            .O(N__6663),
            .I(N__6649));
    LocalMux I__1566 (
            .O(N__6660),
            .I(N__6645));
    InMux I__1565 (
            .O(N__6659),
            .I(N__6642));
    InMux I__1564 (
            .O(N__6658),
            .I(N__6639));
    LocalMux I__1563 (
            .O(N__6649),
            .I(N__6635));
    InMux I__1562 (
            .O(N__6648),
            .I(N__6632));
    Span12Mux_s4_v I__1561 (
            .O(N__6645),
            .I(N__6625));
    LocalMux I__1560 (
            .O(N__6642),
            .I(N__6625));
    LocalMux I__1559 (
            .O(N__6639),
            .I(N__6625));
    InMux I__1558 (
            .O(N__6638),
            .I(N__6622));
    Span4Mux_s2_v I__1557 (
            .O(N__6635),
            .I(N__6619));
    LocalMux I__1556 (
            .O(N__6632),
            .I(N__6616));
    Odrv12 I__1555 (
            .O(N__6625),
            .I(\U400_SDRAM.MA19 ));
    LocalMux I__1554 (
            .O(N__6622),
            .I(\U400_SDRAM.MA19 ));
    Odrv4 I__1553 (
            .O(N__6619),
            .I(\U400_SDRAM.MA19 ));
    Odrv12 I__1552 (
            .O(N__6616),
            .I(\U400_SDRAM.MA19 ));
    IoInMux I__1551 (
            .O(N__6607),
            .I(N__6604));
    LocalMux I__1550 (
            .O(N__6604),
            .I(N__6601));
    Odrv4 I__1549 (
            .O(N__6601),
            .I(MA_c_2));
    CEMux I__1548 (
            .O(N__6598),
            .I(N__6594));
    CEMux I__1547 (
            .O(N__6597),
            .I(N__6589));
    LocalMux I__1546 (
            .O(N__6594),
            .I(N__6585));
    CEMux I__1545 (
            .O(N__6593),
            .I(N__6582));
    CEMux I__1544 (
            .O(N__6592),
            .I(N__6576));
    LocalMux I__1543 (
            .O(N__6589),
            .I(N__6573));
    CEMux I__1542 (
            .O(N__6588),
            .I(N__6570));
    Span4Mux_s3_h I__1541 (
            .O(N__6585),
            .I(N__6564));
    LocalMux I__1540 (
            .O(N__6582),
            .I(N__6564));
    CEMux I__1539 (
            .O(N__6581),
            .I(N__6561));
    CEMux I__1538 (
            .O(N__6580),
            .I(N__6558));
    CEMux I__1537 (
            .O(N__6579),
            .I(N__6555));
    LocalMux I__1536 (
            .O(N__6576),
            .I(N__6547));
    Span4Mux_v I__1535 (
            .O(N__6573),
            .I(N__6547));
    LocalMux I__1534 (
            .O(N__6570),
            .I(N__6547));
    CEMux I__1533 (
            .O(N__6569),
            .I(N__6544));
    Span4Mux_h I__1532 (
            .O(N__6564),
            .I(N__6535));
    LocalMux I__1531 (
            .O(N__6561),
            .I(N__6535));
    LocalMux I__1530 (
            .O(N__6558),
            .I(N__6535));
    LocalMux I__1529 (
            .O(N__6555),
            .I(N__6535));
    CEMux I__1528 (
            .O(N__6554),
            .I(N__6532));
    Sp12to4 I__1527 (
            .O(N__6547),
            .I(N__6527));
    LocalMux I__1526 (
            .O(N__6544),
            .I(N__6527));
    Sp12to4 I__1525 (
            .O(N__6535),
            .I(N__6522));
    LocalMux I__1524 (
            .O(N__6532),
            .I(N__6522));
    Odrv12 I__1523 (
            .O(N__6527),
            .I(\U400_SDRAM.un1_MA20_0_i_0 ));
    Odrv12 I__1522 (
            .O(N__6522),
            .I(\U400_SDRAM.un1_MA20_0_i_0 ));
    CascadeMux I__1521 (
            .O(N__6517),
            .I(N__6514));
    InMux I__1520 (
            .O(N__6514),
            .I(N__6510));
    InMux I__1519 (
            .O(N__6513),
            .I(N__6507));
    LocalMux I__1518 (
            .O(N__6510),
            .I(N__6497));
    LocalMux I__1517 (
            .O(N__6507),
            .I(N__6483));
    SRMux I__1516 (
            .O(N__6506),
            .I(N__6430));
    SRMux I__1515 (
            .O(N__6505),
            .I(N__6430));
    SRMux I__1514 (
            .O(N__6504),
            .I(N__6430));
    SRMux I__1513 (
            .O(N__6503),
            .I(N__6430));
    SRMux I__1512 (
            .O(N__6502),
            .I(N__6430));
    SRMux I__1511 (
            .O(N__6501),
            .I(N__6430));
    SRMux I__1510 (
            .O(N__6500),
            .I(N__6430));
    Glb2LocalMux I__1509 (
            .O(N__6497),
            .I(N__6430));
    SRMux I__1508 (
            .O(N__6496),
            .I(N__6430));
    SRMux I__1507 (
            .O(N__6495),
            .I(N__6430));
    SRMux I__1506 (
            .O(N__6494),
            .I(N__6430));
    SRMux I__1505 (
            .O(N__6493),
            .I(N__6430));
    SRMux I__1504 (
            .O(N__6492),
            .I(N__6430));
    SRMux I__1503 (
            .O(N__6491),
            .I(N__6430));
    SRMux I__1502 (
            .O(N__6490),
            .I(N__6430));
    SRMux I__1501 (
            .O(N__6489),
            .I(N__6430));
    SRMux I__1500 (
            .O(N__6488),
            .I(N__6430));
    SRMux I__1499 (
            .O(N__6487),
            .I(N__6430));
    SRMux I__1498 (
            .O(N__6486),
            .I(N__6430));
    Glb2LocalMux I__1497 (
            .O(N__6483),
            .I(N__6430));
    SRMux I__1496 (
            .O(N__6482),
            .I(N__6430));
    SRMux I__1495 (
            .O(N__6481),
            .I(N__6430));
    SRMux I__1494 (
            .O(N__6480),
            .I(N__6430));
    SRMux I__1493 (
            .O(N__6479),
            .I(N__6430));
    GlobalMux I__1492 (
            .O(N__6430),
            .I(N__6427));
    gio2CtrlBuf I__1491 (
            .O(N__6427),
            .I(RESETn_c_i_g));
    InMux I__1490 (
            .O(N__6424),
            .I(N__6421));
    LocalMux I__1489 (
            .O(N__6421),
            .I(N__6418));
    Span12Mux_s6_h I__1488 (
            .O(N__6418),
            .I(N__6415));
    Odrv12 I__1487 (
            .O(N__6415),
            .I(TA_EN_i_ess));
    IoInMux I__1486 (
            .O(N__6412),
            .I(N__6409));
    LocalMux I__1485 (
            .O(N__6409),
            .I(N__6406));
    Odrv4 I__1484 (
            .O(N__6406),
            .I(N_474_i));
    InMux I__1483 (
            .O(N__6403),
            .I(N__6397));
    InMux I__1482 (
            .O(N__6402),
            .I(N__6394));
    InMux I__1481 (
            .O(N__6401),
            .I(N__6389));
    InMux I__1480 (
            .O(N__6400),
            .I(N__6389));
    LocalMux I__1479 (
            .O(N__6397),
            .I(N__6385));
    LocalMux I__1478 (
            .O(N__6394),
            .I(N__6382));
    LocalMux I__1477 (
            .O(N__6389),
            .I(N__6379));
    InMux I__1476 (
            .O(N__6388),
            .I(N__6376));
    Sp12to4 I__1475 (
            .O(N__6385),
            .I(N__6373));
    Span4Mux_h I__1474 (
            .O(N__6382),
            .I(N__6370));
    Span4Mux_h I__1473 (
            .O(N__6379),
            .I(N__6365));
    LocalMux I__1472 (
            .O(N__6376),
            .I(N__6365));
    Span12Mux_s7_v I__1471 (
            .O(N__6373),
            .I(N__6362));
    Span4Mux_v I__1470 (
            .O(N__6370),
            .I(N__6357));
    Span4Mux_v I__1469 (
            .O(N__6365),
            .I(N__6357));
    Odrv12 I__1468 (
            .O(N__6362),
            .I(SIZ_c_0));
    Odrv4 I__1467 (
            .O(N__6357),
            .I(SIZ_c_0));
    CascadeMux I__1466 (
            .O(N__6352),
            .I(N__6349));
    InMux I__1465 (
            .O(N__6349),
            .I(N__6344));
    CascadeMux I__1464 (
            .O(N__6348),
            .I(N__6341));
    CascadeMux I__1463 (
            .O(N__6347),
            .I(N__6338));
    LocalMux I__1462 (
            .O(N__6344),
            .I(N__6335));
    InMux I__1461 (
            .O(N__6341),
            .I(N__6332));
    InMux I__1460 (
            .O(N__6338),
            .I(N__6329));
    Odrv12 I__1459 (
            .O(N__6335),
            .I(\U400_SDRAM.BURSTZ0Z8 ));
    LocalMux I__1458 (
            .O(N__6332),
            .I(\U400_SDRAM.BURSTZ0Z8 ));
    LocalMux I__1457 (
            .O(N__6329),
            .I(\U400_SDRAM.BURSTZ0Z8 ));
    CascadeMux I__1456 (
            .O(N__6322),
            .I(N__6319));
    InMux I__1455 (
            .O(N__6319),
            .I(N__6316));
    LocalMux I__1454 (
            .O(N__6316),
            .I(N__6313));
    Odrv12 I__1453 (
            .O(N__6313),
            .I(A_c_7));
    CascadeMux I__1452 (
            .O(N__6310),
            .I(N__6302));
    InMux I__1451 (
            .O(N__6309),
            .I(N__6296));
    InMux I__1450 (
            .O(N__6308),
            .I(N__6296));
    InMux I__1449 (
            .O(N__6307),
            .I(N__6293));
    InMux I__1448 (
            .O(N__6306),
            .I(N__6289));
    InMux I__1447 (
            .O(N__6305),
            .I(N__6283));
    InMux I__1446 (
            .O(N__6302),
            .I(N__6280));
    InMux I__1445 (
            .O(N__6301),
            .I(N__6277));
    LocalMux I__1444 (
            .O(N__6296),
            .I(N__6274));
    LocalMux I__1443 (
            .O(N__6293),
            .I(N__6271));
    InMux I__1442 (
            .O(N__6292),
            .I(N__6268));
    LocalMux I__1441 (
            .O(N__6289),
            .I(N__6265));
    InMux I__1440 (
            .O(N__6288),
            .I(N__6262));
    InMux I__1439 (
            .O(N__6287),
            .I(N__6259));
    InMux I__1438 (
            .O(N__6286),
            .I(N__6256));
    LocalMux I__1437 (
            .O(N__6283),
            .I(N__6244));
    LocalMux I__1436 (
            .O(N__6280),
            .I(N__6244));
    LocalMux I__1435 (
            .O(N__6277),
            .I(N__6244));
    Span4Mux_h I__1434 (
            .O(N__6274),
            .I(N__6244));
    Span4Mux_h I__1433 (
            .O(N__6271),
            .I(N__6244));
    LocalMux I__1432 (
            .O(N__6268),
            .I(N__6241));
    Span4Mux_h I__1431 (
            .O(N__6265),
            .I(N__6232));
    LocalMux I__1430 (
            .O(N__6262),
            .I(N__6232));
    LocalMux I__1429 (
            .O(N__6259),
            .I(N__6232));
    LocalMux I__1428 (
            .O(N__6256),
            .I(N__6232));
    InMux I__1427 (
            .O(N__6255),
            .I(N__6229));
    Span4Mux_v I__1426 (
            .O(N__6244),
            .I(N__6226));
    Span4Mux_h I__1425 (
            .O(N__6241),
            .I(N__6221));
    Span4Mux_v I__1424 (
            .O(N__6232),
            .I(N__6221));
    LocalMux I__1423 (
            .O(N__6229),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1422 (
            .O(N__6226),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1421 (
            .O(N__6221),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    CascadeMux I__1420 (
            .O(N__6214),
            .I(N__6211));
    InMux I__1419 (
            .O(N__6211),
            .I(N__6208));
    LocalMux I__1418 (
            .O(N__6208),
            .I(N__6205));
    Span4Mux_h I__1417 (
            .O(N__6205),
            .I(N__6202));
    Odrv4 I__1416 (
            .O(N__6202),
            .I(A_c_3));
    InMux I__1415 (
            .O(N__6199),
            .I(N__6189));
    InMux I__1414 (
            .O(N__6198),
            .I(N__6189));
    InMux I__1413 (
            .O(N__6197),
            .I(N__6184));
    InMux I__1412 (
            .O(N__6196),
            .I(N__6181));
    InMux I__1411 (
            .O(N__6195),
            .I(N__6178));
    InMux I__1410 (
            .O(N__6194),
            .I(N__6175));
    LocalMux I__1409 (
            .O(N__6189),
            .I(N__6172));
    InMux I__1408 (
            .O(N__6188),
            .I(N__6167));
    CascadeMux I__1407 (
            .O(N__6187),
            .I(N__6164));
    LocalMux I__1406 (
            .O(N__6184),
            .I(N__6160));
    LocalMux I__1405 (
            .O(N__6181),
            .I(N__6157));
    LocalMux I__1404 (
            .O(N__6178),
            .I(N__6154));
    LocalMux I__1403 (
            .O(N__6175),
            .I(N__6149));
    Span4Mux_s3_v I__1402 (
            .O(N__6172),
            .I(N__6149));
    InMux I__1401 (
            .O(N__6171),
            .I(N__6146));
    InMux I__1400 (
            .O(N__6170),
            .I(N__6143));
    LocalMux I__1399 (
            .O(N__6167),
            .I(N__6140));
    InMux I__1398 (
            .O(N__6164),
            .I(N__6135));
    InMux I__1397 (
            .O(N__6163),
            .I(N__6135));
    Span4Mux_v I__1396 (
            .O(N__6160),
            .I(N__6132));
    Span4Mux_s3_v I__1395 (
            .O(N__6157),
            .I(N__6123));
    Span4Mux_h I__1394 (
            .O(N__6154),
            .I(N__6123));
    Span4Mux_h I__1393 (
            .O(N__6149),
            .I(N__6123));
    LocalMux I__1392 (
            .O(N__6146),
            .I(N__6123));
    LocalMux I__1391 (
            .O(N__6143),
            .I(N__6117));
    Span4Mux_h I__1390 (
            .O(N__6140),
            .I(N__6117));
    LocalMux I__1389 (
            .O(N__6135),
            .I(N__6110));
    Span4Mux_h I__1388 (
            .O(N__6132),
            .I(N__6110));
    Span4Mux_v I__1387 (
            .O(N__6123),
            .I(N__6110));
    InMux I__1386 (
            .O(N__6122),
            .I(N__6107));
    Span4Mux_v I__1385 (
            .O(N__6117),
            .I(N__6104));
    Span4Mux_v I__1384 (
            .O(N__6110),
            .I(N__6101));
    LocalMux I__1383 (
            .O(N__6107),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1382 (
            .O(N__6104),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1381 (
            .O(N__6101),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    InMux I__1380 (
            .O(N__6094),
            .I(N__6091));
    LocalMux I__1379 (
            .O(N__6091),
            .I(N__6088));
    IoSpan4Mux I__1378 (
            .O(N__6088),
            .I(N__6085));
    Odrv4 I__1377 (
            .O(N__6085),
            .I(A_c_15));
    InMux I__1376 (
            .O(N__6082),
            .I(N__6079));
    LocalMux I__1375 (
            .O(N__6079),
            .I(\U400_SDRAM.MA_5_iv_0_5 ));
    IoInMux I__1374 (
            .O(N__6076),
            .I(N__6073));
    LocalMux I__1373 (
            .O(N__6073),
            .I(N__6070));
    IoSpan4Mux I__1372 (
            .O(N__6070),
            .I(N__6067));
    IoSpan4Mux I__1371 (
            .O(N__6067),
            .I(N__6064));
    Odrv4 I__1370 (
            .O(N__6064),
            .I(MA_c_5));
    InMux I__1369 (
            .O(N__6061),
            .I(N__6058));
    LocalMux I__1368 (
            .O(N__6058),
            .I(N__6055));
    Odrv4 I__1367 (
            .O(N__6055),
            .I(A_c_5));
    CascadeMux I__1366 (
            .O(N__6052),
            .I(N__6049));
    InMux I__1365 (
            .O(N__6049),
            .I(N__6046));
    LocalMux I__1364 (
            .O(N__6046),
            .I(N__6043));
    Span4Mux_v I__1363 (
            .O(N__6043),
            .I(N__6040));
    Odrv4 I__1362 (
            .O(N__6040),
            .I(A_c_13));
    IoInMux I__1361 (
            .O(N__6037),
            .I(N__6034));
    LocalMux I__1360 (
            .O(N__6034),
            .I(N__6031));
    IoSpan4Mux I__1359 (
            .O(N__6031),
            .I(N__6028));
    Span4Mux_s3_h I__1358 (
            .O(N__6028),
            .I(N__6025));
    Span4Mux_h I__1357 (
            .O(N__6025),
            .I(N__6022));
    Odrv4 I__1356 (
            .O(N__6022),
            .I(MA_c_3));
    InMux I__1355 (
            .O(N__6019),
            .I(N__6016));
    LocalMux I__1354 (
            .O(N__6016),
            .I(N__6013));
    Span4Mux_s3_v I__1353 (
            .O(N__6013),
            .I(N__6010));
    Odrv4 I__1352 (
            .O(N__6010),
            .I(A_c_6));
    CascadeMux I__1351 (
            .O(N__6007),
            .I(N__6004));
    InMux I__1350 (
            .O(N__6004),
            .I(N__6001));
    LocalMux I__1349 (
            .O(N__6001),
            .I(N__5998));
    IoSpan4Mux I__1348 (
            .O(N__5998),
            .I(N__5995));
    Odrv4 I__1347 (
            .O(N__5995),
            .I(A_c_14));
    IoInMux I__1346 (
            .O(N__5992),
            .I(N__5989));
    LocalMux I__1345 (
            .O(N__5989),
            .I(N__5986));
    IoSpan4Mux I__1344 (
            .O(N__5986),
            .I(N__5983));
    Span4Mux_s1_v I__1343 (
            .O(N__5983),
            .I(N__5980));
    Span4Mux_h I__1342 (
            .O(N__5980),
            .I(N__5977));
    Odrv4 I__1341 (
            .O(N__5977),
            .I(MA_c_4));
    InMux I__1340 (
            .O(N__5974),
            .I(N__5971));
    LocalMux I__1339 (
            .O(N__5971),
            .I(N__5968));
    Span4Mux_h I__1338 (
            .O(N__5968),
            .I(N__5965));
    Odrv4 I__1337 (
            .O(N__5965),
            .I(A_c_2));
    CascadeMux I__1336 (
            .O(N__5962),
            .I(N__5959));
    InMux I__1335 (
            .O(N__5959),
            .I(N__5956));
    LocalMux I__1334 (
            .O(N__5956),
            .I(N__5953));
    Odrv4 I__1333 (
            .O(N__5953),
            .I(A_c_10));
    IoInMux I__1332 (
            .O(N__5950),
            .I(N__5947));
    LocalMux I__1331 (
            .O(N__5947),
            .I(N__5944));
    Span4Mux_s1_v I__1330 (
            .O(N__5944),
            .I(N__5941));
    Odrv4 I__1329 (
            .O(N__5941),
            .I(MA_c_0));
    InMux I__1328 (
            .O(N__5938),
            .I(N__5935));
    LocalMux I__1327 (
            .O(N__5935),
            .I(N__5932));
    Odrv4 I__1326 (
            .O(N__5932),
            .I(A_c_11));
    InMux I__1325 (
            .O(N__5929),
            .I(N__5926));
    LocalMux I__1324 (
            .O(N__5926),
            .I(\U400_SDRAM.MA_5_iv_0_1 ));
    InMux I__1323 (
            .O(N__5923),
            .I(N__5920));
    LocalMux I__1322 (
            .O(N__5920),
            .I(N__5917));
    Odrv4 I__1321 (
            .O(N__5917),
            .I(\U400_SDRAM.N_270 ));
    CascadeMux I__1320 (
            .O(N__5914),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_0_0_cascade_ ));
    InMux I__1319 (
            .O(N__5911),
            .I(N__5908));
    LocalMux I__1318 (
            .O(N__5908),
            .I(N__5905));
    Span4Mux_h I__1317 (
            .O(N__5905),
            .I(N__5900));
    InMux I__1316 (
            .O(N__5904),
            .I(N__5897));
    InMux I__1315 (
            .O(N__5903),
            .I(N__5894));
    Odrv4 I__1314 (
            .O(N__5900),
            .I(\U400_SDRAM.N_43 ));
    LocalMux I__1313 (
            .O(N__5897),
            .I(\U400_SDRAM.N_43 ));
    LocalMux I__1312 (
            .O(N__5894),
            .I(\U400_SDRAM.N_43 ));
    CascadeMux I__1311 (
            .O(N__5887),
            .I(N__5884));
    InMux I__1310 (
            .O(N__5884),
            .I(N__5881));
    LocalMux I__1309 (
            .O(N__5881),
            .I(N__5878));
    Span12Mux_v I__1308 (
            .O(N__5878),
            .I(N__5875));
    Odrv12 I__1307 (
            .O(N__5875),
            .I(A_c_25));
    IoInMux I__1306 (
            .O(N__5872),
            .I(N__5869));
    LocalMux I__1305 (
            .O(N__5869),
            .I(N__5866));
    Odrv12 I__1304 (
            .O(N__5866),
            .I(MA_c_11));
    IoInMux I__1303 (
            .O(N__5863),
            .I(N__5860));
    LocalMux I__1302 (
            .O(N__5860),
            .I(N__5857));
    Odrv4 I__1301 (
            .O(N__5857),
            .I(U400_BYTE_ENABLE_un1_UMBEn_i));
    IoInMux I__1300 (
            .O(N__5854),
            .I(N__5851));
    LocalMux I__1299 (
            .O(N__5851),
            .I(N__5848));
    Span4Mux_s2_v I__1298 (
            .O(N__5848),
            .I(N__5845));
    Odrv4 I__1297 (
            .O(N__5845),
            .I(U400_BYTE_ENABLE_un1_LMBEn_i));
    InMux I__1296 (
            .O(N__5842),
            .I(N__5832));
    InMux I__1295 (
            .O(N__5841),
            .I(N__5832));
    InMux I__1294 (
            .O(N__5840),
            .I(N__5832));
    InMux I__1293 (
            .O(N__5839),
            .I(N__5829));
    LocalMux I__1292 (
            .O(N__5832),
            .I(RAM_SPACEm));
    LocalMux I__1291 (
            .O(N__5829),
            .I(RAM_SPACEm));
    IoInMux I__1290 (
            .O(N__5824),
            .I(N__5821));
    LocalMux I__1289 (
            .O(N__5821),
            .I(N__5818));
    Span12Mux_s2_v I__1288 (
            .O(N__5818),
            .I(N__5815));
    Odrv12 I__1287 (
            .O(N__5815),
            .I(U400_BYTE_ENABLE_un1_UUBEn_i));
    InMux I__1286 (
            .O(N__5812),
            .I(N__5808));
    CascadeMux I__1285 (
            .O(N__5811),
            .I(N__5805));
    LocalMux I__1284 (
            .O(N__5808),
            .I(N__5800));
    InMux I__1283 (
            .O(N__5805),
            .I(N__5795));
    InMux I__1282 (
            .O(N__5804),
            .I(N__5795));
    InMux I__1281 (
            .O(N__5803),
            .I(N__5792));
    Span4Mux_v I__1280 (
            .O(N__5800),
            .I(N__5789));
    LocalMux I__1279 (
            .O(N__5795),
            .I(N__5784));
    LocalMux I__1278 (
            .O(N__5792),
            .I(N__5784));
    Sp12to4 I__1277 (
            .O(N__5789),
            .I(N__5781));
    Span4Mux_h I__1276 (
            .O(N__5784),
            .I(N__5778));
    Span12Mux_s6_h I__1275 (
            .O(N__5781),
            .I(N__5773));
    Sp12to4 I__1274 (
            .O(N__5778),
            .I(N__5773));
    Span12Mux_v I__1273 (
            .O(N__5773),
            .I(N__5770));
    Odrv12 I__1272 (
            .O(N__5770),
            .I(A_c_0));
    CascadeMux I__1271 (
            .O(N__5767),
            .I(N__5761));
    InMux I__1270 (
            .O(N__5766),
            .I(N__5752));
    InMux I__1269 (
            .O(N__5765),
            .I(N__5752));
    InMux I__1268 (
            .O(N__5764),
            .I(N__5752));
    InMux I__1267 (
            .O(N__5761),
            .I(N__5749));
    InMux I__1266 (
            .O(N__5760),
            .I(N__5744));
    InMux I__1265 (
            .O(N__5759),
            .I(N__5744));
    LocalMux I__1264 (
            .O(N__5752),
            .I(N__5737));
    LocalMux I__1263 (
            .O(N__5749),
            .I(N__5737));
    LocalMux I__1262 (
            .O(N__5744),
            .I(N__5737));
    Sp12to4 I__1261 (
            .O(N__5737),
            .I(N__5734));
    Span12Mux_v I__1260 (
            .O(N__5734),
            .I(N__5731));
    Odrv12 I__1259 (
            .O(N__5731),
            .I(A_c_1));
    InMux I__1258 (
            .O(N__5728),
            .I(N__5725));
    LocalMux I__1257 (
            .O(N__5725),
            .I(\U400_BYTE_ENABLE.un2_UMBEn_0_0 ));
    CascadeMux I__1256 (
            .O(N__5722),
            .I(N__5718));
    InMux I__1255 (
            .O(N__5721),
            .I(N__5713));
    InMux I__1254 (
            .O(N__5718),
            .I(N__5713));
    LocalMux I__1253 (
            .O(N__5713),
            .I(\U400_BYTE_ENABLE.LW_TRANS_0 ));
    CascadeMux I__1252 (
            .O(N__5710),
            .I(N__5706));
    InMux I__1251 (
            .O(N__5709),
            .I(N__5702));
    InMux I__1250 (
            .O(N__5706),
            .I(N__5699));
    InMux I__1249 (
            .O(N__5705),
            .I(N__5696));
    LocalMux I__1248 (
            .O(N__5702),
            .I(N__5693));
    LocalMux I__1247 (
            .O(N__5699),
            .I(N__5690));
    LocalMux I__1246 (
            .O(N__5696),
            .I(N__5687));
    Span4Mux_v I__1245 (
            .O(N__5693),
            .I(N__5684));
    Span4Mux_v I__1244 (
            .O(N__5690),
            .I(N__5681));
    Span12Mux_v I__1243 (
            .O(N__5687),
            .I(N__5676));
    Sp12to4 I__1242 (
            .O(N__5684),
            .I(N__5676));
    Odrv4 I__1241 (
            .O(N__5681),
            .I(U400_ADDRESS_DECODE_RAM_SPACE_3));
    Odrv12 I__1240 (
            .O(N__5676),
            .I(U400_ADDRESS_DECODE_RAM_SPACE_3));
    InMux I__1239 (
            .O(N__5671),
            .I(N__5666));
    InMux I__1238 (
            .O(N__5670),
            .I(N__5663));
    InMux I__1237 (
            .O(N__5669),
            .I(N__5660));
    LocalMux I__1236 (
            .O(N__5666),
            .I(N__5657));
    LocalMux I__1235 (
            .O(N__5663),
            .I(N__5654));
    LocalMux I__1234 (
            .O(N__5660),
            .I(N__5651));
    Span4Mux_h I__1233 (
            .O(N__5657),
            .I(N__5648));
    Span4Mux_v I__1232 (
            .O(N__5654),
            .I(N__5643));
    Span4Mux_h I__1231 (
            .O(N__5651),
            .I(N__5643));
    Span4Mux_h I__1230 (
            .O(N__5648),
            .I(N__5640));
    IoSpan4Mux I__1229 (
            .O(N__5643),
            .I(N__5637));
    Odrv4 I__1228 (
            .O(N__5640),
            .I(A_c_29));
    Odrv4 I__1227 (
            .O(N__5637),
            .I(A_c_29));
    InMux I__1226 (
            .O(N__5632),
            .I(N__5628));
    InMux I__1225 (
            .O(N__5631),
            .I(N__5624));
    LocalMux I__1224 (
            .O(N__5628),
            .I(N__5621));
    InMux I__1223 (
            .O(N__5627),
            .I(N__5618));
    LocalMux I__1222 (
            .O(N__5624),
            .I(N__5615));
    Span4Mux_v I__1221 (
            .O(N__5621),
            .I(N__5610));
    LocalMux I__1220 (
            .O(N__5618),
            .I(N__5610));
    Span12Mux_s8_h I__1219 (
            .O(N__5615),
            .I(N__5607));
    Span4Mux_h I__1218 (
            .O(N__5610),
            .I(N__5604));
    Odrv12 I__1217 (
            .O(N__5607),
            .I(A_c_28));
    Odrv4 I__1216 (
            .O(N__5604),
            .I(A_c_28));
    IoInMux I__1215 (
            .O(N__5599),
            .I(N__5596));
    LocalMux I__1214 (
            .O(N__5596),
            .I(N__5593));
    Span4Mux_s3_h I__1213 (
            .O(N__5593),
            .I(N__5590));
    Odrv4 I__1212 (
            .O(N__5590),
            .I(RAM_SPACEm_i));
    CascadeMux I__1211 (
            .O(N__5587),
            .I(N__5582));
    CascadeMux I__1210 (
            .O(N__5586),
            .I(N__5578));
    CascadeMux I__1209 (
            .O(N__5585),
            .I(N__5574));
    InMux I__1208 (
            .O(N__5582),
            .I(N__5569));
    InMux I__1207 (
            .O(N__5581),
            .I(N__5569));
    InMux I__1206 (
            .O(N__5578),
            .I(N__5566));
    CascadeMux I__1205 (
            .O(N__5577),
            .I(N__5562));
    InMux I__1204 (
            .O(N__5574),
            .I(N__5558));
    LocalMux I__1203 (
            .O(N__5569),
            .I(N__5553));
    LocalMux I__1202 (
            .O(N__5566),
            .I(N__5553));
    InMux I__1201 (
            .O(N__5565),
            .I(N__5548));
    InMux I__1200 (
            .O(N__5562),
            .I(N__5548));
    InMux I__1199 (
            .O(N__5561),
            .I(N__5545));
    LocalMux I__1198 (
            .O(N__5558),
            .I(N__5542));
    Span4Mux_h I__1197 (
            .O(N__5553),
            .I(N__5535));
    LocalMux I__1196 (
            .O(N__5548),
            .I(N__5535));
    LocalMux I__1195 (
            .O(N__5545),
            .I(N__5535));
    Span12Mux_s6_v I__1194 (
            .O(N__5542),
            .I(N__5532));
    Span4Mux_v I__1193 (
            .O(N__5535),
            .I(N__5529));
    Odrv12 I__1192 (
            .O(N__5532),
            .I(SIZ_c_1));
    Odrv4 I__1191 (
            .O(N__5529),
            .I(SIZ_c_1));
    InMux I__1190 (
            .O(N__5524),
            .I(N__5510));
    InMux I__1189 (
            .O(N__5523),
            .I(N__5510));
    InMux I__1188 (
            .O(N__5522),
            .I(N__5510));
    InMux I__1187 (
            .O(N__5521),
            .I(N__5503));
    InMux I__1186 (
            .O(N__5520),
            .I(N__5503));
    InMux I__1185 (
            .O(N__5519),
            .I(N__5503));
    InMux I__1184 (
            .O(N__5518),
            .I(N__5498));
    InMux I__1183 (
            .O(N__5517),
            .I(N__5498));
    LocalMux I__1182 (
            .O(N__5510),
            .I(\U400_SDRAM.N_303_0_i ));
    LocalMux I__1181 (
            .O(N__5503),
            .I(\U400_SDRAM.N_303_0_i ));
    LocalMux I__1180 (
            .O(N__5498),
            .I(\U400_SDRAM.N_303_0_i ));
    InMux I__1179 (
            .O(N__5491),
            .I(N__5485));
    InMux I__1178 (
            .O(N__5490),
            .I(N__5485));
    LocalMux I__1177 (
            .O(N__5485),
            .I(\U400_SDRAM.SDRAM_CMD_5_sqmuxa ));
    InMux I__1176 (
            .O(N__5482),
            .I(N__5479));
    LocalMux I__1175 (
            .O(N__5479),
            .I(N__5476));
    Span4Mux_v I__1174 (
            .O(N__5476),
            .I(N__5473));
    Odrv4 I__1173 (
            .O(N__5473),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_1 ));
    CEMux I__1172 (
            .O(N__5470),
            .I(N__5466));
    CEMux I__1171 (
            .O(N__5469),
            .I(N__5463));
    LocalMux I__1170 (
            .O(N__5466),
            .I(N__5460));
    LocalMux I__1169 (
            .O(N__5463),
            .I(N__5457));
    Span4Mux_h I__1168 (
            .O(N__5460),
            .I(N__5454));
    Span4Mux_v I__1167 (
            .O(N__5457),
            .I(N__5451));
    Odrv4 I__1166 (
            .O(N__5454),
            .I(\U400_SDRAM.SDRAM_COUNTERe_0_i ));
    Odrv4 I__1165 (
            .O(N__5451),
            .I(\U400_SDRAM.SDRAM_COUNTERe_0_i ));
    InMux I__1164 (
            .O(N__5446),
            .I(N__5441));
    InMux I__1163 (
            .O(N__5445),
            .I(N__5436));
    InMux I__1162 (
            .O(N__5444),
            .I(N__5436));
    LocalMux I__1161 (
            .O(N__5441),
            .I(\U400_SDRAM.N_66 ));
    LocalMux I__1160 (
            .O(N__5436),
            .I(\U400_SDRAM.N_66 ));
    InMux I__1159 (
            .O(N__5431),
            .I(N__5427));
    InMux I__1158 (
            .O(N__5430),
            .I(N__5422));
    LocalMux I__1157 (
            .O(N__5427),
            .I(N__5419));
    InMux I__1156 (
            .O(N__5426),
            .I(N__5416));
    InMux I__1155 (
            .O(N__5425),
            .I(N__5413));
    LocalMux I__1154 (
            .O(N__5422),
            .I(\U400_SDRAM.N_55 ));
    Odrv4 I__1153 (
            .O(N__5419),
            .I(\U400_SDRAM.N_55 ));
    LocalMux I__1152 (
            .O(N__5416),
            .I(\U400_SDRAM.N_55 ));
    LocalMux I__1151 (
            .O(N__5413),
            .I(\U400_SDRAM.N_55 ));
    InMux I__1150 (
            .O(N__5404),
            .I(N__5400));
    InMux I__1149 (
            .O(N__5403),
            .I(N__5397));
    LocalMux I__1148 (
            .O(N__5400),
            .I(N__5394));
    LocalMux I__1147 (
            .O(N__5397),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa ));
    Odrv4 I__1146 (
            .O(N__5394),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa ));
    CascadeMux I__1145 (
            .O(N__5389),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_cascade_ ));
    InMux I__1144 (
            .O(N__5386),
            .I(N__5383));
    LocalMux I__1143 (
            .O(N__5383),
            .I(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_1_0 ));
    InMux I__1142 (
            .O(N__5380),
            .I(N__5377));
    LocalMux I__1141 (
            .O(N__5377),
            .I(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_0 ));
    InMux I__1140 (
            .O(N__5374),
            .I(N__5367));
    InMux I__1139 (
            .O(N__5373),
            .I(N__5360));
    InMux I__1138 (
            .O(N__5372),
            .I(N__5360));
    InMux I__1137 (
            .O(N__5371),
            .I(N__5360));
    InMux I__1136 (
            .O(N__5370),
            .I(N__5356));
    LocalMux I__1135 (
            .O(N__5367),
            .I(N__5353));
    LocalMux I__1134 (
            .O(N__5360),
            .I(N__5350));
    InMux I__1133 (
            .O(N__5359),
            .I(N__5347));
    LocalMux I__1132 (
            .O(N__5356),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ));
    Odrv4 I__1131 (
            .O(N__5353),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ));
    Odrv4 I__1130 (
            .O(N__5350),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ));
    LocalMux I__1129 (
            .O(N__5347),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ));
    InMux I__1128 (
            .O(N__5338),
            .I(N__5326));
    InMux I__1127 (
            .O(N__5337),
            .I(N__5321));
    InMux I__1126 (
            .O(N__5336),
            .I(N__5321));
    InMux I__1125 (
            .O(N__5335),
            .I(N__5316));
    InMux I__1124 (
            .O(N__5334),
            .I(N__5316));
    CascadeMux I__1123 (
            .O(N__5333),
            .I(N__5311));
    InMux I__1122 (
            .O(N__5332),
            .I(N__5305));
    CascadeMux I__1121 (
            .O(N__5331),
            .I(N__5300));
    InMux I__1120 (
            .O(N__5330),
            .I(N__5295));
    InMux I__1119 (
            .O(N__5329),
            .I(N__5295));
    LocalMux I__1118 (
            .O(N__5326),
            .I(N__5292));
    LocalMux I__1117 (
            .O(N__5321),
            .I(N__5287));
    LocalMux I__1116 (
            .O(N__5316),
            .I(N__5287));
    InMux I__1115 (
            .O(N__5315),
            .I(N__5282));
    InMux I__1114 (
            .O(N__5314),
            .I(N__5282));
    InMux I__1113 (
            .O(N__5311),
            .I(N__5279));
    InMux I__1112 (
            .O(N__5310),
            .I(N__5276));
    InMux I__1111 (
            .O(N__5309),
            .I(N__5271));
    InMux I__1110 (
            .O(N__5308),
            .I(N__5271));
    LocalMux I__1109 (
            .O(N__5305),
            .I(N__5268));
    InMux I__1108 (
            .O(N__5304),
            .I(N__5261));
    InMux I__1107 (
            .O(N__5303),
            .I(N__5261));
    InMux I__1106 (
            .O(N__5300),
            .I(N__5261));
    LocalMux I__1105 (
            .O(N__5295),
            .I(N__5258));
    Span4Mux_v I__1104 (
            .O(N__5292),
            .I(N__5251));
    Span4Mux_v I__1103 (
            .O(N__5287),
            .I(N__5251));
    LocalMux I__1102 (
            .O(N__5282),
            .I(N__5251));
    LocalMux I__1101 (
            .O(N__5279),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1100 (
            .O(N__5276),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1099 (
            .O(N__5271),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1098 (
            .O(N__5268),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1097 (
            .O(N__5261),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1096 (
            .O(N__5258),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1095 (
            .O(N__5251),
            .I(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__1094 (
            .O(N__5236),
            .I(N__5230));
    InMux I__1093 (
            .O(N__5235),
            .I(N__5224));
    InMux I__1092 (
            .O(N__5234),
            .I(N__5217));
    InMux I__1091 (
            .O(N__5233),
            .I(N__5217));
    InMux I__1090 (
            .O(N__5230),
            .I(N__5217));
    InMux I__1089 (
            .O(N__5229),
            .I(N__5214));
    CascadeMux I__1088 (
            .O(N__5228),
            .I(N__5204));
    InMux I__1087 (
            .O(N__5227),
            .I(N__5200));
    LocalMux I__1086 (
            .O(N__5224),
            .I(N__5193));
    LocalMux I__1085 (
            .O(N__5217),
            .I(N__5193));
    LocalMux I__1084 (
            .O(N__5214),
            .I(N__5193));
    InMux I__1083 (
            .O(N__5213),
            .I(N__5190));
    InMux I__1082 (
            .O(N__5212),
            .I(N__5186));
    InMux I__1081 (
            .O(N__5211),
            .I(N__5183));
    InMux I__1080 (
            .O(N__5210),
            .I(N__5176));
    InMux I__1079 (
            .O(N__5209),
            .I(N__5176));
    InMux I__1078 (
            .O(N__5208),
            .I(N__5171));
    InMux I__1077 (
            .O(N__5207),
            .I(N__5171));
    InMux I__1076 (
            .O(N__5204),
            .I(N__5168));
    InMux I__1075 (
            .O(N__5203),
            .I(N__5165));
    LocalMux I__1074 (
            .O(N__5200),
            .I(N__5161));
    Span4Mux_v I__1073 (
            .O(N__5193),
            .I(N__5156));
    LocalMux I__1072 (
            .O(N__5190),
            .I(N__5156));
    InMux I__1071 (
            .O(N__5189),
            .I(N__5153));
    LocalMux I__1070 (
            .O(N__5186),
            .I(N__5148));
    LocalMux I__1069 (
            .O(N__5183),
            .I(N__5148));
    InMux I__1068 (
            .O(N__5182),
            .I(N__5145));
    InMux I__1067 (
            .O(N__5181),
            .I(N__5142));
    LocalMux I__1066 (
            .O(N__5176),
            .I(N__5135));
    LocalMux I__1065 (
            .O(N__5171),
            .I(N__5135));
    LocalMux I__1064 (
            .O(N__5168),
            .I(N__5135));
    LocalMux I__1063 (
            .O(N__5165),
            .I(N__5132));
    InMux I__1062 (
            .O(N__5164),
            .I(N__5129));
    Span4Mux_v I__1061 (
            .O(N__5161),
            .I(N__5126));
    Span4Mux_v I__1060 (
            .O(N__5156),
            .I(N__5123));
    LocalMux I__1059 (
            .O(N__5153),
            .I(N__5120));
    Span4Mux_v I__1058 (
            .O(N__5148),
            .I(N__5113));
    LocalMux I__1057 (
            .O(N__5145),
            .I(N__5113));
    LocalMux I__1056 (
            .O(N__5142),
            .I(N__5113));
    Span4Mux_h I__1055 (
            .O(N__5135),
            .I(N__5106));
    Span4Mux_h I__1054 (
            .O(N__5132),
            .I(N__5106));
    LocalMux I__1053 (
            .O(N__5129),
            .I(N__5106));
    Span4Mux_h I__1052 (
            .O(N__5126),
            .I(N__5099));
    Span4Mux_h I__1051 (
            .O(N__5123),
            .I(N__5099));
    Span4Mux_v I__1050 (
            .O(N__5120),
            .I(N__5099));
    Span4Mux_v I__1049 (
            .O(N__5113),
            .I(N__5096));
    Span4Mux_v I__1048 (
            .O(N__5106),
            .I(N__5093));
    Span4Mux_h I__1047 (
            .O(N__5099),
            .I(N__5090));
    Span4Mux_h I__1046 (
            .O(N__5096),
            .I(N__5087));
    Span4Mux_h I__1045 (
            .O(N__5093),
            .I(N__5084));
    Odrv4 I__1044 (
            .O(N__5090),
            .I(RESETn_c));
    Odrv4 I__1043 (
            .O(N__5087),
            .I(RESETn_c));
    Odrv4 I__1042 (
            .O(N__5084),
            .I(RESETn_c));
    InMux I__1041 (
            .O(N__5077),
            .I(N__5069));
    InMux I__1040 (
            .O(N__5076),
            .I(N__5069));
    CascadeMux I__1039 (
            .O(N__5075),
            .I(N__5063));
    InMux I__1038 (
            .O(N__5074),
            .I(N__5053));
    LocalMux I__1037 (
            .O(N__5069),
            .I(N__5050));
    InMux I__1036 (
            .O(N__5068),
            .I(N__5047));
    InMux I__1035 (
            .O(N__5067),
            .I(N__5044));
    InMux I__1034 (
            .O(N__5066),
            .I(N__5041));
    InMux I__1033 (
            .O(N__5063),
            .I(N__5036));
    InMux I__1032 (
            .O(N__5062),
            .I(N__5031));
    InMux I__1031 (
            .O(N__5061),
            .I(N__5031));
    InMux I__1030 (
            .O(N__5060),
            .I(N__5024));
    InMux I__1029 (
            .O(N__5059),
            .I(N__5024));
    InMux I__1028 (
            .O(N__5058),
            .I(N__5024));
    InMux I__1027 (
            .O(N__5057),
            .I(N__5021));
    InMux I__1026 (
            .O(N__5056),
            .I(N__5018));
    LocalMux I__1025 (
            .O(N__5053),
            .I(N__5007));
    Span4Mux_v I__1024 (
            .O(N__5050),
            .I(N__5007));
    LocalMux I__1023 (
            .O(N__5047),
            .I(N__5007));
    LocalMux I__1022 (
            .O(N__5044),
            .I(N__5007));
    LocalMux I__1021 (
            .O(N__5041),
            .I(N__5007));
    InMux I__1020 (
            .O(N__5040),
            .I(N__5004));
    InMux I__1019 (
            .O(N__5039),
            .I(N__5001));
    LocalMux I__1018 (
            .O(N__5036),
            .I(N__4994));
    LocalMux I__1017 (
            .O(N__5031),
            .I(N__4994));
    LocalMux I__1016 (
            .O(N__5024),
            .I(N__4994));
    LocalMux I__1015 (
            .O(N__5021),
            .I(N__4991));
    LocalMux I__1014 (
            .O(N__5018),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1013 (
            .O(N__5007),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1012 (
            .O(N__5004),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1011 (
            .O(N__5001),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1010 (
            .O(N__4994),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1009 (
            .O(N__4991),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1008 (
            .O(N__4978),
            .I(N__4968));
    InMux I__1007 (
            .O(N__4977),
            .I(N__4965));
    InMux I__1006 (
            .O(N__4976),
            .I(N__4958));
    InMux I__1005 (
            .O(N__4975),
            .I(N__4953));
    InMux I__1004 (
            .O(N__4974),
            .I(N__4953));
    InMux I__1003 (
            .O(N__4973),
            .I(N__4947));
    InMux I__1002 (
            .O(N__4972),
            .I(N__4947));
    InMux I__1001 (
            .O(N__4971),
            .I(N__4941));
    LocalMux I__1000 (
            .O(N__4968),
            .I(N__4936));
    LocalMux I__999 (
            .O(N__4965),
            .I(N__4936));
    InMux I__998 (
            .O(N__4964),
            .I(N__4929));
    InMux I__997 (
            .O(N__4963),
            .I(N__4929));
    InMux I__996 (
            .O(N__4962),
            .I(N__4929));
    CascadeMux I__995 (
            .O(N__4961),
            .I(N__4926));
    LocalMux I__994 (
            .O(N__4958),
            .I(N__4919));
    LocalMux I__993 (
            .O(N__4953),
            .I(N__4919));
    InMux I__992 (
            .O(N__4952),
            .I(N__4914));
    LocalMux I__991 (
            .O(N__4947),
            .I(N__4911));
    InMux I__990 (
            .O(N__4946),
            .I(N__4904));
    InMux I__989 (
            .O(N__4945),
            .I(N__4904));
    InMux I__988 (
            .O(N__4944),
            .I(N__4904));
    LocalMux I__987 (
            .O(N__4941),
            .I(N__4897));
    Span4Mux_h I__986 (
            .O(N__4936),
            .I(N__4897));
    LocalMux I__985 (
            .O(N__4929),
            .I(N__4897));
    InMux I__984 (
            .O(N__4926),
            .I(N__4890));
    InMux I__983 (
            .O(N__4925),
            .I(N__4890));
    InMux I__982 (
            .O(N__4924),
            .I(N__4890));
    Span4Mux_v I__981 (
            .O(N__4919),
            .I(N__4887));
    InMux I__980 (
            .O(N__4918),
            .I(N__4882));
    InMux I__979 (
            .O(N__4917),
            .I(N__4882));
    LocalMux I__978 (
            .O(N__4914),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__977 (
            .O(N__4911),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__976 (
            .O(N__4904),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__975 (
            .O(N__4897),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__974 (
            .O(N__4890),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__973 (
            .O(N__4887),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__972 (
            .O(N__4882),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__971 (
            .O(N__4867),
            .I(N__4861));
    CascadeMux I__970 (
            .O(N__4866),
            .I(N__4858));
    CascadeMux I__969 (
            .O(N__4865),
            .I(N__4853));
    CascadeMux I__968 (
            .O(N__4864),
            .I(N__4849));
    LocalMux I__967 (
            .O(N__4861),
            .I(N__4842));
    InMux I__966 (
            .O(N__4858),
            .I(N__4839));
    CascadeMux I__965 (
            .O(N__4857),
            .I(N__4834));
    InMux I__964 (
            .O(N__4856),
            .I(N__4828));
    InMux I__963 (
            .O(N__4853),
            .I(N__4828));
    InMux I__962 (
            .O(N__4852),
            .I(N__4825));
    InMux I__961 (
            .O(N__4849),
            .I(N__4822));
    InMux I__960 (
            .O(N__4848),
            .I(N__4819));
    InMux I__959 (
            .O(N__4847),
            .I(N__4814));
    InMux I__958 (
            .O(N__4846),
            .I(N__4814));
    InMux I__957 (
            .O(N__4845),
            .I(N__4811));
    Span4Mux_v I__956 (
            .O(N__4842),
            .I(N__4805));
    LocalMux I__955 (
            .O(N__4839),
            .I(N__4805));
    InMux I__954 (
            .O(N__4838),
            .I(N__4802));
    InMux I__953 (
            .O(N__4837),
            .I(N__4799));
    InMux I__952 (
            .O(N__4834),
            .I(N__4793));
    InMux I__951 (
            .O(N__4833),
            .I(N__4793));
    LocalMux I__950 (
            .O(N__4828),
            .I(N__4785));
    LocalMux I__949 (
            .O(N__4825),
            .I(N__4785));
    LocalMux I__948 (
            .O(N__4822),
            .I(N__4778));
    LocalMux I__947 (
            .O(N__4819),
            .I(N__4778));
    LocalMux I__946 (
            .O(N__4814),
            .I(N__4778));
    LocalMux I__945 (
            .O(N__4811),
            .I(N__4775));
    CascadeMux I__944 (
            .O(N__4810),
            .I(N__4771));
    Span4Mux_v I__943 (
            .O(N__4805),
            .I(N__4763));
    LocalMux I__942 (
            .O(N__4802),
            .I(N__4763));
    LocalMux I__941 (
            .O(N__4799),
            .I(N__4763));
    InMux I__940 (
            .O(N__4798),
            .I(N__4760));
    LocalMux I__939 (
            .O(N__4793),
            .I(N__4757));
    InMux I__938 (
            .O(N__4792),
            .I(N__4750));
    InMux I__937 (
            .O(N__4791),
            .I(N__4750));
    InMux I__936 (
            .O(N__4790),
            .I(N__4750));
    Span4Mux_v I__935 (
            .O(N__4785),
            .I(N__4743));
    Span4Mux_h I__934 (
            .O(N__4778),
            .I(N__4743));
    Span4Mux_v I__933 (
            .O(N__4775),
            .I(N__4743));
    InMux I__932 (
            .O(N__4774),
            .I(N__4736));
    InMux I__931 (
            .O(N__4771),
            .I(N__4736));
    InMux I__930 (
            .O(N__4770),
            .I(N__4736));
    Span4Mux_h I__929 (
            .O(N__4763),
            .I(N__4733));
    LocalMux I__928 (
            .O(N__4760),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__927 (
            .O(N__4757),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__926 (
            .O(N__4750),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__925 (
            .O(N__4743),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__924 (
            .O(N__4736),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__923 (
            .O(N__4733),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ));
    CascadeMux I__922 (
            .O(N__4720),
            .I(N__4708));
    CascadeMux I__921 (
            .O(N__4719),
            .I(N__4705));
    InMux I__920 (
            .O(N__4718),
            .I(N__4702));
    InMux I__919 (
            .O(N__4717),
            .I(N__4699));
    InMux I__918 (
            .O(N__4716),
            .I(N__4694));
    InMux I__917 (
            .O(N__4715),
            .I(N__4694));
    InMux I__916 (
            .O(N__4714),
            .I(N__4688));
    InMux I__915 (
            .O(N__4713),
            .I(N__4684));
    InMux I__914 (
            .O(N__4712),
            .I(N__4681));
    InMux I__913 (
            .O(N__4711),
            .I(N__4674));
    InMux I__912 (
            .O(N__4708),
            .I(N__4674));
    InMux I__911 (
            .O(N__4705),
            .I(N__4674));
    LocalMux I__910 (
            .O(N__4702),
            .I(N__4665));
    LocalMux I__909 (
            .O(N__4699),
            .I(N__4665));
    LocalMux I__908 (
            .O(N__4694),
            .I(N__4665));
    InMux I__907 (
            .O(N__4693),
            .I(N__4660));
    InMux I__906 (
            .O(N__4692),
            .I(N__4660));
    InMux I__905 (
            .O(N__4691),
            .I(N__4657));
    LocalMux I__904 (
            .O(N__4688),
            .I(N__4654));
    InMux I__903 (
            .O(N__4687),
            .I(N__4651));
    LocalMux I__902 (
            .O(N__4684),
            .I(N__4648));
    LocalMux I__901 (
            .O(N__4681),
            .I(N__4643));
    LocalMux I__900 (
            .O(N__4674),
            .I(N__4640));
    InMux I__899 (
            .O(N__4673),
            .I(N__4632));
    InMux I__898 (
            .O(N__4672),
            .I(N__4632));
    Span4Mux_v I__897 (
            .O(N__4665),
            .I(N__4627));
    LocalMux I__896 (
            .O(N__4660),
            .I(N__4627));
    LocalMux I__895 (
            .O(N__4657),
            .I(N__4618));
    Span4Mux_h I__894 (
            .O(N__4654),
            .I(N__4618));
    LocalMux I__893 (
            .O(N__4651),
            .I(N__4618));
    Span4Mux_h I__892 (
            .O(N__4648),
            .I(N__4618));
    InMux I__891 (
            .O(N__4647),
            .I(N__4613));
    InMux I__890 (
            .O(N__4646),
            .I(N__4613));
    Span4Mux_v I__889 (
            .O(N__4643),
            .I(N__4608));
    Span4Mux_h I__888 (
            .O(N__4640),
            .I(N__4608));
    InMux I__887 (
            .O(N__4639),
            .I(N__4603));
    InMux I__886 (
            .O(N__4638),
            .I(N__4603));
    InMux I__885 (
            .O(N__4637),
            .I(N__4600));
    LocalMux I__884 (
            .O(N__4632),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__883 (
            .O(N__4627),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__882 (
            .O(N__4618),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__881 (
            .O(N__4613),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__880 (
            .O(N__4608),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__879 (
            .O(N__4603),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__878 (
            .O(N__4600),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__877 (
            .O(N__4585),
            .I(N__4582));
    LocalMux I__876 (
            .O(N__4582),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_a5_0_0 ));
    CascadeMux I__875 (
            .O(N__4579),
            .I(N__4576));
    InMux I__874 (
            .O(N__4576),
            .I(N__4573));
    LocalMux I__873 (
            .O(N__4573),
            .I(N__4569));
    InMux I__872 (
            .O(N__4572),
            .I(N__4566));
    Span4Mux_h I__871 (
            .O(N__4569),
            .I(N__4563));
    LocalMux I__870 (
            .O(N__4566),
            .I(\U400_SDRAM.N_299_2 ));
    Odrv4 I__869 (
            .O(N__4563),
            .I(\U400_SDRAM.N_299_2 ));
    CascadeMux I__868 (
            .O(N__4558),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_0_tz_cascade_ ));
    CascadeMux I__867 (
            .O(N__4555),
            .I(N__4550));
    CascadeMux I__866 (
            .O(N__4554),
            .I(N__4547));
    InMux I__865 (
            .O(N__4553),
            .I(N__4543));
    InMux I__864 (
            .O(N__4550),
            .I(N__4536));
    InMux I__863 (
            .O(N__4547),
            .I(N__4536));
    InMux I__862 (
            .O(N__4546),
            .I(N__4536));
    LocalMux I__861 (
            .O(N__4543),
            .I(N__4533));
    LocalMux I__860 (
            .O(N__4536),
            .I(N__4530));
    Odrv4 I__859 (
            .O(N__4533),
            .I(\U400_SDRAM.N_266_0 ));
    Odrv4 I__858 (
            .O(N__4530),
            .I(\U400_SDRAM.N_266_0 ));
    CascadeMux I__857 (
            .O(N__4525),
            .I(\U400_BYTE_ENABLE.un2_LLBEn_0_0_cascade_ ));
    IoInMux I__856 (
            .O(N__4522),
            .I(N__4519));
    LocalMux I__855 (
            .O(N__4519),
            .I(N__4516));
    Span4Mux_s2_v I__854 (
            .O(N__4516),
            .I(N__4513));
    Odrv4 I__853 (
            .O(N__4513),
            .I(U400_BYTE_ENABLE_un1_LLBEn_i));
    InMux I__852 (
            .O(N__4510),
            .I(N__4507));
    LocalMux I__851 (
            .O(N__4507),
            .I(N__4504));
    Odrv12 I__850 (
            .O(N__4504),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_76_i_a4_0 ));
    CascadeMux I__849 (
            .O(N__4501),
            .I(\U400_SDRAM.N_321_0_cascade_ ));
    InMux I__848 (
            .O(N__4498),
            .I(N__4495));
    LocalMux I__847 (
            .O(N__4495),
            .I(\U400_SDRAM.N_322_0 ));
    CascadeMux I__846 (
            .O(N__4492),
            .I(N__4485));
    InMux I__845 (
            .O(N__4491),
            .I(N__4480));
    InMux I__844 (
            .O(N__4490),
            .I(N__4477));
    InMux I__843 (
            .O(N__4489),
            .I(N__4474));
    InMux I__842 (
            .O(N__4488),
            .I(N__4469));
    InMux I__841 (
            .O(N__4485),
            .I(N__4469));
    CascadeMux I__840 (
            .O(N__4484),
            .I(N__4466));
    InMux I__839 (
            .O(N__4483),
            .I(N__4463));
    LocalMux I__838 (
            .O(N__4480),
            .I(N__4460));
    LocalMux I__837 (
            .O(N__4477),
            .I(N__4453));
    LocalMux I__836 (
            .O(N__4474),
            .I(N__4453));
    LocalMux I__835 (
            .O(N__4469),
            .I(N__4453));
    InMux I__834 (
            .O(N__4466),
            .I(N__4450));
    LocalMux I__833 (
            .O(N__4463),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    Odrv4 I__832 (
            .O(N__4460),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    Odrv4 I__831 (
            .O(N__4453),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    LocalMux I__830 (
            .O(N__4450),
            .I(\U400_SDRAM.WRITE_CYCLEZ0 ));
    InMux I__829 (
            .O(N__4441),
            .I(N__4438));
    LocalMux I__828 (
            .O(N__4438),
            .I(\U400_SDRAM.N_320_0 ));
    CascadeMux I__827 (
            .O(N__4435),
            .I(N__4432));
    InMux I__826 (
            .O(N__4432),
            .I(N__4429));
    LocalMux I__825 (
            .O(N__4429),
            .I(N__4426));
    Span4Mux_h I__824 (
            .O(N__4426),
            .I(N__4423));
    Odrv4 I__823 (
            .O(N__4423),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_0 ));
    InMux I__822 (
            .O(N__4420),
            .I(N__4417));
    LocalMux I__821 (
            .O(N__4417),
            .I(\U400_SDRAM.N_88 ));
    InMux I__820 (
            .O(N__4414),
            .I(N__4411));
    LocalMux I__819 (
            .O(N__4411),
            .I(N__4408));
    Span4Mux_h I__818 (
            .O(N__4408),
            .I(N__4405));
    Odrv4 I__817 (
            .O(N__4405),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_3 ));
    InMux I__816 (
            .O(N__4402),
            .I(N__4399));
    LocalMux I__815 (
            .O(N__4399),
            .I(N__4396));
    Span4Mux_v I__814 (
            .O(N__4396),
            .I(N__4393));
    Odrv4 I__813 (
            .O(N__4393),
            .I(\U400_SDRAM.N_56 ));
    CascadeMux I__812 (
            .O(N__4390),
            .I(\U400_SDRAM.N_56_cascade_ ));
    InMux I__811 (
            .O(N__4387),
            .I(N__4383));
    InMux I__810 (
            .O(N__4386),
            .I(N__4380));
    LocalMux I__809 (
            .O(N__4383),
            .I(\U400_SDRAM.N_108 ));
    LocalMux I__808 (
            .O(N__4380),
            .I(\U400_SDRAM.N_108 ));
    CascadeMux I__807 (
            .O(N__4375),
            .I(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_o2_0_0_cascade_ ));
    InMux I__806 (
            .O(N__4372),
            .I(N__4368));
    InMux I__805 (
            .O(N__4371),
            .I(N__4362));
    LocalMux I__804 (
            .O(N__4368),
            .I(N__4359));
    InMux I__803 (
            .O(N__4367),
            .I(N__4354));
    InMux I__802 (
            .O(N__4366),
            .I(N__4354));
    InMux I__801 (
            .O(N__4365),
            .I(N__4351));
    LocalMux I__800 (
            .O(N__4362),
            .I(\U400_SDRAM.N_94_1 ));
    Odrv4 I__799 (
            .O(N__4359),
            .I(\U400_SDRAM.N_94_1 ));
    LocalMux I__798 (
            .O(N__4354),
            .I(\U400_SDRAM.N_94_1 ));
    LocalMux I__797 (
            .O(N__4351),
            .I(\U400_SDRAM.N_94_1 ));
    CascadeMux I__796 (
            .O(N__4342),
            .I(\U400_SDRAM.N_275_cascade_ ));
    InMux I__795 (
            .O(N__4339),
            .I(N__4332));
    InMux I__794 (
            .O(N__4338),
            .I(N__4332));
    InMux I__793 (
            .O(N__4337),
            .I(N__4323));
    LocalMux I__792 (
            .O(N__4332),
            .I(N__4320));
    InMux I__791 (
            .O(N__4331),
            .I(N__4315));
    InMux I__790 (
            .O(N__4330),
            .I(N__4315));
    InMux I__789 (
            .O(N__4329),
            .I(N__4312));
    InMux I__788 (
            .O(N__4328),
            .I(N__4307));
    InMux I__787 (
            .O(N__4327),
            .I(N__4307));
    InMux I__786 (
            .O(N__4326),
            .I(N__4304));
    LocalMux I__785 (
            .O(N__4323),
            .I(\U400_SDRAM.N_54 ));
    Odrv4 I__784 (
            .O(N__4320),
            .I(\U400_SDRAM.N_54 ));
    LocalMux I__783 (
            .O(N__4315),
            .I(\U400_SDRAM.N_54 ));
    LocalMux I__782 (
            .O(N__4312),
            .I(\U400_SDRAM.N_54 ));
    LocalMux I__781 (
            .O(N__4307),
            .I(\U400_SDRAM.N_54 ));
    LocalMux I__780 (
            .O(N__4304),
            .I(\U400_SDRAM.N_54 ));
    InMux I__779 (
            .O(N__4291),
            .I(N__4288));
    LocalMux I__778 (
            .O(N__4288),
            .I(\U400_SDRAM.N_276 ));
    InMux I__777 (
            .O(N__4285),
            .I(N__4282));
    LocalMux I__776 (
            .O(N__4282),
            .I(N__4279));
    Span4Mux_h I__775 (
            .O(N__4279),
            .I(N__4276));
    Span4Mux_v I__774 (
            .O(N__4276),
            .I(N__4273));
    Span4Mux_v I__773 (
            .O(N__4273),
            .I(N__4270));
    Odrv4 I__772 (
            .O(N__4270),
            .I(A_c_26));
    IoInMux I__771 (
            .O(N__4267),
            .I(N__4264));
    LocalMux I__770 (
            .O(N__4264),
            .I(N__4261));
    Odrv12 I__769 (
            .O(N__4261),
            .I(MA_c_12));
    CascadeMux I__768 (
            .O(N__4258),
            .I(N__4255));
    InMux I__767 (
            .O(N__4255),
            .I(N__4252));
    LocalMux I__766 (
            .O(N__4252),
            .I(N__4249));
    Span12Mux_v I__765 (
            .O(N__4249),
            .I(N__4246));
    Odrv12 I__764 (
            .O(N__4246),
            .I(A_c_20));
    IoInMux I__763 (
            .O(N__4243),
            .I(N__4240));
    LocalMux I__762 (
            .O(N__4240),
            .I(N__4237));
    Span4Mux_s3_v I__761 (
            .O(N__4237),
            .I(N__4234));
    Odrv4 I__760 (
            .O(N__4234),
            .I(MA_c_10));
    CascadeMux I__759 (
            .O(N__4231),
            .I(N__4228));
    InMux I__758 (
            .O(N__4228),
            .I(N__4225));
    LocalMux I__757 (
            .O(N__4225),
            .I(\U400_SDRAM.N_30_2 ));
    InMux I__756 (
            .O(N__4222),
            .I(N__4219));
    LocalMux I__755 (
            .O(N__4219),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER52_2_i_1 ));
    CascadeMux I__754 (
            .O(N__4216),
            .I(\U400_SDRAM.SDRAM_COUNTER44_5_cascade_ ));
    CascadeMux I__753 (
            .O(N__4213),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER44_0_cascade_ ));
    InMux I__752 (
            .O(N__4210),
            .I(N__4207));
    LocalMux I__751 (
            .O(N__4207),
            .I(N__4204));
    Odrv12 I__750 (
            .O(N__4204),
            .I(\U400_SDRAM.N_117 ));
    CascadeMux I__749 (
            .O(N__4201),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER52_4_i_1_cascade_ ));
    CascadeMux I__748 (
            .O(N__4198),
            .I(N__4195));
    InMux I__747 (
            .O(N__4195),
            .I(N__4192));
    LocalMux I__746 (
            .O(N__4192),
            .I(N__4189));
    Odrv12 I__745 (
            .O(N__4189),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER52_4_i_4 ));
    InMux I__744 (
            .O(N__4186),
            .I(N__4182));
    InMux I__743 (
            .O(N__4185),
            .I(N__4179));
    LocalMux I__742 (
            .O(N__4182),
            .I(\U400_SDRAM.SDRAM_COUNTER42 ));
    LocalMux I__741 (
            .O(N__4179),
            .I(\U400_SDRAM.SDRAM_COUNTER42 ));
    InMux I__740 (
            .O(N__4174),
            .I(N__4170));
    CascadeMux I__739 (
            .O(N__4173),
            .I(N__4167));
    LocalMux I__738 (
            .O(N__4170),
            .I(N__4164));
    InMux I__737 (
            .O(N__4167),
            .I(N__4161));
    Odrv4 I__736 (
            .O(N__4164),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER44_0 ));
    LocalMux I__735 (
            .O(N__4161),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER44_0 ));
    InMux I__734 (
            .O(N__4156),
            .I(N__4153));
    LocalMux I__733 (
            .O(N__4153),
            .I(\U400_SDRAM.TACK_4_m ));
    InMux I__732 (
            .O(N__4150),
            .I(N__4147));
    LocalMux I__731 (
            .O(N__4147),
            .I(N__4144));
    Odrv12 I__730 (
            .O(N__4144),
            .I(\U400_SDRAM.TACK_7_0 ));
    InMux I__729 (
            .O(N__4141),
            .I(N__4138));
    LocalMux I__728 (
            .O(N__4138),
            .I(N__4135));
    Span4Mux_h I__727 (
            .O(N__4135),
            .I(N__4130));
    InMux I__726 (
            .O(N__4134),
            .I(N__4122));
    InMux I__725 (
            .O(N__4133),
            .I(N__4122));
    Span4Mux_h I__724 (
            .O(N__4130),
            .I(N__4119));
    InMux I__723 (
            .O(N__4129),
            .I(N__4116));
    InMux I__722 (
            .O(N__4128),
            .I(N__4111));
    InMux I__721 (
            .O(N__4127),
            .I(N__4111));
    LocalMux I__720 (
            .O(N__4122),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_2 ));
    Odrv4 I__719 (
            .O(N__4119),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_2 ));
    LocalMux I__718 (
            .O(N__4116),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_2 ));
    LocalMux I__717 (
            .O(N__4111),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_2 ));
    InMux I__716 (
            .O(N__4102),
            .I(N__4099));
    LocalMux I__715 (
            .O(N__4099),
            .I(N__4096));
    Odrv12 I__714 (
            .O(N__4096),
            .I(\U400_SDRAM.TA_EN11_m ));
    InMux I__713 (
            .O(N__4093),
            .I(N__4090));
    LocalMux I__712 (
            .O(N__4090),
            .I(N__4087));
    Odrv12 I__711 (
            .O(N__4087),
            .I(\U400_SDRAM.un1_TA_COUNTER26_2_0 ));
    IoInMux I__710 (
            .O(N__4084),
            .I(N__4081));
    LocalMux I__709 (
            .O(N__4081),
            .I(N__4078));
    IoSpan4Mux I__708 (
            .O(N__4078),
            .I(N__4075));
    IoSpan4Mux I__707 (
            .O(N__4075),
            .I(N__4071));
    CascadeMux I__706 (
            .O(N__4074),
            .I(N__4068));
    Span4Mux_s3_v I__705 (
            .O(N__4071),
            .I(N__4065));
    InMux I__704 (
            .O(N__4068),
            .I(N__4062));
    Odrv4 I__703 (
            .O(N__4065),
            .I(TA_OUT));
    LocalMux I__702 (
            .O(N__4062),
            .I(TA_OUT));
    ClkMux I__701 (
            .O(N__4057),
            .I(N__3961));
    ClkMux I__700 (
            .O(N__4056),
            .I(N__3961));
    ClkMux I__699 (
            .O(N__4055),
            .I(N__3961));
    ClkMux I__698 (
            .O(N__4054),
            .I(N__3961));
    ClkMux I__697 (
            .O(N__4053),
            .I(N__3961));
    ClkMux I__696 (
            .O(N__4052),
            .I(N__3961));
    ClkMux I__695 (
            .O(N__4051),
            .I(N__3961));
    ClkMux I__694 (
            .O(N__4050),
            .I(N__3961));
    ClkMux I__693 (
            .O(N__4049),
            .I(N__3961));
    ClkMux I__692 (
            .O(N__4048),
            .I(N__3961));
    ClkMux I__691 (
            .O(N__4047),
            .I(N__3961));
    ClkMux I__690 (
            .O(N__4046),
            .I(N__3961));
    ClkMux I__689 (
            .O(N__4045),
            .I(N__3961));
    ClkMux I__688 (
            .O(N__4044),
            .I(N__3961));
    ClkMux I__687 (
            .O(N__4043),
            .I(N__3961));
    ClkMux I__686 (
            .O(N__4042),
            .I(N__3961));
    ClkMux I__685 (
            .O(N__4041),
            .I(N__3961));
    ClkMux I__684 (
            .O(N__4040),
            .I(N__3961));
    ClkMux I__683 (
            .O(N__4039),
            .I(N__3961));
    ClkMux I__682 (
            .O(N__4038),
            .I(N__3961));
    ClkMux I__681 (
            .O(N__4037),
            .I(N__3961));
    ClkMux I__680 (
            .O(N__4036),
            .I(N__3961));
    ClkMux I__679 (
            .O(N__4035),
            .I(N__3961));
    ClkMux I__678 (
            .O(N__4034),
            .I(N__3961));
    ClkMux I__677 (
            .O(N__4033),
            .I(N__3961));
    ClkMux I__676 (
            .O(N__4032),
            .I(N__3961));
    ClkMux I__675 (
            .O(N__4031),
            .I(N__3961));
    ClkMux I__674 (
            .O(N__4030),
            .I(N__3961));
    ClkMux I__673 (
            .O(N__4029),
            .I(N__3961));
    ClkMux I__672 (
            .O(N__4028),
            .I(N__3961));
    ClkMux I__671 (
            .O(N__4027),
            .I(N__3961));
    ClkMux I__670 (
            .O(N__4026),
            .I(N__3961));
    GlobalMux I__669 (
            .O(N__3961),
            .I(N__3958));
    gio2CtrlBuf I__668 (
            .O(N__3958),
            .I(CLK40_c_g));
    InMux I__667 (
            .O(N__3955),
            .I(N__3951));
    InMux I__666 (
            .O(N__3954),
            .I(N__3948));
    LocalMux I__665 (
            .O(N__3951),
            .I(N__3944));
    LocalMux I__664 (
            .O(N__3948),
            .I(N__3939));
    InMux I__663 (
            .O(N__3947),
            .I(N__3934));
    Span4Mux_v I__662 (
            .O(N__3944),
            .I(N__3931));
    InMux I__661 (
            .O(N__3943),
            .I(N__3926));
    InMux I__660 (
            .O(N__3942),
            .I(N__3926));
    Span4Mux_h I__659 (
            .O(N__3939),
            .I(N__3923));
    InMux I__658 (
            .O(N__3938),
            .I(N__3920));
    InMux I__657 (
            .O(N__3937),
            .I(N__3917));
    LocalMux I__656 (
            .O(N__3934),
            .I(\U400_SDRAM.N_105 ));
    Odrv4 I__655 (
            .O(N__3931),
            .I(\U400_SDRAM.N_105 ));
    LocalMux I__654 (
            .O(N__3926),
            .I(\U400_SDRAM.N_105 ));
    Odrv4 I__653 (
            .O(N__3923),
            .I(\U400_SDRAM.N_105 ));
    LocalMux I__652 (
            .O(N__3920),
            .I(\U400_SDRAM.N_105 ));
    LocalMux I__651 (
            .O(N__3917),
            .I(\U400_SDRAM.N_105 ));
    InMux I__650 (
            .O(N__3904),
            .I(N__3900));
    InMux I__649 (
            .O(N__3903),
            .I(N__3897));
    LocalMux I__648 (
            .O(N__3900),
            .I(N__3892));
    LocalMux I__647 (
            .O(N__3897),
            .I(N__3889));
    InMux I__646 (
            .O(N__3896),
            .I(N__3886));
    InMux I__645 (
            .O(N__3895),
            .I(N__3883));
    Odrv4 I__644 (
            .O(N__3892),
            .I(\U400_SDRAM.N_59 ));
    Odrv12 I__643 (
            .O(N__3889),
            .I(\U400_SDRAM.N_59 ));
    LocalMux I__642 (
            .O(N__3886),
            .I(\U400_SDRAM.N_59 ));
    LocalMux I__641 (
            .O(N__3883),
            .I(\U400_SDRAM.N_59 ));
    CascadeMux I__640 (
            .O(N__3874),
            .I(\U400_SDRAM.SDRAM_CMD_5_sqmuxa_cascade_ ));
    InMux I__639 (
            .O(N__3871),
            .I(N__3868));
    LocalMux I__638 (
            .O(N__3868),
            .I(\U400_SDRAM.N_84 ));
    InMux I__637 (
            .O(N__3865),
            .I(N__3861));
    InMux I__636 (
            .O(N__3864),
            .I(N__3858));
    LocalMux I__635 (
            .O(N__3861),
            .I(N__3855));
    LocalMux I__634 (
            .O(N__3858),
            .I(N__3852));
    Odrv4 I__633 (
            .O(N__3855),
            .I(\U400_SDRAM.RAM_CYCLEZ0 ));
    Odrv4 I__632 (
            .O(N__3852),
            .I(\U400_SDRAM.RAM_CYCLEZ0 ));
    CascadeMux I__631 (
            .O(N__3847),
            .I(\U400_SDRAM.N_30_2_cascade_ ));
    CascadeMux I__630 (
            .O(N__3844),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_1_0_cascade_ ));
    InMux I__629 (
            .O(N__3841),
            .I(N__3838));
    LocalMux I__628 (
            .O(N__3838),
            .I(N__3835));
    Odrv4 I__627 (
            .O(N__3835),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_3_0 ));
    InMux I__626 (
            .O(N__3832),
            .I(N__3828));
    InMux I__625 (
            .O(N__3831),
            .I(N__3825));
    LocalMux I__624 (
            .O(N__3828),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__623 (
            .O(N__3825),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__622 (
            .O(N__3820),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_4 ));
    InMux I__621 (
            .O(N__3817),
            .I(N__3813));
    InMux I__620 (
            .O(N__3816),
            .I(N__3810));
    LocalMux I__619 (
            .O(N__3813),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__618 (
            .O(N__3810),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__617 (
            .O(N__3805),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_5 ));
    InMux I__616 (
            .O(N__3802),
            .I(N__3798));
    InMux I__615 (
            .O(N__3801),
            .I(N__3795));
    LocalMux I__614 (
            .O(N__3798),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__613 (
            .O(N__3795),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__612 (
            .O(N__3790),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_6 ));
    InMux I__611 (
            .O(N__3787),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_7 ));
    SRMux I__610 (
            .O(N__3784),
            .I(N__3780));
    SRMux I__609 (
            .O(N__3783),
            .I(N__3777));
    LocalMux I__608 (
            .O(N__3780),
            .I(\U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1 ));
    LocalMux I__607 (
            .O(N__3777),
            .I(\U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1 ));
    InMux I__606 (
            .O(N__3772),
            .I(N__3769));
    LocalMux I__605 (
            .O(N__3769),
            .I(N__3766));
    Sp12to4 I__604 (
            .O(N__3766),
            .I(N__3763));
    Span12Mux_v I__603 (
            .O(N__3763),
            .I(N__3760));
    Odrv12 I__602 (
            .O(N__3760),
            .I(A_c_24));
    CascadeMux I__601 (
            .O(N__3757),
            .I(N__3754));
    InMux I__600 (
            .O(N__3754),
            .I(N__3751));
    LocalMux I__599 (
            .O(N__3751),
            .I(N__3748));
    Span4Mux_v I__598 (
            .O(N__3748),
            .I(N__3745));
    Span4Mux_h I__597 (
            .O(N__3745),
            .I(N__3742));
    Span4Mux_v I__596 (
            .O(N__3742),
            .I(N__3739));
    Odrv4 I__595 (
            .O(N__3739),
            .I(A_c_18));
    IoInMux I__594 (
            .O(N__3736),
            .I(N__3733));
    LocalMux I__593 (
            .O(N__3733),
            .I(N__3730));
    Odrv12 I__592 (
            .O(N__3730),
            .I(MA_c_8));
    CascadeMux I__591 (
            .O(N__3727),
            .I(N__3724));
    InMux I__590 (
            .O(N__3724),
            .I(N__3721));
    LocalMux I__589 (
            .O(N__3721),
            .I(N__3718));
    Sp12to4 I__588 (
            .O(N__3718),
            .I(N__3715));
    Span12Mux_s10_v I__587 (
            .O(N__3715),
            .I(N__3712));
    Odrv12 I__586 (
            .O(N__3712),
            .I(A_c_19));
    IoInMux I__585 (
            .O(N__3709),
            .I(N__3706));
    LocalMux I__584 (
            .O(N__3706),
            .I(N__3703));
    Odrv4 I__583 (
            .O(N__3703),
            .I(MA_c_9));
    InMux I__582 (
            .O(N__3700),
            .I(N__3697));
    LocalMux I__581 (
            .O(N__3697),
            .I(N__3693));
    InMux I__580 (
            .O(N__3696),
            .I(N__3690));
    Span4Mux_v I__579 (
            .O(N__3693),
            .I(N__3687));
    LocalMux I__578 (
            .O(N__3690),
            .I(N__3684));
    Odrv4 I__577 (
            .O(N__3687),
            .I(\U400_SDRAM.N_110 ));
    Odrv4 I__576 (
            .O(N__3684),
            .I(\U400_SDRAM.N_110 ));
    CascadeMux I__575 (
            .O(N__3679),
            .I(N__3676));
    InMux I__574 (
            .O(N__3676),
            .I(N__3673));
    LocalMux I__573 (
            .O(N__3673),
            .I(N__3670));
    Odrv12 I__572 (
            .O(N__3670),
            .I(RnW_c));
    CascadeMux I__571 (
            .O(N__3667),
            .I(N__3664));
    InMux I__570 (
            .O(N__3664),
            .I(N__3661));
    LocalMux I__569 (
            .O(N__3661),
            .I(\U400_SDRAM.N_57 ));
    InMux I__568 (
            .O(N__3658),
            .I(N__3652));
    InMux I__567 (
            .O(N__3657),
            .I(N__3652));
    LocalMux I__566 (
            .O(N__3652),
            .I(\U400_SDRAM.N_51 ));
    InMux I__565 (
            .O(N__3649),
            .I(N__3645));
    InMux I__564 (
            .O(N__3648),
            .I(N__3642));
    LocalMux I__563 (
            .O(N__3645),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__562 (
            .O(N__3642),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ));
    CascadeMux I__561 (
            .O(N__3637),
            .I(N__3634));
    InMux I__560 (
            .O(N__3634),
            .I(N__3629));
    InMux I__559 (
            .O(N__3633),
            .I(N__3624));
    InMux I__558 (
            .O(N__3632),
            .I(N__3624));
    LocalMux I__557 (
            .O(N__3629),
            .I(N__3621));
    LocalMux I__556 (
            .O(N__3624),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ));
    Odrv4 I__555 (
            .O(N__3621),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ));
    InMux I__554 (
            .O(N__3616),
            .I(N__3613));
    LocalMux I__553 (
            .O(N__3613),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_2 ));
    InMux I__552 (
            .O(N__3610),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_1 ));
    InMux I__551 (
            .O(N__3607),
            .I(N__3603));
    InMux I__550 (
            .O(N__3606),
            .I(N__3600));
    LocalMux I__549 (
            .O(N__3603),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__548 (
            .O(N__3600),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__547 (
            .O(N__3595),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_2 ));
    InMux I__546 (
            .O(N__3592),
            .I(N__3588));
    InMux I__545 (
            .O(N__3591),
            .I(N__3585));
    LocalMux I__544 (
            .O(N__3588),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__543 (
            .O(N__3585),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__542 (
            .O(N__3580),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_3 ));
    InMux I__541 (
            .O(N__3577),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_6 ));
    InMux I__540 (
            .O(N__3574),
            .I(N__3571));
    LocalMux I__539 (
            .O(N__3571),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_76_i_a4_1_1 ));
    InMux I__538 (
            .O(N__3568),
            .I(N__3562));
    InMux I__537 (
            .O(N__3567),
            .I(N__3562));
    LocalMux I__536 (
            .O(N__3562),
            .I(\U400_SDRAM.N_111 ));
    InMux I__535 (
            .O(N__3559),
            .I(N__3556));
    LocalMux I__534 (
            .O(N__3556),
            .I(N__3553));
    Span4Mux_v I__533 (
            .O(N__3553),
            .I(N__3550));
    Span4Mux_h I__532 (
            .O(N__3550),
            .I(N__3547));
    Odrv4 I__531 (
            .O(N__3547),
            .I(TSn_c));
    CascadeMux I__530 (
            .O(N__3544),
            .I(\U400_SDRAM.un3_RAM_CYCLE_START_cascade_ ));
    InMux I__529 (
            .O(N__3541),
            .I(N__3535));
    InMux I__528 (
            .O(N__3540),
            .I(N__3535));
    LocalMux I__527 (
            .O(N__3535),
            .I(N__3532));
    Span4Mux_h I__526 (
            .O(N__3532),
            .I(N__3523));
    InMux I__525 (
            .O(N__3531),
            .I(N__3520));
    InMux I__524 (
            .O(N__3530),
            .I(N__3517));
    InMux I__523 (
            .O(N__3529),
            .I(N__3508));
    InMux I__522 (
            .O(N__3528),
            .I(N__3508));
    InMux I__521 (
            .O(N__3527),
            .I(N__3508));
    InMux I__520 (
            .O(N__3526),
            .I(N__3508));
    Odrv4 I__519 (
            .O(N__3523),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    LocalMux I__518 (
            .O(N__3520),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    LocalMux I__517 (
            .O(N__3517),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    LocalMux I__516 (
            .O(N__3508),
            .I(\U400_SDRAM.RAM_CYCLE_STARTZ0 ));
    InMux I__515 (
            .O(N__3499),
            .I(N__3494));
    InMux I__514 (
            .O(N__3498),
            .I(N__3491));
    InMux I__513 (
            .O(N__3497),
            .I(N__3488));
    LocalMux I__512 (
            .O(N__3494),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__511 (
            .O(N__3491),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__510 (
            .O(N__3488),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__509 (
            .O(N__3481),
            .I(N__3476));
    InMux I__508 (
            .O(N__3480),
            .I(N__3471));
    InMux I__507 (
            .O(N__3479),
            .I(N__3471));
    LocalMux I__506 (
            .O(N__3476),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__505 (
            .O(N__3471),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__504 (
            .O(N__3466),
            .I(N__3461));
    InMux I__503 (
            .O(N__3465),
            .I(N__3458));
    InMux I__502 (
            .O(N__3464),
            .I(N__3455));
    InMux I__501 (
            .O(N__3461),
            .I(N__3452));
    LocalMux I__500 (
            .O(N__3458),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__499 (
            .O(N__3455),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__498 (
            .O(N__3452),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__497 (
            .O(N__3445),
            .I(N__3440));
    InMux I__496 (
            .O(N__3444),
            .I(N__3435));
    InMux I__495 (
            .O(N__3443),
            .I(N__3435));
    LocalMux I__494 (
            .O(N__3440),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__493 (
            .O(N__3435),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ));
    CascadeMux I__492 (
            .O(N__3430),
            .I(\U400_SDRAM.N_54_cascade_ ));
    InMux I__491 (
            .O(N__3427),
            .I(N__3424));
    LocalMux I__490 (
            .O(N__3424),
            .I(N__3421));
    Span12Mux_s11_h I__489 (
            .O(N__3421),
            .I(N__3418));
    Odrv12 I__488 (
            .O(N__3418),
            .I(A_c_9));
    CascadeMux I__487 (
            .O(N__3415),
            .I(N__3412));
    InMux I__486 (
            .O(N__3412),
            .I(N__3409));
    LocalMux I__485 (
            .O(N__3409),
            .I(N__3406));
    Span4Mux_v I__484 (
            .O(N__3406),
            .I(N__3403));
    Odrv4 I__483 (
            .O(N__3403),
            .I(A_c_17));
    IoInMux I__482 (
            .O(N__3400),
            .I(N__3397));
    LocalMux I__481 (
            .O(N__3397),
            .I(N__3394));
    Odrv12 I__480 (
            .O(N__3394),
            .I(MA_c_7));
    InMux I__479 (
            .O(N__3391),
            .I(N__3388));
    LocalMux I__478 (
            .O(N__3388),
            .I(N__3385));
    Odrv12 I__477 (
            .O(N__3385),
            .I(A_c_8));
    CascadeMux I__476 (
            .O(N__3382),
            .I(N__3379));
    InMux I__475 (
            .O(N__3379),
            .I(N__3376));
    LocalMux I__474 (
            .O(N__3376),
            .I(N__3373));
    Span4Mux_v I__473 (
            .O(N__3373),
            .I(N__3370));
    Span4Mux_v I__472 (
            .O(N__3370),
            .I(N__3367));
    Odrv4 I__471 (
            .O(N__3367),
            .I(A_c_16));
    IoInMux I__470 (
            .O(N__3364),
            .I(N__3361));
    LocalMux I__469 (
            .O(N__3361),
            .I(N__3358));
    Odrv12 I__468 (
            .O(N__3358),
            .I(MA_c_6));
    InMux I__467 (
            .O(N__3355),
            .I(bfn_5_4_0_));
    InMux I__466 (
            .O(N__3352),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_0 ));
    InMux I__465 (
            .O(N__3349),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_1 ));
    InMux I__464 (
            .O(N__3346),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_2 ));
    InMux I__463 (
            .O(N__3343),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_3 ));
    InMux I__462 (
            .O(N__3340),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_4 ));
    InMux I__461 (
            .O(N__3337),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_5 ));
    CascadeMux I__460 (
            .O(N__3334),
            .I(\U400_SDRAM.N_57_cascade_ ));
    InMux I__459 (
            .O(N__3331),
            .I(N__3325));
    InMux I__458 (
            .O(N__3330),
            .I(N__3325));
    LocalMux I__457 (
            .O(N__3325),
            .I(\U400_SDRAM.N_46 ));
    CascadeMux I__456 (
            .O(N__3322),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_o5_0_cascade_ ));
    CascadeMux I__455 (
            .O(N__3319),
            .I(\U400_SDRAM.N_266_0_cascade_ ));
    InMux I__454 (
            .O(N__3316),
            .I(N__3312));
    InMux I__453 (
            .O(N__3315),
            .I(N__3309));
    LocalMux I__452 (
            .O(N__3312),
            .I(N__3303));
    LocalMux I__451 (
            .O(N__3309),
            .I(N__3303));
    InMux I__450 (
            .O(N__3308),
            .I(N__3300));
    Odrv12 I__449 (
            .O(N__3303),
            .I(\U400_SDRAM.SDRAM_CMD12 ));
    LocalMux I__448 (
            .O(N__3300),
            .I(\U400_SDRAM.SDRAM_CMD12 ));
    CascadeMux I__447 (
            .O(N__3295),
            .I(\U400_SDRAM.SDRAM_CMD12_cascade_ ));
    CascadeMux I__446 (
            .O(N__3292),
            .I(N__3289));
    InMux I__445 (
            .O(N__3289),
            .I(N__3283));
    InMux I__444 (
            .O(N__3288),
            .I(N__3283));
    LocalMux I__443 (
            .O(N__3283),
            .I(N__3280));
    Odrv4 I__442 (
            .O(N__3280),
            .I(\U400_SDRAM.un1_SDRAM_COUNTER52_0 ));
    InMux I__441 (
            .O(N__3277),
            .I(N__3273));
    InMux I__440 (
            .O(N__3276),
            .I(N__3270));
    LocalMux I__439 (
            .O(N__3273),
            .I(N__3267));
    LocalMux I__438 (
            .O(N__3270),
            .I(\U400_SDRAM.CS0_ENZ0 ));
    Odrv12 I__437 (
            .O(N__3267),
            .I(\U400_SDRAM.CS0_ENZ0 ));
    IoInMux I__436 (
            .O(N__3262),
            .I(N__3259));
    LocalMux I__435 (
            .O(N__3259),
            .I(N__3256));
    IoSpan4Mux I__434 (
            .O(N__3256),
            .I(N__3253));
    Span4Mux_s3_h I__433 (
            .O(N__3253),
            .I(N__3250));
    Odrv4 I__432 (
            .O(N__3250),
            .I(CS0n_c));
    IoInMux I__431 (
            .O(N__3247),
            .I(N__3244));
    LocalMux I__430 (
            .O(N__3244),
            .I(N__3241));
    Odrv12 I__429 (
            .O(N__3241),
            .I(WEn_c));
    IoInMux I__428 (
            .O(N__3238),
            .I(N__3235));
    LocalMux I__427 (
            .O(N__3235),
            .I(N__3232));
    Odrv12 I__426 (
            .O(N__3232),
            .I(CASn_c));
    CascadeMux I__425 (
            .O(N__3229),
            .I(N__3226));
    InMux I__424 (
            .O(N__3226),
            .I(N__3222));
    InMux I__423 (
            .O(N__3225),
            .I(N__3219));
    LocalMux I__422 (
            .O(N__3222),
            .I(N__3216));
    LocalMux I__421 (
            .O(N__3219),
            .I(\U400_SDRAM.CS1_ENZ0 ));
    Odrv12 I__420 (
            .O(N__3216),
            .I(\U400_SDRAM.CS1_ENZ0 ));
    IoInMux I__419 (
            .O(N__3211),
            .I(N__3208));
    LocalMux I__418 (
            .O(N__3208),
            .I(N__3205));
    IoSpan4Mux I__417 (
            .O(N__3205),
            .I(N__3202));
    Span4Mux_s3_v I__416 (
            .O(N__3202),
            .I(N__3199));
    Odrv4 I__415 (
            .O(N__3199),
            .I(CS1n_c));
    CascadeMux I__414 (
            .O(N__3196),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_3_0_cascade_ ));
    CascadeMux I__413 (
            .O(N__3193),
            .I(\U400_SDRAM.N_55_cascade_ ));
    CascadeMux I__412 (
            .O(N__3190),
            .I(\U400_SDRAM.N_105_cascade_ ));
    InMux I__411 (
            .O(N__3187),
            .I(N__3183));
    InMux I__410 (
            .O(N__3186),
            .I(N__3180));
    LocalMux I__409 (
            .O(N__3183),
            .I(\U400_SDRAM.N_68 ));
    LocalMux I__408 (
            .O(N__3180),
            .I(\U400_SDRAM.N_68 ));
    CascadeMux I__407 (
            .O(N__3175),
            .I(\U400_SDRAM.N_62_cascade_ ));
    CascadeMux I__406 (
            .O(N__3172),
            .I(\U400_SDRAM.N_39_cascade_ ));
    InMux I__405 (
            .O(N__3169),
            .I(N__3166));
    LocalMux I__404 (
            .O(N__3166),
            .I(\U400_SDRAM.N_62 ));
    CascadeMux I__403 (
            .O(N__3163),
            .I(N__3160));
    InMux I__402 (
            .O(N__3160),
            .I(N__3154));
    InMux I__401 (
            .O(N__3159),
            .I(N__3154));
    LocalMux I__400 (
            .O(N__3154),
            .I(N__3151));
    Span4Mux_h I__399 (
            .O(N__3151),
            .I(N__3148));
    Span4Mux_v I__398 (
            .O(N__3148),
            .I(N__3145));
    Odrv4 I__397 (
            .O(N__3145),
            .I(A_c_23));
    CascadeMux I__396 (
            .O(N__3142),
            .I(\U400_SDRAM.N_41_cascade_ ));
    InMux I__395 (
            .O(N__3139),
            .I(N__3136));
    LocalMux I__394 (
            .O(N__3136),
            .I(\U400_SDRAM.N_52 ));
    CascadeMux I__393 (
            .O(N__3133),
            .I(\U400_SDRAM.N_295_0_cascade_ ));
    CascadeMux I__392 (
            .O(N__3130),
            .I(\U400_SDRAM.N_300_cascade_ ));
    InMux I__391 (
            .O(N__3127),
            .I(N__3124));
    LocalMux I__390 (
            .O(N__3124),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_0_76_i_0 ));
    CascadeMux I__389 (
            .O(N__3121),
            .I(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_2_0_cascade_ ));
    CascadeMux I__388 (
            .O(N__3118),
            .I(\U400_SDRAM.N_110_cascade_ ));
    CascadeMux I__387 (
            .O(N__3115),
            .I(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_a4_1_0_cascade_ ));
    InMux I__386 (
            .O(N__3112),
            .I(N__3107));
    InMux I__385 (
            .O(N__3111),
            .I(N__3102));
    InMux I__384 (
            .O(N__3110),
            .I(N__3102));
    LocalMux I__383 (
            .O(N__3107),
            .I(\U400_SDRAM.BURSTZ0 ));
    LocalMux I__382 (
            .O(N__3102),
            .I(\U400_SDRAM.BURSTZ0 ));
    InMux I__381 (
            .O(N__3097),
            .I(N__3088));
    InMux I__380 (
            .O(N__3096),
            .I(N__3088));
    InMux I__379 (
            .O(N__3095),
            .I(N__3084));
    InMux I__378 (
            .O(N__3094),
            .I(N__3081));
    InMux I__377 (
            .O(N__3093),
            .I(N__3078));
    LocalMux I__376 (
            .O(N__3088),
            .I(N__3075));
    InMux I__375 (
            .O(N__3087),
            .I(N__3072));
    LocalMux I__374 (
            .O(N__3084),
            .I(\U400_SDRAM.TACKZ0 ));
    LocalMux I__373 (
            .O(N__3081),
            .I(\U400_SDRAM.TACKZ0 ));
    LocalMux I__372 (
            .O(N__3078),
            .I(\U400_SDRAM.TACKZ0 ));
    Odrv4 I__371 (
            .O(N__3075),
            .I(\U400_SDRAM.TACKZ0 ));
    LocalMux I__370 (
            .O(N__3072),
            .I(\U400_SDRAM.TACKZ0 ));
    InMux I__369 (
            .O(N__3061),
            .I(N__3058));
    LocalMux I__368 (
            .O(N__3058),
            .I(N__3055));
    Span4Mux_v I__367 (
            .O(N__3055),
            .I(N__3052));
    Odrv4 I__366 (
            .O(N__3052),
            .I(A_c_22));
    IoInMux I__365 (
            .O(N__3049),
            .I(N__3046));
    LocalMux I__364 (
            .O(N__3046),
            .I(N__3043));
    IoSpan4Mux I__363 (
            .O(N__3043),
            .I(N__3040));
    Span4Mux_s1_h I__362 (
            .O(N__3040),
            .I(N__3036));
    InMux I__361 (
            .O(N__3039),
            .I(N__3033));
    Odrv4 I__360 (
            .O(N__3036),
            .I(BANK1_c));
    LocalMux I__359 (
            .O(N__3033),
            .I(BANK1_c));
    CascadeMux I__358 (
            .O(N__3028),
            .I(N__3025));
    InMux I__357 (
            .O(N__3025),
            .I(N__3022));
    LocalMux I__356 (
            .O(N__3022),
            .I(N__3019));
    Span4Mux_v I__355 (
            .O(N__3019),
            .I(N__3016));
    Odrv4 I__354 (
            .O(N__3016),
            .I(A_c_21));
    IoInMux I__353 (
            .O(N__3013),
            .I(N__3010));
    LocalMux I__352 (
            .O(N__3010),
            .I(N__3007));
    Span12Mux_s1_h I__351 (
            .O(N__3007),
            .I(N__3003));
    InMux I__350 (
            .O(N__3006),
            .I(N__3000));
    Odrv12 I__349 (
            .O(N__3003),
            .I(BANK0_c));
    LocalMux I__348 (
            .O(N__3000),
            .I(BANK0_c));
    IoInMux I__347 (
            .O(N__2995),
            .I(N__2992));
    LocalMux I__346 (
            .O(N__2992),
            .I(N__2989));
    Odrv4 I__345 (
            .O(N__2989),
            .I(RASn_c));
    CascadeMux I__344 (
            .O(N__2986),
            .I(\U400_SDRAM.N_299_cascade_ ));
    CascadeMux I__343 (
            .O(N__2983),
            .I(\U400_SDRAM.un1_TA_COUNTER26_0_cascade_ ));
    CascadeMux I__342 (
            .O(N__2980),
            .I(\U400_SDRAM.TA_COUNTER23_cascade_ ));
    CascadeMux I__341 (
            .O(N__2977),
            .I(\U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_ ));
    InMux I__340 (
            .O(N__2974),
            .I(N__2966));
    InMux I__339 (
            .O(N__2973),
            .I(N__2963));
    InMux I__338 (
            .O(N__2972),
            .I(N__2960));
    InMux I__337 (
            .O(N__2971),
            .I(N__2953));
    InMux I__336 (
            .O(N__2970),
            .I(N__2953));
    InMux I__335 (
            .O(N__2969),
            .I(N__2953));
    LocalMux I__334 (
            .O(N__2966),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_1 ));
    LocalMux I__333 (
            .O(N__2963),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_1 ));
    LocalMux I__332 (
            .O(N__2960),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_1 ));
    LocalMux I__331 (
            .O(N__2953),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_1 ));
    InMux I__330 (
            .O(N__2944),
            .I(N__2932));
    InMux I__329 (
            .O(N__2943),
            .I(N__2932));
    InMux I__328 (
            .O(N__2942),
            .I(N__2929));
    InMux I__327 (
            .O(N__2941),
            .I(N__2918));
    InMux I__326 (
            .O(N__2940),
            .I(N__2918));
    InMux I__325 (
            .O(N__2939),
            .I(N__2918));
    InMux I__324 (
            .O(N__2938),
            .I(N__2918));
    InMux I__323 (
            .O(N__2937),
            .I(N__2918));
    LocalMux I__322 (
            .O(N__2932),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_0 ));
    LocalMux I__321 (
            .O(N__2929),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_0 ));
    LocalMux I__320 (
            .O(N__2918),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_0 ));
    CascadeMux I__319 (
            .O(N__2911),
            .I(N__2905));
    CascadeMux I__318 (
            .O(N__2910),
            .I(N__2901));
    CascadeMux I__317 (
            .O(N__2909),
            .I(N__2898));
    CascadeMux I__316 (
            .O(N__2908),
            .I(N__2895));
    InMux I__315 (
            .O(N__2905),
            .I(N__2892));
    InMux I__314 (
            .O(N__2904),
            .I(N__2889));
    InMux I__313 (
            .O(N__2901),
            .I(N__2886));
    InMux I__312 (
            .O(N__2898),
            .I(N__2881));
    InMux I__311 (
            .O(N__2895),
            .I(N__2881));
    LocalMux I__310 (
            .O(N__2892),
            .I(N__2878));
    LocalMux I__309 (
            .O(N__2889),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_3 ));
    LocalMux I__308 (
            .O(N__2886),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_3 ));
    LocalMux I__307 (
            .O(N__2881),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_3 ));
    Odrv4 I__306 (
            .O(N__2878),
            .I(\U400_SDRAM.TA_COUNTERZ0Z_3 ));
    InMux I__305 (
            .O(N__2869),
            .I(N__2865));
    InMux I__304 (
            .O(N__2868),
            .I(N__2862));
    LocalMux I__303 (
            .O(N__2865),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa ));
    LocalMux I__302 (
            .O(N__2862),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa ));
    InMux I__301 (
            .O(N__2857),
            .I(N__2853));
    CascadeMux I__300 (
            .O(N__2856),
            .I(N__2850));
    LocalMux I__299 (
            .O(N__2853),
            .I(N__2845));
    InMux I__298 (
            .O(N__2850),
            .I(N__2842));
    InMux I__297 (
            .O(N__2849),
            .I(N__2839));
    InMux I__296 (
            .O(N__2848),
            .I(N__2836));
    Odrv4 I__295 (
            .O(N__2845),
            .I(\U400_SDRAM.TA_COUNTER23 ));
    LocalMux I__294 (
            .O(N__2842),
            .I(\U400_SDRAM.TA_COUNTER23 ));
    LocalMux I__293 (
            .O(N__2839),
            .I(\U400_SDRAM.TA_COUNTER23 ));
    LocalMux I__292 (
            .O(N__2836),
            .I(\U400_SDRAM.TA_COUNTER23 ));
    InMux I__291 (
            .O(N__2827),
            .I(N__2823));
    InMux I__290 (
            .O(N__2826),
            .I(N__2820));
    LocalMux I__289 (
            .O(N__2823),
            .I(\U400_SDRAM.TA_COUNTER27 ));
    LocalMux I__288 (
            .O(N__2820),
            .I(\U400_SDRAM.TA_COUNTER27 ));
    CascadeMux I__287 (
            .O(N__2815),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_ ));
    InMux I__286 (
            .O(N__2812),
            .I(N__2809));
    LocalMux I__285 (
            .O(N__2809),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en ));
    InMux I__284 (
            .O(N__2806),
            .I(N__2803));
    LocalMux I__283 (
            .O(N__2803),
            .I(\U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0 ));
    CascadeMux I__282 (
            .O(N__2800),
            .I(N__2797));
    InMux I__281 (
            .O(N__2797),
            .I(N__2791));
    InMux I__280 (
            .O(N__2796),
            .I(N__2791));
    LocalMux I__279 (
            .O(N__2791),
            .I(\U400_SDRAM.CO1 ));
    CascadeMux I__278 (
            .O(N__2788),
            .I(\U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_ ));
    CEMux I__277 (
            .O(N__2785),
            .I(N__2782));
    LocalMux I__276 (
            .O(N__2782),
            .I(N__2779));
    Span4Mux_s1_h I__275 (
            .O(N__2779),
            .I(N__2776));
    Odrv4 I__274 (
            .O(N__2776),
            .I(\U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0 ));
    IoInMux I__273 (
            .O(N__2773),
            .I(N__2770));
    LocalMux I__272 (
            .O(N__2770),
            .I(RESETn_c_i));
    IoInMux I__271 (
            .O(N__2767),
            .I(N__2764));
    LocalMux I__270 (
            .O(N__2764),
            .I(CONSTANT_ONE_NET));
    InMux I__269 (
            .O(N__2761),
            .I(N__2758));
    LocalMux I__268 (
            .O(N__2758),
            .I(N__2755));
    Odrv4 I__267 (
            .O(N__2755),
            .I(A_c_31));
    CascadeMux I__266 (
            .O(N__2752),
            .I(N__2749));
    InMux I__265 (
            .O(N__2749),
            .I(N__2746));
    LocalMux I__264 (
            .O(N__2746),
            .I(N__2743));
    Span4Mux_h I__263 (
            .O(N__2743),
            .I(N__2740));
    Odrv4 I__262 (
            .O(N__2740),
            .I(A_c_30));
    InMux I__261 (
            .O(N__2737),
            .I(N__2734));
    LocalMux I__260 (
            .O(N__2734),
            .I(N__2731));
    Odrv12 I__259 (
            .O(N__2731),
            .I(A_c_27));
    IoInMux I__258 (
            .O(N__2728),
            .I(N__2725));
    LocalMux I__257 (
            .O(N__2725),
            .I(N__2722));
    IoSpan4Mux I__256 (
            .O(N__2722),
            .I(N__2719));
    Span4Mux_s3_h I__255 (
            .O(N__2719),
            .I(N__2716));
    Span4Mux_h I__254 (
            .O(N__2716),
            .I(N__2713));
    Span4Mux_h I__253 (
            .O(N__2713),
            .I(N__2710));
    Span4Mux_v I__252 (
            .O(N__2710),
            .I(N__2707));
    Odrv4 I__251 (
            .O(N__2707),
            .I(CLK40_ibuf_gb_io_gb_input));
    INV \INVU400_SDRAM.MA_nesr_4C  (
            .O(\INVU400_SDRAM.MA_nesr_4C_net ),
            .I(N__4057));
    INV \INVU400_SDRAM.MA_nesr_3C  (
            .O(\INVU400_SDRAM.MA_nesr_3C_net ),
            .I(N__4055));
    INV \INVU400_SDRAM.MA_nesr_5C  (
            .O(\INVU400_SDRAM.MA_nesr_5C_net ),
            .I(N__4056));
    INV \INVU400_SDRAM.MA_nesr_11C  (
            .O(\INVU400_SDRAM.MA_nesr_11C_net ),
            .I(N__4052));
    INV \INVU400_SDRAM.SDRAM_CMD_1C  (
            .O(\INVU400_SDRAM.SDRAM_CMD_1C_net ),
            .I(N__4045));
    INV \INVU400_SDRAM.SDRAM_CONFIGUREDC  (
            .O(\INVU400_SDRAM.SDRAM_CONFIGUREDC_net ),
            .I(N__4050));
    INV \INVU400_SDRAM.SDRAM_COUNTER_0C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_0C_net ),
            .I(N__4053));
    INV \INVU400_SDRAM.MA_nesr_10C  (
            .O(\INVU400_SDRAM.MA_nesr_10C_net ),
            .I(N__4048));
    INV \INVU400_SDRAM.MA_nesr_12C  (
            .O(\INVU400_SDRAM.MA_nesr_12C_net ),
            .I(N__4044));
    INV \INVU400_SDRAM.RAM_CYCLEC  (
            .O(\INVU400_SDRAM.RAM_CYCLEC_net ),
            .I(N__4049));
    INV \INVU400_SDRAM.WRITE_CYCLEC  (
            .O(\INVU400_SDRAM.WRITE_CYCLEC_net ),
            .I(N__4054));
    INV \INVU400_SDRAM.MA_nesr_9C  (
            .O(\INVU400_SDRAM.MA_nesr_9C_net ),
            .I(N__4046));
    INV \INVU400_SDRAM.MA_nesr_8C  (
            .O(\INVU400_SDRAM.MA_nesr_8C_net ),
            .I(N__4039));
    INV \INVU400_SDRAM.REFRESH_COUNTER_2C  (
            .O(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .I(N__4037));
    INV \INVU400_SDRAM.REFRESH_COUNTER_0C  (
            .O(\INVU400_SDRAM.REFRESH_COUNTER_0C_net ),
            .I(N__4040));
    INV \INVU400_SDRAM.SDRAM_COUNTER_2C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .I(N__4047));
    INV \INVU400_SDRAM.MA_nesr_6C  (
            .O(\INVU400_SDRAM.MA_nesr_6C_net ),
            .I(N__4041));
    INV \INVU400_SDRAM.MA_nesr_7C  (
            .O(\INVU400_SDRAM.MA_nesr_7C_net ),
            .I(N__4035));
    INV \INVU400_SDRAM.CS1nC  (
            .O(\INVU400_SDRAM.CS1nC_net ),
            .I(N__4032));
    INV \INVU400_SDRAM.CS0nC  (
            .O(\INVU400_SDRAM.CS0nC_net ),
            .I(N__4027));
    INV \INVU400_SDRAM.CS0_ENC  (
            .O(\INVU400_SDRAM.CS0_ENC_net ),
            .I(N__4036));
    INV \INVU400_SDRAM.SDRAM_CMD_0C  (
            .O(\INVU400_SDRAM.SDRAM_CMD_0C_net ),
            .I(N__4038));
    INV \INVU400_SDRAM.SDRAM_CMD_2C  (
            .O(\INVU400_SDRAM.SDRAM_CMD_2C_net ),
            .I(N__4042));
    INV \INVU400_SDRAM.RASnC  (
            .O(\INVU400_SDRAM.RASnC_net ),
            .I(N__4026));
    INV \INVU400_SDRAM.BANK1C  (
            .O(\INVU400_SDRAM.BANK1C_net ),
            .I(N__4029));
    INV \INVU400_SDRAM.TACKC  (
            .O(\INVU400_SDRAM.TACKC_net ),
            .I(N__4031));
    INV \INVU400_SDRAM.BURSTC  (
            .O(\INVU400_SDRAM.BURSTC_net ),
            .I(N__4033));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_5_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_4_0_));
    ICE_GB CLK40_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__2728),
            .GLOBALBUFFEROUTPUT(CLK40_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__2773),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_1_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_1_5_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_1_5_1  (
            .in0(_gnd_net_),
            .in1(N__6513),
            .in2(_gnd_net_),
            .in3(N__2812),
            .lcout(\U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_1_LC_1_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_1_LC_1_5_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_1_LC_1_5_2 .LUT_INIT=16'b0110000000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_1_LC_1_5_2  (
            .in0(N__2974),
            .in1(N__2944),
            .in2(N__5236),
            .in3(N__2806),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4030),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_3_LC_1_5_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_3_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_3_LC_1_5_3 .LUT_INIT=16'b0100110010000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_3_LC_1_5_3  (
            .in0(N__4134),
            .in1(N__5234),
            .in2(N__2800),
            .in3(N__2904),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4030),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_1_5_4 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_1_5_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(N__2973),
            .in2(_gnd_net_),
            .in3(N__2943),
            .lcout(\U400_SDRAM.CO1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNI0LUG4_LC_1_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNI0LUG4_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNI0LUG4_LC_1_5_5 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \U400_SDRAM.TACK_RNI0LUG4_LC_1_5_5  (
            .in0(N__3093),
            .in1(N__2827),
            .in2(N__2856),
            .in3(N__2868),
            .lcout(\U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0 ),
            .ltout(\U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_2_LC_1_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_2_LC_1_5_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_2_LC_1_5_6 .LUT_INIT=16'b0010000010000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_2_LC_1_5_6  (
            .in0(N__5233),
            .in1(N__2796),
            .in2(N__2788),
            .in3(N__4133),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4030),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_EN_i_ess_LC_1_6_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_EN_i_ess_LC_1_6_3 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.TA_EN_i_ess_LC_1_6_3 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U400_SDRAM.TA_EN_i_ess_LC_1_6_3  (
            .in0(N__2857),
            .in1(N__5227),
            .in2(_gnd_net_),
            .in3(N__3094),
            .lcout(TA_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4028),
            .ce(N__2785),
            .sr(N__6479));
    defparam RESETn_ibuf_RNIM9SF_LC_1_8_3.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_1_8_3.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_1_8_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_1_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5213),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_1_14_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_14_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_14_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_3_LC_2_2_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_3_LC_2_2_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_3_LC_2_2_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U400_ADDRESS_DECODE.RAM_SPACE_3_LC_2_2_2  (
            .in0(N__5235),
            .in1(N__2761),
            .in2(N__2752),
            .in3(N__2737),
            .lcout(U400_ADDRESS_DECODE_RAM_SPACE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_2_4_0 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_2_4_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_2_4_0  (
            .in0(N__2969),
            .in1(N__4127),
            .in2(N__2908),
            .in3(N__2937),
            .lcout(\U400_SDRAM.TA_COUNTER27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_OUT_RNO_2_LC_2_4_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_RNO_2_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_OUT_RNO_2_LC_2_4_2 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \U400_SDRAM.TA_OUT_RNO_2_LC_2_4_2  (
            .in0(N__2971),
            .in1(N__4128),
            .in2(N__2909),
            .in3(N__2939),
            .lcout(),
            .ltout(\U400_SDRAM.un1_TA_COUNTER26_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_OUT_RNO_1_LC_2_4_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_RNO_1_LC_2_4_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_OUT_RNO_1_LC_2_4_3 .LUT_INIT=16'b0000101000001111;
    LogicCell40 \U400_SDRAM.TA_OUT_RNO_1_LC_2_4_3  (
            .in0(N__3097),
            .in1(_gnd_net_),
            .in2(N__2983),
            .in3(N__2849),
            .lcout(\U400_SDRAM.un1_TA_COUNTER26_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_OUT_RNO_0_LC_2_4_4 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_RNO_0_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_OUT_RNO_0_LC_2_4_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U400_SDRAM.TA_OUT_RNO_0_LC_2_4_4  (
            .in0(_gnd_net_),
            .in1(N__2940),
            .in2(_gnd_net_),
            .in3(N__3112),
            .lcout(\U400_SDRAM.TA_EN11_m ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_2_4_5 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_2_4_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_2_4_5  (
            .in0(N__2938),
            .in1(N__4129),
            .in2(N__2910),
            .in3(N__2970),
            .lcout(\U400_SDRAM.TA_COUNTER23 ),
            .ltout(\U400_SDRAM.TA_COUNTER23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_2_4_6 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_2_4_6 .LUT_INIT=16'b0000110000111100;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_2_4_6  (
            .in0(_gnd_net_),
            .in1(N__2941),
            .in2(N__2980),
            .in3(N__3096),
            .lcout(),
            .ltout(\U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_0_LC_2_4_7 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_0_LC_2_4_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_0_LC_2_4_7 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_0_LC_2_4_7  (
            .in0(_gnd_net_),
            .in1(N__2869),
            .in2(N__2977),
            .in3(N__5229),
            .lcout(\U400_SDRAM.TA_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4034),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.BURST_RNISKH51_LC_2_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.BURST_RNISKH51_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.BURST_RNISKH51_LC_2_5_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U400_SDRAM.BURST_RNISKH51_LC_2_5_0  (
            .in0(N__2972),
            .in1(N__2942),
            .in2(N__2911),
            .in3(N__3110),
            .lcout(\U400_SDRAM.TA_COUNTER_0_sqmuxa ),
            .ltout(\U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_2_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_2_5_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_2_5_1  (
            .in0(N__2848),
            .in1(N__2826),
            .in2(N__2815),
            .in3(N__3087),
            .lcout(\U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.BURST_LC_2_5_3 .C_ON=1'b0;
    defparam \U400_SDRAM.BURST_LC_2_5_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BURST_LC_2_5_3 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \U400_SDRAM.BURST_LC_2_5_3  (
            .in0(N__3111),
            .in1(N__3696),
            .in2(N__6352),
            .in3(N__3903),
            .lcout(\U400_SDRAM.BURSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BURSTC_net ),
            .ce(),
            .sr(N__6486));
    defparam \U400_SDRAM.TACK_LC_2_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_LC_2_6_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TACK_LC_2_6_1 .LUT_INIT=16'b1111101100000001;
    LogicCell40 \U400_SDRAM.TACK_LC_2_6_1  (
            .in0(N__4210),
            .in1(N__4150),
            .in2(N__4198),
            .in3(N__3095),
            .lcout(\U400_SDRAM.TACKZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.TACKC_net ),
            .ce(),
            .sr(N__6482));
    defparam \U400_SDRAM.BANK1_LC_2_7_2 .C_ON=1'b0;
    defparam \U400_SDRAM.BANK1_LC_2_7_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BANK1_LC_2_7_2 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \U400_SDRAM.BANK1_LC_2_7_2  (
            .in0(N__3541),
            .in1(N__3061),
            .in2(N__3292),
            .in3(N__3039),
            .lcout(BANK1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK1C_net ),
            .ce(),
            .sr(N__6480));
    defparam \U400_SDRAM.BANK0_LC_2_7_5 .C_ON=1'b0;
    defparam \U400_SDRAM.BANK0_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BANK0_LC_2_7_5 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \U400_SDRAM.BANK0_LC_2_7_5  (
            .in0(N__3006),
            .in1(N__3288),
            .in2(N__3028),
            .in3(N__3540),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK1C_net ),
            .ce(),
            .sr(N__6480));
    defparam \U400_SDRAM.RASn_LC_2_10_1 .C_ON=1'b0;
    defparam \U400_SDRAM.RASn_LC_2_10_1 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.RASn_LC_2_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.RASn_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6835),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.RASnC_net ),
            .ce(),
            .sr(N__6481));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_4_4_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_4_4_1 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_4_4_1  (
            .in0(N__4402),
            .in1(N__3315),
            .in2(N__4579),
            .in3(N__3530),
            .lcout(),
            .ltout(\U400_SDRAM.N_299_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_4_4_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_4_4_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_4_4_2 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_2_LC_4_4_2  (
            .in0(N__6753),
            .in1(N__3127),
            .in2(N__2986),
            .in3(N__5904),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_2_LC_4_4_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_2_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_2_LC_4_4_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_4_2_LC_4_4_3  (
            .in0(N__3464),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3498),
            .lcout(\U400_SDRAM.N_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_5_2_LC_4_4_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_5_2_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_5_2_LC_4_4_5 .LUT_INIT=16'b1111111011011010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_5_2_LC_4_4_5  (
            .in0(N__5068),
            .in1(N__4977),
            .in2(N__4866),
            .in3(N__4714),
            .lcout(),
            .ltout(\U400_SDRAM.N_295_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_4_4_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_4_4_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_4_4_6  (
            .in0(N__3574),
            .in1(N__3139),
            .in2(N__3133),
            .in3(N__5336),
            .lcout(),
            .ltout(\U400_SDRAM.N_300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_4_4_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_4_4_7 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_4_4_7  (
            .in0(N__5337),
            .in1(N__5074),
            .in2(N__3130),
            .in3(N__4510),
            .lcout(\U400_SDRAM.SDRAM_CMD_cnst_0_76_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_2_LC_4_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_2_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_2_LC_4_5_0 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_2_LC_4_5_0  (
            .in0(N__4846),
            .in1(N__5040),
            .in2(_gnd_net_),
            .in3(N__4327),
            .lcout(\U400_SDRAM.N_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_4_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_4_5_1 .LUT_INIT=16'b0010000011111110;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_4_5_1  (
            .in0(N__4973),
            .in1(N__5430),
            .in2(N__4864),
            .in3(N__5335),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_0_LC_4_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_0_LC_4_5_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_0_LC_4_5_2 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_0_LC_4_5_2  (
            .in0(N__6122),
            .in1(N__5903),
            .in2(N__3121),
            .in3(N__3841),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITAGQ1_1_LC_4_5_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITAGQ1_1_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITAGQ1_1_LC_4_5_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNITAGQ1_1_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(N__4693),
            .in2(_gnd_net_),
            .in3(N__3938),
            .lcout(\U400_SDRAM.N_110 ),
            .ltout(\U400_SDRAM.N_110_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIFGBJ4_LC_4_5_4 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIFGBJ4_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNIFGBJ4_LC_4_5_4 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNIFGBJ4_LC_4_5_4  (
            .in0(N__5209),
            .in1(N__3316),
            .in2(N__3118),
            .in3(N__3531),
            .lcout(\U400_SDRAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI5LLK_3_LC_4_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI5LLK_3_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI5LLK_3_LC_4_5_5 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI5LLK_3_LC_4_5_5  (
            .in0(N__4972),
            .in1(N__4847),
            .in2(_gnd_net_),
            .in3(N__4692),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_a4_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITM402_3_LC_4_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITM402_3_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNITM402_3_LC_4_5_6 .LUT_INIT=16'b0101010111110101;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNITM402_3_LC_4_5_6  (
            .in0(N__5210),
            .in1(_gnd_net_),
            .in2(N__3115),
            .in3(N__4328),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI0TRC3_LC_4_5_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI0TRC3_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI0TRC3_LC_4_5_7 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNI0TRC3_LC_4_5_7  (
            .in0(_gnd_net_),
            .in1(N__5334),
            .in2(N__3196),
            .in3(N__3187),
            .lcout(\U400_SDRAM.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIFAF21_2_LC_4_6_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIFAF21_2_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIFAF21_2_LC_4_6_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIFAF21_2_LC_4_6_0  (
            .in0(N__5057),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4326),
            .lcout(\U400_SDRAM.N_55 ),
            .ltout(\U400_SDRAM.N_55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIHPJJ1_LC_4_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIHPJJ1_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIHPJJ1_LC_4_6_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIHPJJ1_LC_4_6_1  (
            .in0(N__5314),
            .in1(N__4837),
            .in2(N__3193),
            .in3(N__4974),
            .lcout(\U400_SDRAM.N_105 ),
            .ltout(\U400_SDRAM.N_105_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI2J773_LC_4_6_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI2J773_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI2J773_LC_4_6_2 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNI2J773_LC_4_6_2  (
            .in0(N__4975),
            .in1(N__5315),
            .in2(N__3190),
            .in3(N__3186),
            .lcout(\U400_SDRAM.N_62 ),
            .ltout(\U400_SDRAM.N_62_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS0_EN_RNO_0_LC_4_6_3 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0_EN_RNO_0_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.CS0_EN_RNO_0_LC_4_6_3 .LUT_INIT=16'b1111111111010101;
    LogicCell40 \U400_SDRAM.CS0_EN_RNO_0_LC_4_6_3  (
            .in0(N__3159),
            .in1(N__4718),
            .in2(N__3175),
            .in3(N__3567),
            .lcout(),
            .ltout(\U400_SDRAM.N_39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS0_EN_LC_4_6_4 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0_EN_LC_4_6_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.CS0_EN_LC_4_6_4 .LUT_INIT=16'b0011111110111011;
    LogicCell40 \U400_SDRAM.CS0_EN_LC_4_6_4  (
            .in0(N__3276),
            .in1(N__3330),
            .in2(N__3172),
            .in3(N__3657),
            .lcout(\U400_SDRAM.CS0_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0_ENC_net ),
            .ce(),
            .sr(N__6489));
    defparam \U400_SDRAM.CS1_EN_RNO_0_LC_4_6_5 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1_EN_RNO_0_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.CS1_EN_RNO_0_LC_4_6_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U400_SDRAM.CS1_EN_RNO_0_LC_4_6_5  (
            .in0(N__4717),
            .in1(N__3169),
            .in2(N__3163),
            .in3(N__3568),
            .lcout(),
            .ltout(\U400_SDRAM.N_41_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS1_EN_LC_4_6_6 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1_EN_LC_4_6_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.CS1_EN_LC_4_6_6 .LUT_INIT=16'b0011111110111011;
    LogicCell40 \U400_SDRAM.CS1_EN_LC_4_6_6  (
            .in0(N__3225),
            .in1(N__3331),
            .in2(N__3142),
            .in3(N__3658),
            .lcout(\U400_SDRAM.CS1_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0_ENC_net ),
            .ce(),
            .sr(N__6489));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_3_LC_4_7_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_3_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_3_LC_4_7_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_3_LC_4_7_2  (
            .in0(N__4867),
            .in1(N__4976),
            .in2(_gnd_net_),
            .in3(N__5425),
            .lcout(\U400_SDRAM.N_57 ),
            .ltout(\U400_SDRAM.N_57_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIG9NQ3_LC_4_7_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIG9NQ3_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIG9NQ3_LC_4_7_3 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIG9NQ3_LC_4_7_3  (
            .in0(N__5338),
            .in1(N__3308),
            .in2(N__3334),
            .in3(N__4716),
            .lcout(\U400_SDRAM.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIJ1DL_6_LC_4_7_4 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIJ1DL_6_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIJ1DL_6_LC_4_7_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNIJ1DL_6_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(N__3801),
            .in2(_gnd_net_),
            .in3(N__3816),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_o5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNI8CGL1_3_LC_4_7_5 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNI8CGL1_3_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNI8CGL1_3_LC_4_7_5 .LUT_INIT=16'b0011000001110000;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNI8CGL1_3_LC_4_7_5  (
            .in0(N__3606),
            .in1(N__3831),
            .in2(N__3322),
            .in3(N__3591),
            .lcout(\U400_SDRAM.N_266_0 ),
            .ltout(\U400_SDRAM.N_266_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_4_7_6 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_4_7_6 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3319),
            .in3(N__5359),
            .lcout(\U400_SDRAM.SDRAM_CMD12 ),
            .ltout(\U400_SDRAM.SDRAM_CMD12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIG9NQ3_1_LC_4_7_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIG9NQ3_1_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIG9NQ3_1_LC_4_7_7 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIG9NQ3_1_LC_4_7_7  (
            .in0(_gnd_net_),
            .in1(N__4715),
            .in2(N__3295),
            .in3(N__3947),
            .lcout(\U400_SDRAM.un1_SDRAM_COUNTER52_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS0n_LC_4_9_0 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0n_LC_4_9_0 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CS0n_LC_4_9_0 .LUT_INIT=16'b1000000011111111;
    LogicCell40 \U400_SDRAM.CS0n_LC_4_9_0  (
            .in0(N__6770),
            .in1(N__6308),
            .in2(N__6187),
            .in3(N__3277),
            .lcout(CS0n_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0nC_net ),
            .ce(),
            .sr(N__6487));
    defparam \U400_SDRAM.WEn_LC_4_9_3 .C_ON=1'b0;
    defparam \U400_SDRAM.WEn_LC_4_9_3 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.WEn_LC_4_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.WEn_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6163),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0nC_net ),
            .ce(),
            .sr(N__6487));
    defparam \U400_SDRAM.CASn_LC_4_9_5 .C_ON=1'b0;
    defparam \U400_SDRAM.CASn_LC_4_9_5 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CASn_LC_4_9_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U400_SDRAM.CASn_LC_4_9_5  (
            .in0(N__6309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0nC_net ),
            .ce(),
            .sr(N__6487));
    defparam \U400_SDRAM.CS1n_LC_4_10_2 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1n_LC_4_10_2 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CS1n_LC_4_10_2 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \U400_SDRAM.CS1n_LC_4_10_2  (
            .in0(N__6771),
            .in1(N__6292),
            .in2(N__3229),
            .in3(N__6170),
            .lcout(CS1n_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS1nC_net ),
            .ce(),
            .sr(N__6488));
    defparam \U400_SDRAM.MA_nesr_7_LC_4_12_6 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_7_LC_4_12_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_7_LC_4_12_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_7_LC_4_12_6  (
            .in0(N__3427),
            .in1(N__6772),
            .in2(N__3415),
            .in3(N__6659),
            .lcout(MA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_7C_net ),
            .ce(N__6580),
            .sr(N__6490));
    defparam \U400_SDRAM.MA_nesr_6_LC_4_14_0 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_6_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_6_LC_4_14_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_6_LC_4_14_0  (
            .in0(N__3391),
            .in1(N__6776),
            .in2(N__3382),
            .in3(N__6667),
            .lcout(MA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_6C_net ),
            .ce(N__6581),
            .sr(N__6494));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_5_4_0 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_5_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_5_4_0  (
            .in0(_gnd_net_),
            .in1(N__4845),
            .in2(_gnd_net_),
            .in3(N__3355),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(bfn_5_4_0_),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_4_1 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(N__4713),
            .in2(_gnd_net_),
            .in3(N__3352),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_1 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_5_4_2 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_5_4_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_5_4_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_2_LC_5_4_2  (
            .in0(N__5522),
            .in1(N__5067),
            .in2(_gnd_net_),
            .in3(N__3349),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_2 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__5469),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_5_4_3 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_5_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_5_4_3  (
            .in0(_gnd_net_),
            .in1(N__4978),
            .in2(_gnd_net_),
            .in3(N__3346),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_3 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_5_4_4 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_5_4_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_4_LC_5_4_4  (
            .in0(N__5523),
            .in1(N__3481),
            .in2(_gnd_net_),
            .in3(N__3343),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_4 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__5469),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_5_4_5 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_5_4_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_5_4_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_5_LC_5_4_5  (
            .in0(N__5517),
            .in1(N__3465),
            .in2(_gnd_net_),
            .in3(N__3340),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_5 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__5469),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_5_4_6 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_5_4_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_5_4_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_6_LC_5_4_6  (
            .in0(N__5524),
            .in1(N__3499),
            .in2(_gnd_net_),
            .in3(N__3337),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_6 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__5469),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_5_4_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_5_4_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_7_LC_5_4_7  (
            .in0(N__5518),
            .in1(N__3445),
            .in2(_gnd_net_),
            .in3(N__3577),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__5469),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNISRU82_8_LC_5_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNISRU82_8_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNISRU82_8_LC_5_5_0 .LUT_INIT=16'b0010001011111111;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNISRU82_8_LC_5_5_0  (
            .in0(N__5371),
            .in1(N__4546),
            .in2(_gnd_net_),
            .in3(N__3526),
            .lcout(\U400_SDRAM.N_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_RNO_0_LC_5_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_0_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_0_LC_5_5_1 .LUT_INIT=16'b0101110100000000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_RNO_0_LC_5_5_1  (
            .in0(N__3528),
            .in1(N__5373),
            .in2(N__4555),
            .in3(N__4367),
            .lcout(\U400_SDRAM.N_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_6_2_LC_5_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_6_2_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_6_2_LC_5_5_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_6_2_LC_5_5_2  (
            .in0(N__5208),
            .in1(N__3480),
            .in2(_gnd_net_),
            .in3(N__3444),
            .lcout(\U400_SDRAM.SDRAM_CMD_cnst_0_76_i_a4_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIDLIS3_8_LC_5_5_3 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIDLIS3_8_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIDLIS3_8_LC_5_5_3 .LUT_INIT=16'b0101000100000000;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNIDLIS3_8_LC_5_5_3  (
            .in0(N__3527),
            .in1(N__5372),
            .in2(N__4554),
            .in3(N__3937),
            .lcout(\U400_SDRAM.N_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_5_5_4 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_5_5_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_5_5_4  (
            .in0(N__3559),
            .in1(N__5670),
            .in2(N__5710),
            .in3(N__5631),
            .lcout(),
            .ltout(\U400_SDRAM.un3_RAM_CYCLE_START_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_5_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_5_5_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_5_5_5 .LUT_INIT=16'b1111001000000000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_LC_5_5_5  (
            .in0(N__3529),
            .in1(N__3864),
            .in2(N__3544),
            .in3(N__5207),
            .lcout(\U400_SDRAM.RAM_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4043),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_5_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_5_6  (
            .in0(N__3497),
            .in1(N__3479),
            .in2(N__3466),
            .in3(N__3443),
            .lcout(\U400_SDRAM.N_54 ),
            .ltout(\U400_SDRAM.N_54_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_2_LC_5_5_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_2_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_2_LC_5_5_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_2_LC_5_5_7  (
            .in0(N__4848),
            .in1(N__5039),
            .in2(N__3430),
            .in3(N__4366),
            .lcout(\U400_SDRAM.SDRAM_COUNTER42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI24955_1_LC_5_6_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI24955_1_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI24955_1_LC_5_6_2 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI24955_1_LC_5_6_2  (
            .in0(N__5404),
            .in1(N__3942),
            .in2(N__3667),
            .in3(N__4711),
            .lcout(\U400_SDRAM.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_3_LC_5_6_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_3_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_3_LC_5_6_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U400_SDRAM.TACK_RNO_3_LC_5_6_3  (
            .in0(N__4838),
            .in1(N__5426),
            .in2(N__4719),
            .in3(N__4489),
            .lcout(\U400_SDRAM.TACK_4_m ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_1_LC_5_6_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_1_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_1_LC_5_6_5 .LUT_INIT=16'b1011001110110011;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_1_LC_5_6_5  (
            .in0(N__3943),
            .in1(N__5189),
            .in2(N__4720),
            .in3(_gnd_net_),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_5_6_6 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_5_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_0_LC_5_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3632),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_0C_net ),
            .ce(),
            .sr(N__3783));
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_5_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_5_6_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_1_LC_5_6_7  (
            .in0(N__3633),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3649),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_0C_net ),
            .ce(),
            .sr(N__3783));
    defparam \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_5_7_0 .C_ON=1'b1;
    defparam \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_5_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(N__3648),
            .in2(N__3637),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_5_7_1 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_5_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_2_LC_5_7_1  (
            .in0(_gnd_net_),
            .in1(N__3616),
            .in2(_gnd_net_),
            .in3(N__3610),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_1 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_2 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3784));
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_5_7_2 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_5_7_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_5_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_3_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(N__3607),
            .in2(_gnd_net_),
            .in3(N__3595),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_2 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_3 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3784));
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_5_7_3 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_5_7_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_5_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_4_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(N__3592),
            .in2(_gnd_net_),
            .in3(N__3580),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_3 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_4 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3784));
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_5_7_4 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_5_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_5_LC_5_7_4  (
            .in0(_gnd_net_),
            .in1(N__3832),
            .in2(_gnd_net_),
            .in3(N__3820),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_4 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_5 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3784));
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_5_7_5 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_5_7_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_5_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_6_LC_5_7_5  (
            .in0(_gnd_net_),
            .in1(N__3817),
            .in2(_gnd_net_),
            .in3(N__3805),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_5 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_6 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3784));
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_5_7_6 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_5_7_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_5_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_7_LC_5_7_6  (
            .in0(_gnd_net_),
            .in1(N__3802),
            .in2(_gnd_net_),
            .in3(N__3790),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_6 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_7 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3784));
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_5_7_7 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_5_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_8_LC_5_7_7  (
            .in0(_gnd_net_),
            .in1(N__5370),
            .in2(_gnd_net_),
            .in3(N__3787),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3784));
    defparam \U400_SDRAM.MA_nesr_8_LC_5_12_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_8_LC_5_12_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_8_LC_5_12_7 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_8_LC_5_12_7  (
            .in0(N__3772),
            .in1(N__6823),
            .in2(N__3757),
            .in3(N__6658),
            .lcout(MA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_8C_net ),
            .ce(N__6554),
            .sr(N__6491));
    defparam \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_5_13_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_5_13_0 .LUT_INIT=16'b1111011011110111;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_5_13_0  (
            .in0(N__6821),
            .in1(N__6307),
            .in2(N__6517),
            .in3(N__6171),
            .lcout(\U400_SDRAM.un1_MA20_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_9_LC_5_14_2 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_9_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_9_LC_5_14_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.MA_nesr_9_LC_5_14_2  (
            .in0(N__6822),
            .in1(N__6306),
            .in2(N__3727),
            .in3(N__6196),
            .lcout(MA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_9C_net ),
            .ce(N__6579),
            .sr(N__6500));
    defparam \U400_SDRAM.WRITE_CYCLE_LC_6_3_5 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_LC_6_3_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.WRITE_CYCLE_LC_6_3_5 .LUT_INIT=16'b1010101000101110;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_LC_6_3_5  (
            .in0(N__4483),
            .in1(N__3700),
            .in2(N__3679),
            .in3(N__3904),
            .lcout(\U400_SDRAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.WRITE_CYCLEC_net ),
            .ce(),
            .sr(N__6502));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_6_4_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_6_4_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_6_4_0  (
            .in0(N__6402),
            .in1(N__3954),
            .in2(N__5585),
            .in3(N__3895),
            .lcout(\U400_SDRAM.N_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_OUT_LC_6_4_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_LC_6_4_3 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.TA_OUT_LC_6_4_3 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \U400_SDRAM.TA_OUT_LC_6_4_3  (
            .in0(N__4141),
            .in1(N__4102),
            .in2(N__4074),
            .in3(N__4093),
            .lcout(TA_OUT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4051),
            .ce(),
            .sr(N__6496));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI8O963_LC_6_4_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI8O963_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNI8O963_LC_6_4_7 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNI8O963_LC_6_4_7  (
            .in0(N__5212),
            .in1(N__4498),
            .in2(_gnd_net_),
            .in3(N__4337),
            .lcout(\U400_SDRAM.N_303_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIFGBJ4_1_LC_6_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIFGBJ4_1_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIFGBJ4_1_LC_6_5_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIFGBJ4_1_LC_6_5_0  (
            .in0(N__4672),
            .in1(N__3955),
            .in2(N__5228),
            .in3(N__3896),
            .lcout(\U400_SDRAM.SDRAM_CMD_5_sqmuxa ),
            .ltout(\U400_SDRAM.SDRAM_CMD_5_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_LC_6_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_LC_6_5_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.RAM_CYCLE_LC_6_5_1 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_LC_6_5_1  (
            .in0(N__4222),
            .in1(N__3865),
            .in2(N__3874),
            .in3(N__3871),
            .lcout(\U400_SDRAM.RAM_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.RAM_CYCLEC_net ),
            .ce(),
            .sr(N__6492));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIQ4PD_3_LC_6_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIQ4PD_3_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIQ4PD_3_LC_6_5_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIQ4PD_3_LC_6_5_2  (
            .in0(_gnd_net_),
            .in1(N__4917),
            .in2(_gnd_net_),
            .in3(N__4637),
            .lcout(\U400_SDRAM.N_94_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIOLQ51_LC_6_5_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIOLQ51_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIOLQ51_LC_6_5_4 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIOLQ51_LC_6_5_4  (
            .in0(N__5056),
            .in1(N__5308),
            .in2(_gnd_net_),
            .in3(N__4329),
            .lcout(\U400_SDRAM.N_30_2 ),
            .ltout(\U400_SDRAM.N_30_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_5_5 .LUT_INIT=16'b1101111111011101;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_5_5  (
            .in0(N__5203),
            .in1(N__4185),
            .in2(N__3847),
            .in3(N__4371),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_6_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_6_5_6 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_6_5_6  (
            .in0(N__4174),
            .in1(N__4490),
            .in2(N__3844),
            .in3(N__5309),
            .lcout(\U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_RNO_1_LC_6_5_7 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_1_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.RAM_CYCLE_RNO_1_LC_6_5_7 .LUT_INIT=16'b1111101111111100;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_RNO_1_LC_6_5_7  (
            .in0(N__4918),
            .in1(N__4798),
            .in2(N__4231),
            .in3(N__4673),
            .lcout(\U400_SDRAM.un1_SDRAM_COUNTER52_2_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIN1PD_0_LC_6_6_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIN1PD_0_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIN1PD_0_LC_6_6_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIN1PD_0_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__4770),
            .in2(_gnd_net_),
            .in3(N__4638),
            .lcout(\U400_SDRAM.N_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNII7IR_2_LC_6_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNII7IR_2_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNII7IR_2_LC_6_6_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNII7IR_2_LC_6_6_1  (
            .in0(N__4639),
            .in1(N__5058),
            .in2(N__4810),
            .in3(N__4944),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_COUNTER44_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIPKQB2_3_LC_6_6_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIPKQB2_3_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIPKQB2_3_LC_6_6_2 .LUT_INIT=16'b1111111100001110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIPKQB2_3_LC_6_6_2  (
            .in0(N__4945),
            .in1(N__5444),
            .in2(N__4216),
            .in3(N__4330),
            .lcout(\U400_SDRAM.un1_SDRAM_COUNTER44_0 ),
            .ltout(\U400_SDRAM.un1_SDRAM_COUNTER44_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_0_LC_6_6_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_0_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_0_LC_6_6_3 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \U400_SDRAM.TACK_RNO_0_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4213),
            .in3(N__4488),
            .lcout(\U400_SDRAM.N_117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.WRITE_CYCLE_RNIPAEV_LC_6_6_4 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_RNIPAEV_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.WRITE_CYCLE_RNIPAEV_LC_6_6_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_RNIPAEV_LC_6_6_4  (
            .in0(N__5059),
            .in1(N__4774),
            .in2(N__4492),
            .in3(N__4365),
            .lcout(\U400_SDRAM.N_108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_4_LC_6_6_5 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_4_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_4_LC_6_6_5 .LUT_INIT=16'b1100111100101111;
    LogicCell40 \U400_SDRAM.TACK_RNO_4_LC_6_6_5  (
            .in0(N__5445),
            .in1(N__5060),
            .in2(N__5333),
            .in3(N__4946),
            .lcout(),
            .ltout(\U400_SDRAM.un1_SDRAM_COUNTER52_4_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_2_LC_6_6_6 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_2_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_2_LC_6_6_6 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \U400_SDRAM.TACK_RNO_2_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(N__4387),
            .in2(N__4201),
            .in3(N__4331),
            .lcout(\U400_SDRAM.un1_SDRAM_COUNTER52_4_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TACK_RNO_1_LC_6_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_RNO_1_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TACK_RNO_1_LC_6_6_7 .LUT_INIT=16'b0000000010110001;
    LogicCell40 \U400_SDRAM.TACK_RNO_1_LC_6_6_7  (
            .in0(N__4491),
            .in1(N__4186),
            .in2(N__4173),
            .in3(N__4156),
            .lcout(\U400_SDRAM.TACK_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIP3PD_3_LC_6_7_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIP3PD_3_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNIP3PD_3_LC_6_7_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNIP3PD_3_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(N__4852),
            .in2(_gnd_net_),
            .in3(N__4962),
            .lcout(\U400_SDRAM.N_56 ),
            .ltout(\U400_SDRAM.N_56_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_7_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_7_1 .LUT_INIT=16'b0000111110001000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_7_1  (
            .in0(N__4964),
            .in1(N__5062),
            .in2(N__4390),
            .in3(N__4712),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_o2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_6_7_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_6_7_2 .LUT_INIT=16'b0000000011111100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(N__4386),
            .in2(N__4375),
            .in3(N__4338),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_6_7_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_6_7_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_6_7_3  (
            .in0(N__5332),
            .in1(N__4856),
            .in2(N__5075),
            .in3(N__4372),
            .lcout(),
            .ltout(\U400_SDRAM.N_275_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_6_7_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_6_7_4 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_6_7_4  (
            .in0(N__5181),
            .in1(N__4291),
            .in2(N__4342),
            .in3(N__4339),
            .lcout(\U400_SDRAM.N_270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_6_7_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_6_7_6 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_6_7_6  (
            .in0(N__5061),
            .in1(N__4963),
            .in2(N__4865),
            .in3(N__4687),
            .lcout(\U400_SDRAM.N_276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_12_LC_6_12_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_12_LC_6_12_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_12_LC_6_12_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U400_SDRAM.MA_nesr_12_LC_6_12_7  (
            .in0(N__6188),
            .in1(N__4285),
            .in2(N__6310),
            .in3(N__6834),
            .lcout(MA_c_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_12C_net ),
            .ce(N__6597),
            .sr(N__6495));
    defparam \U400_SDRAM.MA_nesr_10_LC_6_13_4 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_10_LC_6_13_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_10_LC_6_13_4 .LUT_INIT=16'b0100000001000100;
    LogicCell40 \U400_SDRAM.MA_nesr_10_LC_6_13_4  (
            .in0(N__6847),
            .in1(N__6305),
            .in2(N__4258),
            .in3(N__6195),
            .lcout(MA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_10C_net ),
            .ce(N__6569),
            .sr(N__6501));
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_LC_7_3_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.RAM_SPACE_LC_7_3_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U400_ADDRESS_DECODE.RAM_SPACE_LC_7_3_2  (
            .in0(N__5627),
            .in1(N__5669),
            .in2(_gnd_net_),
            .in3(N__5709),
            .lcout(RAM_SPACEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un2_LLBEn_0_LC_7_3_6 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un2_LLBEn_0_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un2_LLBEn_0_LC_7_3_6 .LUT_INIT=16'b0001010000111100;
    LogicCell40 \U400_BYTE_ENABLE.un2_LLBEn_0_LC_7_3_6  (
            .in0(N__5760),
            .in1(N__6403),
            .in2(N__5587),
            .in3(N__5803),
            .lcout(),
            .ltout(\U400_BYTE_ENABLE.un2_LLBEn_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_LC_7_3_7 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_LLBEn_i_LC_7_3_7 .LUT_INIT=16'b0111010111110101;
    LogicCell40 \U400_BYTE_ENABLE.un1_LLBEn_i_LC_7_3_7  (
            .in0(N__5839),
            .in1(N__5759),
            .in2(N__4525),
            .in3(N__5581),
            .lcout(U400_BYTE_ENABLE_un1_LLBEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_2_LC_7_4_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_2_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_3_2_LC_7_4_0 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_3_2_LC_7_4_0  (
            .in0(N__4925),
            .in1(N__4792),
            .in2(_gnd_net_),
            .in3(N__5211),
            .lcout(\U400_SDRAM.SDRAM_CMD_cnst_0_76_i_a4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIE01O_LC_7_4_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIE01O_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIE01O_LC_7_4_2 .LUT_INIT=16'b1111110001111110;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIE01O_LC_7_4_2  (
            .in0(N__4647),
            .in1(N__4791),
            .in2(N__4961),
            .in3(N__5329),
            .lcout(),
            .ltout(\U400_SDRAM.N_321_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIGMQQ1_LC_7_4_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIGMQQ1_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIGMQQ1_LC_7_4_3 .LUT_INIT=16'b1101110111110000;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIGMQQ1_LC_7_4_3  (
            .in0(N__5330),
            .in1(N__4441),
            .in2(N__4501),
            .in3(N__5066),
            .lcout(\U400_SDRAM.N_322_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_7_4_7 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_7_4_7 .LUT_INIT=16'b1100110000010011;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_7_4_7  (
            .in0(N__4790),
            .in1(N__4924),
            .in2(N__4484),
            .in3(N__4646),
            .lcout(\U400_SDRAM.N_320_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_7_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_7_5_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_7_5_1 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_0_LC_7_5_1  (
            .in0(N__5519),
            .in1(N__5380),
            .in2(N__4435),
            .in3(N__4420),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_0C_net ),
            .ce(N__5470),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_7_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_7_5_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_7_5_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_3_LC_7_5_6  (
            .in0(N__5491),
            .in1(N__4414),
            .in2(N__6348),
            .in3(N__5521),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_0C_net ),
            .ce(N__5470),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_7_5_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_7_5_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_7_5_7 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_1_LC_7_5_7  (
            .in0(N__5520),
            .in1(N__5490),
            .in2(N__6347),
            .in3(N__5482),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_0C_net ),
            .ce(N__5470),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_7_6_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_7_6_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_LC_7_6_4  (
            .in0(N__5304),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5403),
            .lcout(\U400_SDRAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CONFIGUREDC_net ),
            .ce(),
            .sr(N__6493));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_7_6_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_7_6_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_7_6_6  (
            .in0(N__5446),
            .in1(N__4952),
            .in2(N__5331),
            .in3(N__5431),
            .lcout(\U400_SDRAM.SDRAM_CMD_3_sqmuxa ),
            .ltout(\U400_SDRAM.SDRAM_CMD_3_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_7_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_7_6_7 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_7_6_7  (
            .in0(N__5182),
            .in1(N__5303),
            .in2(N__5389),
            .in3(N__5386),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_5_1_LC_7_7_2 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_5_1_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_5_1_LC_7_7_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_5_1_LC_7_7_2  (
            .in0(N__5374),
            .in1(N__4833),
            .in2(_gnd_net_),
            .in3(N__5076),
            .lcout(\U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_a5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_LC_7_7_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_LC_7_7_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_LC_7_7_3  (
            .in0(N__5310),
            .in1(N__5164),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U400_SDRAM.N_299_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_7_7_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_7_7_5 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_7_7_5  (
            .in0(N__5077),
            .in1(N__4971),
            .in2(N__4857),
            .in3(N__4691),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_0_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_7_7_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_7_7_6 .LUT_INIT=16'b1111001101110011;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_7_7_6  (
            .in0(N__4585),
            .in1(N__4572),
            .in2(N__4558),
            .in3(N__4553),
            .lcout(),
            .ltout(\U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_7_7_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_7_7_7 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_1_LC_7_7_7  (
            .in0(N__6255),
            .in1(N__5923),
            .in2(N__5914),
            .in3(N__5911),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_11_LC_7_13_6 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_11_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_11_LC_7_13_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.MA_nesr_11_LC_7_13_6  (
            .in0(N__6842),
            .in1(N__6301),
            .in2(N__5887),
            .in3(N__6194),
            .lcout(MA_c_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_11C_net ),
            .ce(N__6588),
            .sr(N__6503));
    defparam \U400_BYTE_ENABLE.un1_UMBEn_i_LC_8_3_3 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_UMBEn_i_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_UMBEn_i_LC_8_3_3 .LUT_INIT=16'b1011111100110011;
    LogicCell40 \U400_BYTE_ENABLE.un1_UMBEn_i_LC_8_3_3  (
            .in0(N__5765),
            .in1(N__5841),
            .in2(N__5586),
            .in3(N__5728),
            .lcout(U400_BYTE_ENABLE_un1_UMBEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_LMBEn_i_LC_8_3_4 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_LMBEn_i_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_LMBEn_i_LC_8_3_4 .LUT_INIT=16'b1111010101110101;
    LogicCell40 \U400_BYTE_ENABLE.un1_LMBEn_i_LC_8_3_4  (
            .in0(N__5840),
            .in1(N__5764),
            .in2(N__5722),
            .in3(N__5804),
            .lcout(U400_BYTE_ENABLE_un1_LMBEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un1_UUBEn_i_LC_8_3_5 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un1_UUBEn_i_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un1_UUBEn_i_LC_8_3_5 .LUT_INIT=16'b1111101100110011;
    LogicCell40 \U400_BYTE_ENABLE.un1_UUBEn_i_LC_8_3_5  (
            .in0(N__5766),
            .in1(N__5842),
            .in2(N__5811),
            .in3(N__5721),
            .lcout(U400_BYTE_ENABLE_un1_UUBEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.un2_UMBEn_0_LC_8_4_4 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.un2_UMBEn_0_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.un2_UMBEn_0_LC_8_4_4 .LUT_INIT=16'b0011000111000100;
    LogicCell40 \U400_BYTE_ENABLE.un2_UMBEn_0_LC_8_4_4  (
            .in0(N__5812),
            .in1(N__6401),
            .in2(N__5767),
            .in3(N__5565),
            .lcout(\U400_BYTE_ENABLE.un2_UMBEn_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_BYTE_ENABLE.LW_TRANS_LC_8_4_5 .C_ON=1'b0;
    defparam \U400_BYTE_ENABLE.LW_TRANS_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \U400_BYTE_ENABLE.LW_TRANS_LC_8_4_5 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \U400_BYTE_ENABLE.LW_TRANS_LC_8_4_5  (
            .in0(N__6400),
            .in1(_gnd_net_),
            .in2(N__5577),
            .in3(_gnd_net_),
            .lcout(\U400_BYTE_ENABLE.LW_TRANS_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.RAM_SPACEm_i_LC_8_4_7 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.RAM_SPACEm_i_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.RAM_SPACEm_i_LC_8_4_7 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U400_ADDRESS_DECODE.RAM_SPACEm_i_LC_8_4_7  (
            .in0(N__5705),
            .in1(N__5671),
            .in2(_gnd_net_),
            .in3(N__5632),
            .lcout(RAM_SPACEm_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.BURST8_LC_8_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.BURST8_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.BURST8_LC_8_5_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U400_SDRAM.BURST8_LC_8_5_6  (
            .in0(N__5561),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6388),
            .lcout(\U400_SDRAM.BURSTZ0Z8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_8_12_0 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_8_12_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_8_12_0  (
            .in0(N__6839),
            .in1(N__6286),
            .in2(_gnd_net_),
            .in3(N__6197),
            .lcout(\U400_SDRAM.MA19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_RNO_0_5_LC_8_14_1 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_RNO_0_5_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.MA_nesr_RNO_0_5_LC_8_14_1 .LUT_INIT=16'b0011111100101110;
    LogicCell40 \U400_SDRAM.MA_nesr_RNO_0_5_LC_8_14_1  (
            .in0(N__6198),
            .in1(N__6841),
            .in2(N__6322),
            .in3(N__6288),
            .lcout(\U400_SDRAM.MA_5_iv_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_RNO_0_1_LC_8_14_6 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_RNO_0_1_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.MA_nesr_RNO_0_1_LC_8_14_6 .LUT_INIT=16'b0101111101001110;
    LogicCell40 \U400_SDRAM.MA_nesr_RNO_0_1_LC_8_14_6  (
            .in0(N__6840),
            .in1(N__6287),
            .in2(N__6214),
            .in3(N__6199),
            .lcout(\U400_SDRAM.MA_5_iv_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_5_LC_8_15_4 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_5_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_5_LC_8_15_4 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \U400_SDRAM.MA_nesr_5_LC_8_15_4  (
            .in0(N__6094),
            .in1(N__6082),
            .in2(_gnd_net_),
            .in3(N__6648),
            .lcout(MA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_5C_net ),
            .ce(N__6593),
            .sr(N__6505));
    defparam \U400_SDRAM.MA_nesr_3_LC_9_13_2 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_3_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_3_LC_9_13_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_3_LC_9_13_2  (
            .in0(N__6061),
            .in1(N__6843),
            .in2(N__6052),
            .in3(N__6638),
            .lcout(MA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_3C_net ),
            .ce(N__6592),
            .sr(N__6504));
    defparam \U400_SDRAM.MA_nesr_4_LC_9_15_0 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_4_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_4_LC_9_15_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_4_LC_9_15_0  (
            .in0(N__6846),
            .in1(N__6019),
            .in2(N__6007),
            .in3(N__6666),
            .lcout(MA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_4C_net ),
            .ce(N__6598),
            .sr(N__6506));
    defparam \U400_SDRAM.MA_nesr_0_LC_9_15_1 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_0_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_0_LC_9_15_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \U400_SDRAM.MA_nesr_0_LC_9_15_1  (
            .in0(N__6664),
            .in1(N__5974),
            .in2(N__5962),
            .in3(N__6844),
            .lcout(MA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_4C_net ),
            .ce(N__6598),
            .sr(N__6506));
    defparam \U400_SDRAM.MA_nesr_1_LC_9_15_4 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_1_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_1_LC_9_15_4 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \U400_SDRAM.MA_nesr_1_LC_9_15_4  (
            .in0(N__5938),
            .in1(N__5929),
            .in2(_gnd_net_),
            .in3(N__6663),
            .lcout(MA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_4C_net ),
            .ce(N__6598),
            .sr(N__6506));
    defparam \U400_SDRAM.MA_nesr_2_LC_9_15_6 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_2_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_2_LC_9_15_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_2_LC_9_15_6  (
            .in0(N__6845),
            .in1(N__6691),
            .in2(N__6679),
            .in3(N__6665),
            .lcout(MA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_4C_net ),
            .ce(N__6598),
            .sr(N__6506));
    defparam TAn_obuft_RNO_LC_11_6_6.C_ON=1'b0;
    defparam TAn_obuft_RNO_LC_11_6_6.SEQ_MODE=4'b0000;
    defparam TAn_obuft_RNO_LC_11_6_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 TAn_obuft_RNO_LC_11_6_6 (
            .in0(N__6424),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_474_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U400_TOP

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Sep 14 2025 20:14:53

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    DRA,
    CMA,
    DA,
    A,
    TBIn,
    RAMSPACEn,
    DBRn,
    RAMENn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    PRnW,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    BLSn,
    TCIn,
    WEn,
    REGENn,
    LLBEn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    input [1:0] SIZ;
    input [9:0] DRA;
    output [10:0] CMA;
    output [2:0] DA;
    input [20:0] A;
    output TBIn;
    input RAMSPACEn;
    input DBRn;
    output RAMENn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output PRnW;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    output BLSn;
    output TCIn;
    output WEn;
    output REGENn;
    output LLBEn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__13239;
    wire N__13238;
    wire N__13237;
    wire N__13230;
    wire N__13229;
    wire N__13228;
    wire N__13221;
    wire N__13220;
    wire N__13219;
    wire N__13212;
    wire N__13211;
    wire N__13210;
    wire N__13203;
    wire N__13202;
    wire N__13201;
    wire N__13194;
    wire N__13193;
    wire N__13192;
    wire N__13185;
    wire N__13184;
    wire N__13183;
    wire N__13176;
    wire N__13175;
    wire N__13174;
    wire N__13167;
    wire N__13166;
    wire N__13165;
    wire N__13158;
    wire N__13157;
    wire N__13156;
    wire N__13149;
    wire N__13148;
    wire N__13147;
    wire N__13140;
    wire N__13139;
    wire N__13138;
    wire N__13131;
    wire N__13130;
    wire N__13129;
    wire N__13122;
    wire N__13121;
    wire N__13120;
    wire N__13113;
    wire N__13112;
    wire N__13111;
    wire N__13104;
    wire N__13103;
    wire N__13102;
    wire N__13095;
    wire N__13094;
    wire N__13093;
    wire N__13086;
    wire N__13085;
    wire N__13084;
    wire N__13077;
    wire N__13076;
    wire N__13075;
    wire N__13068;
    wire N__13067;
    wire N__13066;
    wire N__13059;
    wire N__13058;
    wire N__13057;
    wire N__13050;
    wire N__13049;
    wire N__13048;
    wire N__13041;
    wire N__13040;
    wire N__13039;
    wire N__13032;
    wire N__13031;
    wire N__13030;
    wire N__13023;
    wire N__13022;
    wire N__13021;
    wire N__13014;
    wire N__13013;
    wire N__13012;
    wire N__13005;
    wire N__13004;
    wire N__13003;
    wire N__12996;
    wire N__12995;
    wire N__12994;
    wire N__12987;
    wire N__12986;
    wire N__12985;
    wire N__12978;
    wire N__12977;
    wire N__12976;
    wire N__12969;
    wire N__12968;
    wire N__12967;
    wire N__12960;
    wire N__12959;
    wire N__12958;
    wire N__12951;
    wire N__12950;
    wire N__12949;
    wire N__12942;
    wire N__12941;
    wire N__12940;
    wire N__12933;
    wire N__12932;
    wire N__12931;
    wire N__12924;
    wire N__12923;
    wire N__12922;
    wire N__12915;
    wire N__12914;
    wire N__12913;
    wire N__12906;
    wire N__12905;
    wire N__12904;
    wire N__12897;
    wire N__12896;
    wire N__12895;
    wire N__12888;
    wire N__12887;
    wire N__12886;
    wire N__12879;
    wire N__12878;
    wire N__12877;
    wire N__12870;
    wire N__12869;
    wire N__12868;
    wire N__12861;
    wire N__12860;
    wire N__12859;
    wire N__12852;
    wire N__12851;
    wire N__12850;
    wire N__12843;
    wire N__12842;
    wire N__12841;
    wire N__12834;
    wire N__12833;
    wire N__12832;
    wire N__12825;
    wire N__12824;
    wire N__12823;
    wire N__12816;
    wire N__12815;
    wire N__12814;
    wire N__12807;
    wire N__12806;
    wire N__12805;
    wire N__12798;
    wire N__12797;
    wire N__12796;
    wire N__12789;
    wire N__12788;
    wire N__12787;
    wire N__12780;
    wire N__12779;
    wire N__12778;
    wire N__12771;
    wire N__12770;
    wire N__12769;
    wire N__12762;
    wire N__12761;
    wire N__12760;
    wire N__12753;
    wire N__12752;
    wire N__12751;
    wire N__12744;
    wire N__12743;
    wire N__12742;
    wire N__12735;
    wire N__12734;
    wire N__12733;
    wire N__12726;
    wire N__12725;
    wire N__12724;
    wire N__12717;
    wire N__12716;
    wire N__12715;
    wire N__12708;
    wire N__12707;
    wire N__12706;
    wire N__12699;
    wire N__12698;
    wire N__12697;
    wire N__12690;
    wire N__12689;
    wire N__12688;
    wire N__12681;
    wire N__12680;
    wire N__12679;
    wire N__12672;
    wire N__12671;
    wire N__12670;
    wire N__12663;
    wire N__12662;
    wire N__12661;
    wire N__12654;
    wire N__12653;
    wire N__12652;
    wire N__12645;
    wire N__12644;
    wire N__12643;
    wire N__12636;
    wire N__12635;
    wire N__12634;
    wire N__12627;
    wire N__12626;
    wire N__12625;
    wire N__12618;
    wire N__12617;
    wire N__12616;
    wire N__12609;
    wire N__12608;
    wire N__12607;
    wire N__12600;
    wire N__12599;
    wire N__12598;
    wire N__12591;
    wire N__12590;
    wire N__12589;
    wire N__12582;
    wire N__12581;
    wire N__12580;
    wire N__12573;
    wire N__12572;
    wire N__12571;
    wire N__12564;
    wire N__12563;
    wire N__12562;
    wire N__12555;
    wire N__12554;
    wire N__12553;
    wire N__12546;
    wire N__12545;
    wire N__12544;
    wire N__12537;
    wire N__12536;
    wire N__12535;
    wire N__12528;
    wire N__12527;
    wire N__12526;
    wire N__12519;
    wire N__12518;
    wire N__12517;
    wire N__12510;
    wire N__12509;
    wire N__12508;
    wire N__12501;
    wire N__12500;
    wire N__12499;
    wire N__12492;
    wire N__12491;
    wire N__12490;
    wire N__12483;
    wire N__12482;
    wire N__12481;
    wire N__12474;
    wire N__12473;
    wire N__12472;
    wire N__12465;
    wire N__12464;
    wire N__12463;
    wire N__12456;
    wire N__12455;
    wire N__12454;
    wire N__12447;
    wire N__12446;
    wire N__12445;
    wire N__12438;
    wire N__12437;
    wire N__12436;
    wire N__12429;
    wire N__12428;
    wire N__12427;
    wire N__12420;
    wire N__12419;
    wire N__12418;
    wire N__12411;
    wire N__12410;
    wire N__12409;
    wire N__12402;
    wire N__12401;
    wire N__12400;
    wire N__12393;
    wire N__12392;
    wire N__12391;
    wire N__12384;
    wire N__12383;
    wire N__12382;
    wire N__12375;
    wire N__12374;
    wire N__12373;
    wire N__12366;
    wire N__12365;
    wire N__12364;
    wire N__12347;
    wire N__12344;
    wire N__12341;
    wire N__12338;
    wire N__12335;
    wire N__12334;
    wire N__12333;
    wire N__12332;
    wire N__12329;
    wire N__12326;
    wire N__12323;
    wire N__12320;
    wire N__12313;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12301;
    wire N__12300;
    wire N__12299;
    wire N__12296;
    wire N__12293;
    wire N__12290;
    wire N__12287;
    wire N__12280;
    wire N__12277;
    wire N__12274;
    wire N__12271;
    wire N__12268;
    wire N__12265;
    wire N__12262;
    wire N__12259;
    wire N__12256;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12238;
    wire N__12235;
    wire N__12234;
    wire N__12233;
    wire N__12230;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12194;
    wire N__12191;
    wire N__12188;
    wire N__12185;
    wire N__12182;
    wire N__12179;
    wire N__12176;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12160;
    wire N__12157;
    wire N__12152;
    wire N__12149;
    wire N__12146;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12130;
    wire N__12129;
    wire N__12128;
    wire N__12127;
    wire N__12126;
    wire N__12125;
    wire N__12124;
    wire N__12123;
    wire N__12122;
    wire N__12121;
    wire N__12120;
    wire N__12119;
    wire N__12118;
    wire N__12117;
    wire N__12116;
    wire N__12115;
    wire N__12114;
    wire N__12113;
    wire N__12112;
    wire N__12111;
    wire N__12110;
    wire N__12109;
    wire N__12108;
    wire N__12107;
    wire N__12106;
    wire N__12105;
    wire N__12104;
    wire N__12103;
    wire N__12102;
    wire N__12101;
    wire N__12100;
    wire N__12099;
    wire N__12098;
    wire N__12097;
    wire N__12096;
    wire N__12095;
    wire N__12094;
    wire N__12093;
    wire N__12092;
    wire N__12089;
    wire N__12088;
    wire N__12087;
    wire N__12086;
    wire N__12085;
    wire N__12084;
    wire N__12083;
    wire N__12082;
    wire N__12081;
    wire N__12080;
    wire N__12079;
    wire N__12078;
    wire N__11975;
    wire N__11972;
    wire N__11971;
    wire N__11968;
    wire N__11965;
    wire N__11962;
    wire N__11959;
    wire N__11956;
    wire N__11953;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11939;
    wire N__11936;
    wire N__11933;
    wire N__11930;
    wire N__11929;
    wire N__11928;
    wire N__11927;
    wire N__11926;
    wire N__11925;
    wire N__11924;
    wire N__11923;
    wire N__11920;
    wire N__11919;
    wire N__11918;
    wire N__11913;
    wire N__11910;
    wire N__11907;
    wire N__11904;
    wire N__11903;
    wire N__11902;
    wire N__11899;
    wire N__11896;
    wire N__11895;
    wire N__11894;
    wire N__11893;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11876;
    wire N__11871;
    wire N__11870;
    wire N__11869;
    wire N__11866;
    wire N__11863;
    wire N__11858;
    wire N__11855;
    wire N__11852;
    wire N__11849;
    wire N__11840;
    wire N__11837;
    wire N__11834;
    wire N__11831;
    wire N__11818;
    wire N__11817;
    wire N__11816;
    wire N__11815;
    wire N__11810;
    wire N__11803;
    wire N__11798;
    wire N__11795;
    wire N__11790;
    wire N__11785;
    wire N__11782;
    wire N__11779;
    wire N__11776;
    wire N__11773;
    wire N__11768;
    wire N__11765;
    wire N__11764;
    wire N__11763;
    wire N__11760;
    wire N__11755;
    wire N__11754;
    wire N__11749;
    wire N__11746;
    wire N__11741;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11723;
    wire N__11722;
    wire N__11721;
    wire N__11720;
    wire N__11719;
    wire N__11718;
    wire N__11717;
    wire N__11702;
    wire N__11699;
    wire N__11696;
    wire N__11695;
    wire N__11694;
    wire N__11693;
    wire N__11692;
    wire N__11691;
    wire N__11690;
    wire N__11689;
    wire N__11688;
    wire N__11687;
    wire N__11686;
    wire N__11685;
    wire N__11684;
    wire N__11683;
    wire N__11682;
    wire N__11651;
    wire N__11648;
    wire N__11645;
    wire N__11644;
    wire N__11643;
    wire N__11642;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11632;
    wire N__11629;
    wire N__11626;
    wire N__11625;
    wire N__11624;
    wire N__11623;
    wire N__11622;
    wire N__11621;
    wire N__11620;
    wire N__11619;
    wire N__11618;
    wire N__11617;
    wire N__11616;
    wire N__11615;
    wire N__11612;
    wire N__11611;
    wire N__11610;
    wire N__11609;
    wire N__11608;
    wire N__11607;
    wire N__11606;
    wire N__11605;
    wire N__11604;
    wire N__11603;
    wire N__11602;
    wire N__11601;
    wire N__11600;
    wire N__11599;
    wire N__11598;
    wire N__11597;
    wire N__11596;
    wire N__11595;
    wire N__11594;
    wire N__11593;
    wire N__11592;
    wire N__11591;
    wire N__11590;
    wire N__11587;
    wire N__11586;
    wire N__11585;
    wire N__11584;
    wire N__11581;
    wire N__11580;
    wire N__11579;
    wire N__11578;
    wire N__11577;
    wire N__11576;
    wire N__11575;
    wire N__11574;
    wire N__11573;
    wire N__11572;
    wire N__11571;
    wire N__11570;
    wire N__11569;
    wire N__11568;
    wire N__11565;
    wire N__11564;
    wire N__11563;
    wire N__11562;
    wire N__11559;
    wire N__11558;
    wire N__11557;
    wire N__11556;
    wire N__11435;
    wire N__11432;
    wire N__11429;
    wire N__11426;
    wire N__11425;
    wire N__11424;
    wire N__11421;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11411;
    wire N__11408;
    wire N__11405;
    wire N__11402;
    wire N__11399;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11389;
    wire N__11386;
    wire N__11383;
    wire N__11378;
    wire N__11375;
    wire N__11370;
    wire N__11367;
    wire N__11362;
    wire N__11357;
    wire N__11354;
    wire N__11353;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11335;
    wire N__11332;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11315;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11286;
    wire N__11281;
    wire N__11280;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11256;
    wire N__11253;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11241;
    wire N__11234;
    wire N__11231;
    wire N__11228;
    wire N__11225;
    wire N__11224;
    wire N__11223;
    wire N__11220;
    wire N__11219;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11204;
    wire N__11199;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11182;
    wire N__11177;
    wire N__11174;
    wire N__11171;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11151;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11139;
    wire N__11132;
    wire N__11131;
    wire N__11130;
    wire N__11129;
    wire N__11126;
    wire N__11125;
    wire N__11124;
    wire N__11123;
    wire N__11120;
    wire N__11119;
    wire N__11116;
    wire N__11115;
    wire N__11114;
    wire N__11113;
    wire N__11112;
    wire N__11109;
    wire N__11108;
    wire N__11105;
    wire N__11104;
    wire N__11103;
    wire N__11102;
    wire N__11101;
    wire N__11100;
    wire N__11097;
    wire N__11096;
    wire N__11095;
    wire N__11094;
    wire N__11093;
    wire N__11090;
    wire N__11085;
    wire N__11082;
    wire N__11077;
    wire N__11072;
    wire N__11067;
    wire N__11066;
    wire N__11065;
    wire N__11062;
    wire N__11059;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11048;
    wire N__11045;
    wire N__11044;
    wire N__11041;
    wire N__11038;
    wire N__11033;
    wire N__11028;
    wire N__11025;
    wire N__11022;
    wire N__11019;
    wire N__11012;
    wire N__11005;
    wire N__11002;
    wire N__11001;
    wire N__10998;
    wire N__10997;
    wire N__10996;
    wire N__10995;
    wire N__10994;
    wire N__10993;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10973;
    wire N__10970;
    wire N__10963;
    wire N__10962;
    wire N__10961;
    wire N__10960;
    wire N__10959;
    wire N__10948;
    wire N__10945;
    wire N__10942;
    wire N__10939;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10900;
    wire N__10891;
    wire N__10888;
    wire N__10873;
    wire N__10868;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10838;
    wire N__10837;
    wire N__10834;
    wire N__10833;
    wire N__10830;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10806;
    wire N__10803;
    wire N__10798;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10750;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10739;
    wire N__10736;
    wire N__10731;
    wire N__10728;
    wire N__10725;
    wire N__10720;
    wire N__10717;
    wire N__10714;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10657;
    wire N__10654;
    wire N__10651;
    wire N__10646;
    wire N__10645;
    wire N__10644;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10573;
    wire N__10572;
    wire N__10571;
    wire N__10570;
    wire N__10569;
    wire N__10568;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10558;
    wire N__10557;
    wire N__10554;
    wire N__10553;
    wire N__10550;
    wire N__10549;
    wire N__10548;
    wire N__10545;
    wire N__10544;
    wire N__10543;
    wire N__10542;
    wire N__10541;
    wire N__10540;
    wire N__10539;
    wire N__10536;
    wire N__10535;
    wire N__10534;
    wire N__10531;
    wire N__10530;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10517;
    wire N__10512;
    wire N__10505;
    wire N__10502;
    wire N__10497;
    wire N__10492;
    wire N__10491;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10476;
    wire N__10471;
    wire N__10462;
    wire N__10461;
    wire N__10460;
    wire N__10457;
    wire N__10452;
    wire N__10451;
    wire N__10450;
    wire N__10443;
    wire N__10442;
    wire N__10441;
    wire N__10440;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10425;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10401;
    wire N__10398;
    wire N__10393;
    wire N__10388;
    wire N__10385;
    wire N__10374;
    wire N__10371;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10327;
    wire N__10326;
    wire N__10325;
    wire N__10322;
    wire N__10321;
    wire N__10320;
    wire N__10319;
    wire N__10316;
    wire N__10315;
    wire N__10312;
    wire N__10309;
    wire N__10306;
    wire N__10303;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10293;
    wire N__10290;
    wire N__10287;
    wire N__10284;
    wire N__10279;
    wire N__10272;
    wire N__10269;
    wire N__10266;
    wire N__10261;
    wire N__10258;
    wire N__10255;
    wire N__10244;
    wire N__10243;
    wire N__10242;
    wire N__10241;
    wire N__10238;
    wire N__10235;
    wire N__10234;
    wire N__10233;
    wire N__10232;
    wire N__10229;
    wire N__10228;
    wire N__10227;
    wire N__10226;
    wire N__10225;
    wire N__10224;
    wire N__10221;
    wire N__10218;
    wire N__10215;
    wire N__10212;
    wire N__10205;
    wire N__10198;
    wire N__10193;
    wire N__10188;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10153;
    wire N__10150;
    wire N__10147;
    wire N__10146;
    wire N__10145;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10131;
    wire N__10128;
    wire N__10125;
    wire N__10122;
    wire N__10117;
    wire N__10114;
    wire N__10111;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10078;
    wire N__10075;
    wire N__10072;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10045;
    wire N__10042;
    wire N__10039;
    wire N__10038;
    wire N__10035;
    wire N__10034;
    wire N__10033;
    wire N__10032;
    wire N__10029;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10021;
    wire N__10020;
    wire N__10017;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__10000;
    wire N__9997;
    wire N__9994;
    wire N__9987;
    wire N__9980;
    wire N__9971;
    wire N__9970;
    wire N__9969;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9946;
    wire N__9943;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9922;
    wire N__9919;
    wire N__9916;
    wire N__9915;
    wire N__9914;
    wire N__9909;
    wire N__9906;
    wire N__9903;
    wire N__9898;
    wire N__9895;
    wire N__9892;
    wire N__9889;
    wire N__9886;
    wire N__9883;
    wire N__9880;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9863;
    wire N__9860;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9823;
    wire N__9818;
    wire N__9815;
    wire N__9814;
    wire N__9813;
    wire N__9810;
    wire N__9809;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9790;
    wire N__9787;
    wire N__9784;
    wire N__9783;
    wire N__9782;
    wire N__9781;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9767;
    wire N__9762;
    wire N__9759;
    wire N__9746;
    wire N__9743;
    wire N__9742;
    wire N__9739;
    wire N__9736;
    wire N__9733;
    wire N__9730;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9685;
    wire N__9680;
    wire N__9679;
    wire N__9678;
    wire N__9677;
    wire N__9676;
    wire N__9675;
    wire N__9674;
    wire N__9673;
    wire N__9672;
    wire N__9671;
    wire N__9670;
    wire N__9669;
    wire N__9668;
    wire N__9667;
    wire N__9666;
    wire N__9663;
    wire N__9660;
    wire N__9655;
    wire N__9652;
    wire N__9647;
    wire N__9642;
    wire N__9635;
    wire N__9634;
    wire N__9633;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9623;
    wire N__9622;
    wire N__9621;
    wire N__9620;
    wire N__9619;
    wire N__9616;
    wire N__9613;
    wire N__9602;
    wire N__9595;
    wire N__9590;
    wire N__9587;
    wire N__9580;
    wire N__9577;
    wire N__9570;
    wire N__9567;
    wire N__9566;
    wire N__9565;
    wire N__9564;
    wire N__9563;
    wire N__9560;
    wire N__9553;
    wire N__9548;
    wire N__9545;
    wire N__9540;
    wire N__9537;
    wire N__9532;
    wire N__9529;
    wire N__9520;
    wire N__9515;
    wire N__9512;
    wire N__9511;
    wire N__9510;
    wire N__9509;
    wire N__9508;
    wire N__9505;
    wire N__9496;
    wire N__9491;
    wire N__9490;
    wire N__9487;
    wire N__9486;
    wire N__9483;
    wire N__9478;
    wire N__9473;
    wire N__9472;
    wire N__9471;
    wire N__9468;
    wire N__9463;
    wire N__9462;
    wire N__9457;
    wire N__9454;
    wire N__9451;
    wire N__9446;
    wire N__9445;
    wire N__9442;
    wire N__9441;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9429;
    wire N__9426;
    wire N__9423;
    wire N__9420;
    wire N__9417;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9406;
    wire N__9403;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9377;
    wire N__9368;
    wire N__9365;
    wire N__9364;
    wire N__9363;
    wire N__9362;
    wire N__9361;
    wire N__9360;
    wire N__9357;
    wire N__9356;
    wire N__9355;
    wire N__9352;
    wire N__9351;
    wire N__9350;
    wire N__9349;
    wire N__9342;
    wire N__9341;
    wire N__9340;
    wire N__9339;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9316;
    wire N__9313;
    wire N__9304;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9100;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9073;
    wire N__9072;
    wire N__9069;
    wire N__9066;
    wire N__9063;
    wire N__9060;
    wire N__9057;
    wire N__9054;
    wire N__9053;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9043;
    wire N__9038;
    wire N__9037;
    wire N__9028;
    wire N__9025;
    wire N__9020;
    wire N__9017;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9007;
    wire N__9004;
    wire N__9001;
    wire N__8998;
    wire N__8995;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8962;
    wire N__8959;
    wire N__8958;
    wire N__8957;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8949;
    wire N__8946;
    wire N__8943;
    wire N__8940;
    wire N__8935;
    wire N__8928;
    wire N__8925;
    wire N__8922;
    wire N__8915;
    wire N__8912;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8898;
    wire N__8895;
    wire N__8892;
    wire N__8889;
    wire N__8886;
    wire N__8883;
    wire N__8880;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8864;
    wire N__8861;
    wire N__8856;
    wire N__8853;
    wire N__8846;
    wire N__8845;
    wire N__8842;
    wire N__8841;
    wire N__8840;
    wire N__8839;
    wire N__8838;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8824;
    wire N__8817;
    wire N__8814;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8792;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8782;
    wire N__8779;
    wire N__8774;
    wire N__8773;
    wire N__8770;
    wire N__8767;
    wire N__8766;
    wire N__8761;
    wire N__8758;
    wire N__8755;
    wire N__8750;
    wire N__8749;
    wire N__8748;
    wire N__8745;
    wire N__8744;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8731;
    wire N__8728;
    wire N__8725;
    wire N__8722;
    wire N__8719;
    wire N__8716;
    wire N__8711;
    wire N__8706;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8617;
    wire N__8616;
    wire N__8613;
    wire N__8610;
    wire N__8607;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8521;
    wire N__8518;
    wire N__8515;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8491;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8464;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8446;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8431;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8372;
    wire N__8369;
    wire N__8366;
    wire N__8363;
    wire N__8362;
    wire N__8361;
    wire N__8358;
    wire N__8355;
    wire N__8354;
    wire N__8351;
    wire N__8350;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8321;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8285;
    wire N__8282;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8267;
    wire N__8266;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8219;
    wire N__8216;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8197;
    wire N__8192;
    wire N__8191;
    wire N__8188;
    wire N__8185;
    wire N__8180;
    wire N__8179;
    wire N__8178;
    wire N__8177;
    wire N__8172;
    wire N__8169;
    wire N__8166;
    wire N__8159;
    wire N__8156;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8144;
    wire N__8141;
    wire N__8138;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8126;
    wire N__8125;
    wire N__8124;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8113;
    wire N__8110;
    wire N__8109;
    wire N__8108;
    wire N__8107;
    wire N__8106;
    wire N__8101;
    wire N__8098;
    wire N__8097;
    wire N__8096;
    wire N__8095;
    wire N__8094;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8078;
    wire N__8073;
    wire N__8068;
    wire N__8061;
    wire N__8048;
    wire N__8045;
    wire N__8044;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8029;
    wire N__8026;
    wire N__8023;
    wire N__8020;
    wire N__8017;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7984;
    wire N__7981;
    wire N__7978;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7844;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7825;
    wire N__7822;
    wire N__7819;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7804;
    wire N__7803;
    wire N__7802;
    wire N__7801;
    wire N__7800;
    wire N__7797;
    wire N__7792;
    wire N__7785;
    wire N__7778;
    wire N__7777;
    wire N__7776;
    wire N__7775;
    wire N__7770;
    wire N__7765;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7751;
    wire N__7750;
    wire N__7747;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7737;
    wire N__7730;
    wire N__7729;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7672;
    wire N__7669;
    wire N__7666;
    wire N__7663;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7642;
    wire N__7639;
    wire N__7636;
    wire N__7633;
    wire N__7630;
    wire N__7627;
    wire N__7624;
    wire N__7621;
    wire N__7618;
    wire N__7613;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7601;
    wire N__7598;
    wire N__7595;
    wire N__7592;
    wire N__7591;
    wire N__7588;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7570;
    wire N__7567;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7532;
    wire N__7531;
    wire N__7528;
    wire N__7525;
    wire N__7522;
    wire N__7517;
    wire N__7516;
    wire N__7513;
    wire N__7510;
    wire N__7507;
    wire N__7502;
    wire N__7501;
    wire N__7498;
    wire N__7495;
    wire N__7490;
    wire N__7489;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7465;
    wire N__7462;
    wire N__7459;
    wire N__7454;
    wire N__7453;
    wire N__7452;
    wire N__7449;
    wire N__7446;
    wire N__7443;
    wire N__7442;
    wire N__7441;
    wire N__7440;
    wire N__7437;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7414;
    wire N__7411;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7391;
    wire N__7390;
    wire N__7389;
    wire N__7386;
    wire N__7383;
    wire N__7376;
    wire N__7373;
    wire N__7370;
    wire N__7367;
    wire N__7366;
    wire N__7365;
    wire N__7364;
    wire N__7359;
    wire N__7356;
    wire N__7353;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7321;
    wire N__7320;
    wire N__7319;
    wire N__7318;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7303;
    wire N__7300;
    wire N__7293;
    wire N__7290;
    wire N__7287;
    wire N__7282;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7267;
    wire N__7264;
    wire N__7261;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7241;
    wire N__7238;
    wire N__7235;
    wire N__7232;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7219;
    wire N__7216;
    wire N__7213;
    wire N__7210;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7181;
    wire N__7180;
    wire N__7177;
    wire N__7176;
    wire N__7173;
    wire N__7170;
    wire N__7167;
    wire N__7164;
    wire N__7161;
    wire N__7158;
    wire N__7155;
    wire N__7152;
    wire N__7149;
    wire N__7146;
    wire N__7143;
    wire N__7140;
    wire N__7137;
    wire N__7134;
    wire N__7131;
    wire N__7128;
    wire N__7123;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7109;
    wire N__7106;
    wire N__7103;
    wire N__7100;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7070;
    wire N__7067;
    wire N__7064;
    wire N__7063;
    wire N__7062;
    wire N__7061;
    wire N__7058;
    wire N__7057;
    wire N__7052;
    wire N__7049;
    wire N__7044;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7024;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7003;
    wire N__7002;
    wire N__6999;
    wire N__6996;
    wire N__6995;
    wire N__6992;
    wire N__6989;
    wire N__6984;
    wire N__6977;
    wire N__6974;
    wire N__6973;
    wire N__6972;
    wire N__6971;
    wire N__6968;
    wire N__6965;
    wire N__6960;
    wire N__6953;
    wire N__6950;
    wire N__6947;
    wire N__6944;
    wire N__6941;
    wire N__6940;
    wire N__6939;
    wire N__6938;
    wire N__6937;
    wire N__6936;
    wire N__6935;
    wire N__6934;
    wire N__6933;
    wire N__6932;
    wire N__6911;
    wire N__6908;
    wire N__6905;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6892;
    wire N__6889;
    wire N__6886;
    wire N__6881;
    wire N__6880;
    wire N__6877;
    wire N__6874;
    wire N__6869;
    wire N__6868;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6854;
    wire N__6853;
    wire N__6850;
    wire N__6847;
    wire N__6842;
    wire N__6841;
    wire N__6838;
    wire N__6835;
    wire N__6830;
    wire N__6829;
    wire N__6826;
    wire N__6823;
    wire N__6818;
    wire N__6815;
    wire N__6814;
    wire N__6811;
    wire N__6808;
    wire N__6803;
    wire N__6802;
    wire N__6799;
    wire N__6798;
    wire N__6795;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6781;
    wire N__6778;
    wire N__6771;
    wire N__6768;
    wire N__6765;
    wire N__6762;
    wire N__6755;
    wire N__6752;
    wire N__6749;
    wire N__6746;
    wire N__6745;
    wire N__6742;
    wire N__6739;
    wire N__6734;
    wire N__6731;
    wire N__6730;
    wire N__6727;
    wire N__6724;
    wire N__6721;
    wire N__6718;
    wire N__6717;
    wire N__6712;
    wire N__6709;
    wire N__6708;
    wire N__6705;
    wire N__6702;
    wire N__6699;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6655;
    wire N__6652;
    wire N__6651;
    wire N__6650;
    wire N__6649;
    wire N__6648;
    wire N__6647;
    wire N__6644;
    wire N__6643;
    wire N__6640;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6619;
    wire N__6612;
    wire N__6609;
    wire N__6606;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6584;
    wire N__6581;
    wire N__6578;
    wire N__6577;
    wire N__6576;
    wire N__6573;
    wire N__6568;
    wire N__6563;
    wire N__6560;
    wire N__6557;
    wire N__6554;
    wire N__6551;
    wire N__6550;
    wire N__6547;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6502;
    wire N__6501;
    wire N__6500;
    wire N__6499;
    wire N__6498;
    wire N__6497;
    wire N__6496;
    wire N__6495;
    wire N__6494;
    wire N__6493;
    wire N__6492;
    wire N__6489;
    wire N__6488;
    wire N__6485;
    wire N__6482;
    wire N__6481;
    wire N__6478;
    wire N__6471;
    wire N__6470;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6462;
    wire N__6459;
    wire N__6450;
    wire N__6449;
    wire N__6448;
    wire N__6447;
    wire N__6446;
    wire N__6445;
    wire N__6444;
    wire N__6443;
    wire N__6442;
    wire N__6439;
    wire N__6434;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6417;
    wire N__6414;
    wire N__6409;
    wire N__6404;
    wire N__6397;
    wire N__6390;
    wire N__6381;
    wire N__6362;
    wire N__6361;
    wire N__6360;
    wire N__6357;
    wire N__6356;
    wire N__6353;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6329;
    wire N__6328;
    wire N__6327;
    wire N__6326;
    wire N__6325;
    wire N__6324;
    wire N__6323;
    wire N__6322;
    wire N__6319;
    wire N__6318;
    wire N__6317;
    wire N__6316;
    wire N__6313;
    wire N__6312;
    wire N__6311;
    wire N__6304;
    wire N__6301;
    wire N__6296;
    wire N__6295;
    wire N__6292;
    wire N__6291;
    wire N__6290;
    wire N__6289;
    wire N__6288;
    wire N__6287;
    wire N__6280;
    wire N__6279;
    wire N__6278;
    wire N__6277;
    wire N__6270;
    wire N__6269;
    wire N__6268;
    wire N__6267;
    wire N__6264;
    wire N__6259;
    wire N__6258;
    wire N__6255;
    wire N__6252;
    wire N__6247;
    wire N__6240;
    wire N__6237;
    wire N__6230;
    wire N__6227;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6188;
    wire N__6185;
    wire N__6182;
    wire N__6181;
    wire N__6180;
    wire N__6177;
    wire N__6176;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6133;
    wire N__6132;
    wire N__6131;
    wire N__6130;
    wire N__6129;
    wire N__6128;
    wire N__6125;
    wire N__6124;
    wire N__6123;
    wire N__6120;
    wire N__6117;
    wire N__6114;
    wire N__6111;
    wire N__6110;
    wire N__6105;
    wire N__6102;
    wire N__6101;
    wire N__6098;
    wire N__6097;
    wire N__6096;
    wire N__6093;
    wire N__6086;
    wire N__6083;
    wire N__6082;
    wire N__6081;
    wire N__6080;
    wire N__6077;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6059;
    wire N__6052;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6008;
    wire N__6007;
    wire N__6006;
    wire N__6005;
    wire N__6002;
    wire N__5999;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5958;
    wire N__5957;
    wire N__5956;
    wire N__5955;
    wire N__5954;
    wire N__5949;
    wire N__5948;
    wire N__5947;
    wire N__5944;
    wire N__5941;
    wire N__5940;
    wire N__5939;
    wire N__5936;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5924;
    wire N__5923;
    wire N__5920;
    wire N__5917;
    wire N__5910;
    wire N__5905;
    wire N__5900;
    wire N__5895;
    wire N__5882;
    wire N__5881;
    wire N__5880;
    wire N__5879;
    wire N__5876;
    wire N__5875;
    wire N__5874;
    wire N__5873;
    wire N__5870;
    wire N__5869;
    wire N__5864;
    wire N__5863;
    wire N__5858;
    wire N__5857;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5834;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5809;
    wire N__5806;
    wire N__5805;
    wire N__5802;
    wire N__5801;
    wire N__5800;
    wire N__5799;
    wire N__5798;
    wire N__5797;
    wire N__5796;
    wire N__5793;
    wire N__5790;
    wire N__5787;
    wire N__5780;
    wire N__5775;
    wire N__5772;
    wire N__5759;
    wire N__5756;
    wire N__5753;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5729;
    wire N__5728;
    wire N__5727;
    wire N__5726;
    wire N__5723;
    wire N__5720;
    wire N__5715;
    wire N__5708;
    wire N__5705;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5653;
    wire N__5648;
    wire N__5645;
    wire N__5644;
    wire N__5643;
    wire N__5636;
    wire N__5635;
    wire N__5634;
    wire N__5633;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5596;
    wire N__5593;
    wire N__5592;
    wire N__5591;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5577;
    wire N__5570;
    wire N__5569;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5559;
    wire N__5558;
    wire N__5557;
    wire N__5552;
    wire N__5545;
    wire N__5540;
    wire N__5539;
    wire N__5536;
    wire N__5535;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5519;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5470;
    wire N__5465;
    wire N__5462;
    wire N__5459;
    wire N__5458;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5450;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5440;
    wire N__5435;
    wire N__5426;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5414;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5399;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5387;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5375;
    wire N__5374;
    wire N__5373;
    wire N__5372;
    wire N__5367;
    wire N__5364;
    wire N__5361;
    wire N__5358;
    wire N__5355;
    wire N__5352;
    wire N__5349;
    wire N__5342;
    wire N__5341;
    wire N__5340;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5242;
    wire N__5239;
    wire N__5236;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5189;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5164;
    wire N__5161;
    wire N__5160;
    wire N__5157;
    wire N__5152;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5126;
    wire N__5123;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5115;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5107;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4927;
    wire N__4926;
    wire N__4925;
    wire N__4924;
    wire N__4923;
    wire N__4922;
    wire N__4921;
    wire N__4920;
    wire N__4907;
    wire N__4902;
    wire N__4899;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4864;
    wire N__4859;
    wire N__4858;
    wire N__4857;
    wire N__4856;
    wire N__4855;
    wire N__4854;
    wire N__4853;
    wire N__4850;
    wire N__4841;
    wire N__4836;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4804;
    wire N__4801;
    wire N__4798;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4732;
    wire N__4729;
    wire N__4726;
    wire N__4721;
    wire N__4720;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4708;
    wire N__4707;
    wire N__4704;
    wire N__4699;
    wire N__4694;
    wire N__4691;
    wire N__4688;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4618;
    wire N__4615;
    wire N__4612;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_PLL_i_i;
    wire DBRn_c_i_0;
    wire A_c_8;
    wire LATCH_CLK_c;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.m104_ns_1_cascade_ ;
    wire \U712_CHIP_RAM.N_105_0_cascade_ ;
    wire \U712_CHIP_RAM.N_106_0 ;
    wire \U712_CHIP_RAM.N_106_0_cascade_ ;
    wire \U712_CHIP_RAM.DBENn_8_0 ;
    wire \U712_CHIP_RAM.N_233 ;
    wire DBDIR_c;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ;
    wire AWEn_c;
    wire A_c_18;
    wire A_c_20;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0 ;
    wire CONSTANT_ONE_NET;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ;
    wire bfn_7_11_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.N_206_0_cascade_ ;
    wire \U712_CHIP_RAM.N_214_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.N_216_0_i_cascade_ ;
    wire \U712_CHIP_RAM.N_217_0 ;
    wire \U712_CHIP_RAM.N_216_0_i ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire \U712_CHIP_RAM.N_195_0_cascade_ ;
    wire \U712_CHIP_RAM.N_213_0 ;
    wire \U712_CHIP_RAM.N_189_0 ;
    wire \U712_CHIP_RAM.N_195_0 ;
    wire VBENn_c;
    wire A_c_2;
    wire A_c_5;
    wire A_c_6;
    wire A_c_3;
    wire A_c_7;
    wire A_c_4;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_111_0_cascade_ ;
    wire \U712_CHIP_RAM.N_50 ;
    wire \U712_CHIP_RAM.m138_0 ;
    wire \U712_CHIP_RAM.N_352_mux_cascade_ ;
    wire \U712_CHIP_RAM.N_183_0 ;
    wire \U712_CHIP_RAM.N_137_0_cascade_ ;
    wire \U712_CHIP_RAM.N_178_0 ;
    wire \U712_CHIP_RAM.N_94_0_cascade_ ;
    wire \U712_CHIP_RAM.N_96_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.m92_0_cascade_ ;
    wire \U712_CHIP_RAM.N_190_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_222_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_358_cascade_ ;
    wire \U712_CHIP_RAM.m219_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_2_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2 ;
    wire \U712_CHIP_RAM.N_137_0 ;
    wire \U712_CHIP_RAM.N_142_0_cascade_ ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.SDRAM_COUNTER43 ;
    wire \U712_CHIP_RAM.m207_ns_1_cascade_ ;
    wire \U712_CHIP_RAM.N_206_0 ;
    wire \U712_CHIP_RAM.N_208_0 ;
    wire \U712_CHIP_RAM.m141_ns_1 ;
    wire \U712_CHIP_RAM.N_140_0 ;
    wire \U712_CHIP_RAM.N_140_0_cascade_ ;
    wire \U712_CHIP_RAM.N_103_0 ;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.N_358 ;
    wire \U712_CHIP_RAM.N_188_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0 ;
    wire \U712_CHIP_RAM.N_344 ;
    wire \U712_CHIP_RAM.N_96_0 ;
    wire \U712_CHIP_RAM.m123_0_cascade_ ;
    wire \U712_CHIP_RAM.N_117_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.m92_0 ;
    wire \U712_CHIP_RAM.N_130_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5Z0Z_3_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNIG3845Z0Z_0 ;
    wire \U712_CHIP_RAM.m203_ns_1 ;
    wire \U712_CHIP_RAM.N_363_mux_cascade_ ;
    wire \U712_CHIP_RAM.m186_0 ;
    wire \U712_CHIP_RAM.N_363 ;
    wire \U712_CHIP_RAM.m225_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.N_110_0 ;
    wire \U712_CHIP_RAM.N_112_0 ;
    wire \U712_CHIP_RAM.N_112_0_cascade_ ;
    wire \U712_CHIP_RAM.N_94_0 ;
    wire RAMENn_c;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire REGSPACEn_c;
    wire TSn_c;
    wire U712_REG_SM_START_RST;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_111_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.N_359_cascade_ ;
    wire \U712_CHIP_RAM.N_130_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1 ;
    wire \U712_CHIP_RAM.N_135_0_cascade_ ;
    wire \U712_CHIP_RAM.N_125_0 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_3 ;
    wire \U712_CHIP_RAM.N_204_0 ;
    wire \U712_CHIP_RAM.N_120_0_cascade_ ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ;
    wire C3_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.N_28_0_cascade_ ;
    wire \U712_CHIP_RAM.N_16_0 ;
    wire \U712_CHIP_RAM.N_16_0_cascade_ ;
    wire \U712_CHIP_RAM.N_66_0_cascade_ ;
    wire A_c_0;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_11_8_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH5lt7_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.N_168_0 ;
    wire CPU_TACKm;
    wire \U712_CYCLE_TERM.TACK_RST_0_i ;
    wire U712_REG_SM_STATE_COUNT_5;
    wire \U712_REG_SM.STATE_COUNTZ0Z_6 ;
    wire N_10_0_cascade_;
    wire U712_REG_SM_REG_CYCLE_START;
    wire \U712_CHIP_RAM.N_84_0_cascade_ ;
    wire U712_REG_SM_STATE_COUNT_0;
    wire i66_mux_cascade_;
    wire \U712_CHIP_RAM.m40_nsZ0Z_1 ;
    wire N_10_0;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire U712_REG_SM_STATE_COUNT_7;
    wire \U712_CHIP_RAM.N_21_0 ;
    wire \U712_CHIP_RAM.N_21_0_cascade_ ;
    wire \U712_CHIP_RAM.N_31_0 ;
    wire \U712_CHIP_RAM.N_329 ;
    wire U712_REG_SM_STATE_COUNT_1;
    wire N_20_0_cascade_;
    wire U712_REG_SM_STATE_COUNT_2;
    wire \U712_CHIP_RAM.N_37_0 ;
    wire N_174_0;
    wire UDSn_c;
    wire SIZ_c_0;
    wire \U712_CHIP_RAM.N_326_mux ;
    wire A_c_1;
    wire SIZ_c_1;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire CLK40_PLL;
    wire CLK40_PLL_iso_i;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.m154_0_2 ;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.m154_0_0 ;
    wire A_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire A_c_11;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire \U712_CHIP_RAM.m157_xx_mm_0_0_cascade_ ;
    wire \U712_CHIP_RAM.m157_xx_mm_0_2 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ;
    wire A_c_17;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8 ;
    wire \U712_CHIP_RAM.m162_xx_mm_0_0_cascade_ ;
    wire \U712_CHIP_RAM.m162_xx_mm_0_2_cascade_ ;
    wire CMA_c_8;
    wire U712_CHIP_RAM_m45_0;
    wire REG_TACK;
    wire U712_REG_SM_REG_TACK_7_0;
    wire U712_REG_SM_STATE_COUNT_8;
    wire U712_REG_SM_STATE_COUNT_3;
    wire N_44_0;
    wire N_175_0;
    wire DBRn_c;
    wire DBR_SYNCZ0Z_0;
    wire U712_REG_SM_WRITE_CYCLE;
    wire N_20_0;
    wire PRnW_c;
    wire U712_REG_SM_C3_SYNC_1;
    wire BLSn_c;
    wire \U712_REG_SM.N_20_0_0 ;
    wire N_172_0;
    wire LDSn_c;
    wire RESETn_c_i;
    wire WEn_c;
    wire A_c_16;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.m161_xx_mm_0_0_cascade_ ;
    wire A_c_13;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire \U712_CHIP_RAM.m159_xx_mm_0_0_cascade_ ;
    wire A_c_15;
    wire \U712_CHIP_RAM.m156_xx_mm_0_2 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire A_c_9;
    wire \U712_CHIP_RAM.N_3_0_cascade_ ;
    wire \U712_CHIP_RAM.m156_xx_mm_0_0 ;
    wire N_144_0;
    wire CLMBEn_c;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ;
    wire bfn_13_13_0_;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ;
    wire \U712_CHIP_RAM.N_325 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_1 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ;
    wire DBR_SYNCZ0Z_1;
    wire DBR_SYNC_i_1;
    wire N_33_0;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire \U712_CHIP_RAM.m160_xx_mm_0_0 ;
    wire \U712_CHIP_RAM.m164_0 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.m159_xx_mm_0_2 ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.m161_xx_mm_0_2 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ;
    wire A_c_14;
    wire \U712_CHIP_RAM.m155_0_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_ ;
    wire \U712_CHIP_RAM.m155_0_2 ;
    wire N_68_0;
    wire CUUBEn_c;
    wire N_145_0;
    wire CLLBEn_c;
    wire DBENn_c;
    wire N_71_0;
    wire CUMBEn_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CYCLE_TERM.N_36_0_cascade_ ;
    wire TACK_OUT;
    wire RESETn_c;
    wire \INVU712_CYCLE_TERM.TACK_OUTC_net ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STARTZ0 ;
    wire TACK_EN;
    wire \INVU712_CYCLE_TERM.TACK_ENC_net ;
    wire U712_REG_SM_C1_SYNC_1;
    wire ASn_c;
    wire \U712_REG_SM.N_33_0_0 ;
    wire DMA_LATCH_EN_c;
    wire \U712_CHIP_RAM.m160_xx_mm_0_2 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire \U712_CHIP_RAM.m228_0 ;
    wire \U712_CHIP_RAM.N_343 ;
    wire \U712_CHIP_RAM.DMA_CYCLEm ;
    wire \U712_CHIP_RAM.N_342 ;
    wire A_c_12;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire \U712_CHIP_RAM.N_3_0 ;
    wire CMA_c_10;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_2 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_5 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_3 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_4 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire \U712_CHIP_RAM.m158_xx_mm_0_0 ;
    wire \U712_CHIP_RAM.m154_a2_0 ;
    wire DRA_c_7;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire CASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.m158_xx_mm_0_2 ;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.N_168_0_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DRA_c_3;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire RAS1n_c;
    wire RAS0n_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire CLK80_PLL;
    wire DRA_c_0;
    wire AGNUS_REV_c;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire RnW_c;
    wire \U712_CHIP_RAM.DMA_WRITE_CYCLEZ0 ;
    wire N_323_mux;
    wire CASLn_c;
    wire CASUn_c;
    wire REG_CYCLEm;
    wire \U712_CHIP_RAM.CPU_CYCLEm ;
    wire N_333_mux;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL),
            .REFERENCECLK(N__4517),
            .RESETB(N__4634),
            .BYPASS(GNDG0),
            .PLLOUTCOREA(),
            .SDI(GNDG0),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(GNDG0),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK(GNDG0));
    IO_PAD DBENn_obuf_iopad (
            .OE(N__13239),
            .DIN(N__13238),
            .DOUT(N__13237),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__13239),
            .PADOUT(N__13238),
            .PADIN(N__13237),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9074),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__13230),
            .DIN(N__13229),
            .DOUT(N__13228),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__13230),
            .PADOUT(N__13229),
            .PADIN(N__13228),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__13221),
            .DIN(N__13220),
            .DOUT(N__13219),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__13221),
            .PADOUT(N__13220),
            .PADIN(N__13219),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10595),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__13212),
            .DIN(N__13211),
            .DOUT(N__13210),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__13212),
            .PADOUT(N__13211),
            .PADIN(N__13210),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11315),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__13203),
            .DIN(N__13202),
            .DOUT(N__13201),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__13203),
            .PADOUT(N__13202),
            .PADIN(N__13201),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__13194),
            .DIN(N__13193),
            .DOUT(N__13192),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__13194),
            .PADOUT(N__13193),
            .PADIN(N__13192),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__13185),
            .DIN(N__13184),
            .DOUT(N__13183),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__13185),
            .PADOUT(N__13184),
            .PADIN(N__13183),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__13176),
            .DIN(N__13175),
            .DOUT(N__13174),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__13176),
            .PADOUT(N__13175),
            .PADIN(N__13174),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__13167),
            .DIN(N__13166),
            .DOUT(N__13165),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__13167),
            .PADOUT(N__13166),
            .PADIN(N__13165),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__13158),
            .DIN(N__13157),
            .DOUT(N__13156),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__13158),
            .PADOUT(N__13157),
            .PADIN(N__13156),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__13149),
            .DIN(N__13148),
            .DOUT(N__13147),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__13149),
            .PADOUT(N__13148),
            .PADIN(N__13147),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__13140),
            .DIN(N__13139),
            .DOUT(N__13138),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__13140),
            .PADOUT(N__13139),
            .PADIN(N__13138),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8543),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__13131),
            .DIN(N__13130),
            .DOUT(N__13129),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__13131),
            .PADOUT(N__13130),
            .PADIN(N__13129),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9176),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__13122),
            .DIN(N__13121),
            .DOUT(N__13120),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__13122),
            .PADOUT(N__13121),
            .PADIN(N__13120),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__13113),
            .DIN(N__13112),
            .DOUT(N__13111),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__13113),
            .PADOUT(N__13112),
            .PADIN(N__13111),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5752),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__13104),
            .DIN(N__13103),
            .DOUT(N__13102),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__13104),
            .PADOUT(N__13103),
            .PADIN(N__13102),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__13095),
            .DIN(N__13094),
            .DOUT(N__13093),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__13095),
            .PADOUT(N__13094),
            .PADIN(N__13093),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__13086),
            .DIN(N__13085),
            .DOUT(N__13084),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__13086),
            .PADOUT(N__13085),
            .PADIN(N__13084),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5042),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__13077),
            .DIN(N__13076),
            .DOUT(N__13075),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__13077),
            .PADOUT(N__13076),
            .PADIN(N__13075),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__13068),
            .DIN(N__13067),
            .DOUT(N__13066),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__13068),
            .PADOUT(N__13067),
            .PADIN(N__13066),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__13059),
            .DIN(N__13058),
            .DOUT(N__13057),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__13059),
            .PADOUT(N__13058),
            .PADIN(N__13057),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8384),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__13050),
            .DIN(N__13049),
            .DOUT(N__13048),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__13050),
            .PADOUT(N__13049),
            .PADIN(N__13048),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__13041),
            .DIN(N__13040),
            .DOUT(N__13039),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__13041),
            .PADOUT(N__13040),
            .PADIN(N__13039),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10613),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__13032),
            .DIN(N__13031),
            .DOUT(N__13030),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__13032),
            .PADOUT(N__13031),
            .PADIN(N__13030),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__13023),
            .DIN(N__13022),
            .DOUT(N__13021),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__13023),
            .PADOUT(N__13022),
            .PADIN(N__13021),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9121),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__13014),
            .DIN(N__13013),
            .DOUT(N__13012),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__13014),
            .PADOUT(N__13013),
            .PADIN(N__13012),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9441),
            .DIN0(),
            .DOUT0(N__8898),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__13005),
            .DIN(N__13004),
            .DOUT(N__13003),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__13005),
            .PADOUT(N__13004),
            .PADIN(N__13003),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__12996),
            .DIN(N__12995),
            .DOUT(N__12994),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__12996),
            .PADOUT(N__12995),
            .PADIN(N__12994),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__12987),
            .DIN(N__12986),
            .DOUT(N__12985),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__12987),
            .PADOUT(N__12986),
            .PADIN(N__12985),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__12978),
            .DIN(N__12977),
            .DOUT(N__12976),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__12978),
            .PADOUT(N__12977),
            .PADIN(N__12976),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__12969),
            .DIN(N__12968),
            .DOUT(N__12967),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__12969),
            .PADOUT(N__12968),
            .PADIN(N__12967),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__12960),
            .DIN(N__12959),
            .DOUT(N__12958),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__12960),
            .PADOUT(N__12959),
            .PADIN(N__12958),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9260),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__12951),
            .DIN(N__12950),
            .DOUT(N__12949),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__12951),
            .PADOUT(N__12950),
            .PADIN(N__12949),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__12942),
            .DIN(N__12941),
            .DOUT(N__12940),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__12942),
            .PADOUT(N__12941),
            .PADIN(N__12940),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__12933),
            .DIN(N__12932),
            .DOUT(N__12931),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__12933),
            .PADOUT(N__12932),
            .PADIN(N__12931),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__12924),
            .DIN(N__12923),
            .DOUT(N__12922),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__12924),
            .PADOUT(N__12923),
            .PADIN(N__12922),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__12915),
            .DIN(N__12914),
            .DOUT(N__12913),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__12915),
            .PADOUT(N__12914),
            .PADIN(N__12913),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__12906),
            .DIN(N__12905),
            .DOUT(N__12904),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__12906),
            .PADOUT(N__12905),
            .PADIN(N__12904),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8699),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__12897),
            .DIN(N__12896),
            .DOUT(N__12895),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__12897),
            .PADOUT(N__12896),
            .PADIN(N__12895),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__12888),
            .DIN(N__12887),
            .DOUT(N__12886),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__12888),
            .PADOUT(N__12887),
            .PADIN(N__12886),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__12879),
            .DIN(N__12878),
            .DOUT(N__12877),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__12879),
            .PADOUT(N__12878),
            .PADIN(N__12877),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9287),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_0_iopad (
            .OE(N__12870),
            .DIN(N__12869),
            .DOUT(N__12868),
            .PACKAGEPIN(DA[0]));
    defparam DA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_0_preio (
            .PADOEN(N__12870),
            .PADOUT(N__12869),
            .PADIN(N__12868),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8321),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__12861),
            .DIN(N__12860),
            .DOUT(N__12859),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__12861),
            .PADOUT(N__12860),
            .PADIN(N__12859),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__12852),
            .DIN(N__12851),
            .DOUT(N__12850),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__12852),
            .PADOUT(N__12851),
            .PADIN(N__12850),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10175),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__12843),
            .DIN(N__12842),
            .DOUT(N__12841),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__12843),
            .PADOUT(N__12842),
            .PADIN(N__12841),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8570),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__12834),
            .DIN(N__12833),
            .DOUT(N__12832),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__12834),
            .PADOUT(N__12833),
            .PADIN(N__12832),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8048),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__12825),
            .DIN(N__12824),
            .DOUT(N__12823),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__12825),
            .PADOUT(N__12824),
            .PADIN(N__12823),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__12816),
            .DIN(N__12815),
            .DOUT(N__12814),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__12816),
            .PADOUT(N__12815),
            .PADIN(N__12814),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8240),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__12807),
            .DIN(N__12806),
            .DOUT(N__12805),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__12807),
            .PADOUT(N__12806),
            .PADIN(N__12805),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9445),
            .DIN0(),
            .DOUT0(N__8912),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__12798),
            .DIN(N__12797),
            .DOUT(N__12796),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__12798),
            .PADOUT(N__12797),
            .PADIN(N__12796),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7961),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__12789),
            .DIN(N__12788),
            .DOUT(N__12787),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__12789),
            .PADOUT(N__12788),
            .PADIN(N__12787),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4748),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__12780),
            .DIN(N__12779),
            .DOUT(N__12778),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__12780),
            .PADOUT(N__12779),
            .PADIN(N__12778),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8990),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__12771),
            .DIN(N__12770),
            .DOUT(N__12769),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__12771),
            .PADOUT(N__12770),
            .PADIN(N__12769),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__12762),
            .DIN(N__12761),
            .DOUT(N__12760),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__12762),
            .PADOUT(N__12761),
            .PADIN(N__12760),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_2_iopad (
            .OE(N__12753),
            .DIN(N__12752),
            .DOUT(N__12751),
            .PACKAGEPIN(DA[2]));
    defparam DA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_2_preio (
            .PADOEN(N__12753),
            .PADOUT(N__12752),
            .PADIN(N__12751),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7604),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__12744),
            .DIN(N__12743),
            .DOUT(N__12742),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__12744),
            .PADOUT(N__12743),
            .PADIN(N__12742),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__12735),
            .DIN(N__12734),
            .DOUT(N__12733),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__12735),
            .PADOUT(N__12734),
            .PADIN(N__12733),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__12726),
            .DIN(N__12725),
            .DOUT(N__12724),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__12726),
            .PADOUT(N__12725),
            .PADIN(N__12724),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7694),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__12717),
            .DIN(N__12716),
            .DOUT(N__12715),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__12717),
            .PADOUT(N__12716),
            .PADIN(N__12715),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8273),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__12708),
            .DIN(N__12707),
            .DOUT(N__12706),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__12708),
            .PADOUT(N__12707),
            .PADIN(N__12706),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__12699),
            .DIN(N__12698),
            .DOUT(N__12697),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__12699),
            .PADOUT(N__12698),
            .PADIN(N__12697),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9143),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__12690),
            .DIN(N__12689),
            .DOUT(N__12688),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__12690),
            .PADOUT(N__12689),
            .PADIN(N__12688),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9446),
            .DIN0(),
            .DOUT0(N__8911),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__12681),
            .DIN(N__12680),
            .DOUT(N__12679),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__12681),
            .PADOUT(N__12680),
            .PADIN(N__12679),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6686),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__12672),
            .DIN(N__12671),
            .DOUT(N__12670),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__12672),
            .PADOUT(N__12671),
            .PADIN(N__12670),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__12663),
            .DIN(N__12662),
            .DOUT(N__12661),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__12663),
            .PADOUT(N__12662),
            .PADIN(N__12661),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__12654),
            .DIN(N__12653),
            .DOUT(N__12652),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__12654),
            .PADOUT(N__12653),
            .PADIN(N__12652),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7859),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__12645),
            .DIN(N__12644),
            .DOUT(N__12643),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__12645),
            .PADOUT(N__12644),
            .PADIN(N__12643),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__12636),
            .DIN(N__12635),
            .DOUT(N__12634),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__12636),
            .PADOUT(N__12635),
            .PADIN(N__12634),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_1_iopad (
            .OE(N__12627),
            .DIN(N__12626),
            .DOUT(N__12625),
            .PACKAGEPIN(DA[1]));
    defparam DA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_1_preio (
            .PADOEN(N__12627),
            .PADOUT(N__12626),
            .PADIN(N__12625),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7652),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__12618),
            .DIN(N__12617),
            .DOUT(N__12616),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__12618),
            .PADOUT(N__12617),
            .PADIN(N__12616),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__12609),
            .DIN(N__12608),
            .DOUT(N__12607),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__12609),
            .PADOUT(N__12608),
            .PADIN(N__12607),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__12600),
            .DIN(N__12599),
            .DOUT(N__12598),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__12600),
            .PADOUT(N__12599),
            .PADIN(N__12598),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8600),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__12591),
            .DIN(N__12590),
            .DOUT(N__12589),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__12591),
            .PADOUT(N__12590),
            .PADIN(N__12589),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7475),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__12582),
            .DIN(N__12581),
            .DOUT(N__12580),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__12582),
            .PADOUT(N__12581),
            .PADIN(N__12580),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9016),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__12573),
            .DIN(N__12572),
            .DOUT(N__12571),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__12573),
            .PADOUT(N__12572),
            .PADIN(N__12571),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5258),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__12564),
            .DIN(N__12563),
            .DOUT(N__12562),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__12564),
            .PADOUT(N__12563),
            .PADIN(N__12562),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__12555),
            .DIN(N__12554),
            .DOUT(N__12553),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__12555),
            .PADOUT(N__12554),
            .PADIN(N__12553),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__12546),
            .DIN(N__12545),
            .DOUT(N__12544),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__12546),
            .PADOUT(N__12545),
            .PADIN(N__12544),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9233),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__12537),
            .DIN(N__12536),
            .DOUT(N__12535),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__12537),
            .PADOUT(N__12536),
            .PADIN(N__12535),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__12528),
            .DIN(N__12527),
            .DOUT(N__12526),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__12528),
            .PADOUT(N__12527),
            .PADIN(N__12526),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__12519),
            .DIN(N__12518),
            .DOUT(N__12517),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__12519),
            .PADOUT(N__12518),
            .PADIN(N__12517),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4544),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__12510),
            .DIN(N__12509),
            .DOUT(N__12508),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__12510),
            .PADOUT(N__12509),
            .PADIN(N__12508),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7994),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__12501),
            .DIN(N__12500),
            .DOUT(N__12499),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__12501),
            .PADOUT(N__12500),
            .PADIN(N__12499),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7180),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PRnW_obuf_iopad (
            .OE(N__12492),
            .DIN(N__12491),
            .DOUT(N__12490),
            .PACKAGEPIN(PRnW));
    defparam PRnW_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PRnW_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PRnW_obuf_preio (
            .PADOEN(N__12492),
            .PADOUT(N__12491),
            .PADIN(N__12490),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8150),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__12483),
            .DIN(N__12482),
            .DOUT(N__12481),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__12483),
            .PADOUT(N__12482),
            .PADIN(N__12481),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__12474),
            .DIN(N__12473),
            .DOUT(N__12472),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__12474),
            .PADOUT(N__12473),
            .PADIN(N__12472),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7181),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__12465),
            .DIN(N__12464),
            .DOUT(N__12463),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__12465),
            .PADOUT(N__12464),
            .PADIN(N__12463),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4583),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__12456),
            .DIN(N__12455),
            .DOUT(N__12454),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__12456),
            .PADOUT(N__12455),
            .PADIN(N__12454),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10346),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__12447),
            .DIN(N__12446),
            .DOUT(N__12445),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__12447),
            .PADOUT(N__12446),
            .PADIN(N__12445),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__12438),
            .DIN(N__12437),
            .DOUT(N__12436),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__12438),
            .PADOUT(N__12437),
            .PADIN(N__12436),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__12429),
            .DIN(N__12428),
            .DOUT(N__12427),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__12429),
            .PADOUT(N__12428),
            .PADIN(N__12427),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BLSn_obuf_iopad (
            .OE(N__12420),
            .DIN(N__12419),
            .DOUT(N__12418),
            .PACKAGEPIN(BLSn));
    defparam BLSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BLSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BLSn_obuf_preio (
            .PADOEN(N__12420),
            .PADOUT(N__12419),
            .PADIN(N__12418),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8044),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__12411),
            .DIN(N__12410),
            .DOUT(N__12409),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__12411),
            .PADOUT(N__12410),
            .PADIN(N__12409),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__12402),
            .DIN(N__12401),
            .DOUT(N__12400),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__12402),
            .PADOUT(N__12401),
            .PADIN(N__12400),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7176),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__12393),
            .DIN(N__12392),
            .DOUT(N__12391),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__12393),
            .PADOUT(N__12392),
            .PADIN(N__12391),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10853),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__12384),
            .DIN(N__12383),
            .DOUT(N__12382),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__12384),
            .PADOUT(N__12383),
            .PADIN(N__12382),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9095),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__12375),
            .DIN(N__12374),
            .DOUT(N__12373),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__12375),
            .PADOUT(N__12374),
            .PADIN(N__12373),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8660),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__12366),
            .DIN(N__12365),
            .DOUT(N__12364),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__12366),
            .PADOUT(N__12365),
            .PADIN(N__12364),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__3007 (
            .O(N__12347),
            .I(N__12344));
    LocalMux I__3006 (
            .O(N__12344),
            .I(N__12341));
    Odrv12 I__3005 (
            .O(N__12341),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__3004 (
            .O(N__12338),
            .I(N__12335));
    LocalMux I__3003 (
            .O(N__12335),
            .I(N__12329));
    InMux I__3002 (
            .O(N__12334),
            .I(N__12326));
    InMux I__3001 (
            .O(N__12333),
            .I(N__12323));
    InMux I__3000 (
            .O(N__12332),
            .I(N__12320));
    Span4Mux_h I__2999 (
            .O(N__12329),
            .I(N__12313));
    LocalMux I__2998 (
            .O(N__12326),
            .I(N__12313));
    LocalMux I__2997 (
            .O(N__12323),
            .I(N__12313));
    LocalMux I__2996 (
            .O(N__12320),
            .I(N__12308));
    Sp12to4 I__2995 (
            .O(N__12313),
            .I(N__12308));
    Span12Mux_v I__2994 (
            .O(N__12308),
            .I(N__12305));
    Odrv12 I__2993 (
            .O(N__12305),
            .I(DRA_c_3));
    InMux I__2992 (
            .O(N__12302),
            .I(N__12296));
    InMux I__2991 (
            .O(N__12301),
            .I(N__12293));
    InMux I__2990 (
            .O(N__12300),
            .I(N__12290));
    InMux I__2989 (
            .O(N__12299),
            .I(N__12287));
    LocalMux I__2988 (
            .O(N__12296),
            .I(N__12280));
    LocalMux I__2987 (
            .O(N__12293),
            .I(N__12280));
    LocalMux I__2986 (
            .O(N__12290),
            .I(N__12280));
    LocalMux I__2985 (
            .O(N__12287),
            .I(N__12277));
    Span4Mux_v I__2984 (
            .O(N__12280),
            .I(N__12274));
    Span4Mux_v I__2983 (
            .O(N__12277),
            .I(N__12271));
    Span4Mux_v I__2982 (
            .O(N__12274),
            .I(N__12268));
    Span4Mux_v I__2981 (
            .O(N__12271),
            .I(N__12265));
    Sp12to4 I__2980 (
            .O(N__12268),
            .I(N__12262));
    Sp12to4 I__2979 (
            .O(N__12265),
            .I(N__12259));
    Span12Mux_h I__2978 (
            .O(N__12262),
            .I(N__12256));
    Odrv12 I__2977 (
            .O(N__12259),
            .I(DRA_c_4));
    Odrv12 I__2976 (
            .O(N__12256),
            .I(DRA_c_4));
    InMux I__2975 (
            .O(N__12251),
            .I(N__12248));
    LocalMux I__2974 (
            .O(N__12248),
            .I(N__12245));
    Odrv4 I__2973 (
            .O(N__12245),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2972 (
            .O(N__12242),
            .I(N__12239));
    LocalMux I__2971 (
            .O(N__12239),
            .I(N__12235));
    InMux I__2970 (
            .O(N__12238),
            .I(N__12230));
    Span4Mux_h I__2969 (
            .O(N__12235),
            .I(N__12227));
    InMux I__2968 (
            .O(N__12234),
            .I(N__12224));
    InMux I__2967 (
            .O(N__12233),
            .I(N__12221));
    LocalMux I__2966 (
            .O(N__12230),
            .I(N__12218));
    Sp12to4 I__2965 (
            .O(N__12227),
            .I(N__12209));
    LocalMux I__2964 (
            .O(N__12224),
            .I(N__12209));
    LocalMux I__2963 (
            .O(N__12221),
            .I(N__12209));
    Sp12to4 I__2962 (
            .O(N__12218),
            .I(N__12209));
    Span12Mux_v I__2961 (
            .O(N__12209),
            .I(N__12206));
    Odrv12 I__2960 (
            .O(N__12206),
            .I(DRA_c_2));
    InMux I__2959 (
            .O(N__12203),
            .I(N__12200));
    LocalMux I__2958 (
            .O(N__12200),
            .I(N__12197));
    Span4Mux_h I__2957 (
            .O(N__12197),
            .I(N__12194));
    Span4Mux_h I__2956 (
            .O(N__12194),
            .I(N__12191));
    Odrv4 I__2955 (
            .O(N__12191),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__2954 (
            .O(N__12188),
            .I(N__12185));
    LocalMux I__2953 (
            .O(N__12185),
            .I(N__12182));
    Span12Mux_h I__2952 (
            .O(N__12182),
            .I(N__12179));
    Odrv12 I__2951 (
            .O(N__12179),
            .I(RAS1n_c));
    InMux I__2950 (
            .O(N__12176),
            .I(N__12172));
    InMux I__2949 (
            .O(N__12175),
            .I(N__12169));
    LocalMux I__2948 (
            .O(N__12172),
            .I(N__12166));
    LocalMux I__2947 (
            .O(N__12169),
            .I(N__12163));
    Span12Mux_v I__2946 (
            .O(N__12166),
            .I(N__12160));
    Span12Mux_h I__2945 (
            .O(N__12163),
            .I(N__12157));
    Odrv12 I__2944 (
            .O(N__12160),
            .I(RAS0n_c));
    Odrv12 I__2943 (
            .O(N__12157),
            .I(RAS0n_c));
    InMux I__2942 (
            .O(N__12152),
            .I(N__12149));
    LocalMux I__2941 (
            .O(N__12149),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2940 (
            .O(N__12146),
            .I(N__12143));
    LocalMux I__2939 (
            .O(N__12143),
            .I(N__12140));
    Span4Mux_v I__2938 (
            .O(N__12140),
            .I(N__12137));
    Odrv4 I__2937 (
            .O(N__12137),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    InMux I__2936 (
            .O(N__12134),
            .I(N__12131));
    LocalMux I__2935 (
            .O(N__12131),
            .I(N__12089));
    ClkMux I__2934 (
            .O(N__12130),
            .I(N__11975));
    ClkMux I__2933 (
            .O(N__12129),
            .I(N__11975));
    ClkMux I__2932 (
            .O(N__12128),
            .I(N__11975));
    ClkMux I__2931 (
            .O(N__12127),
            .I(N__11975));
    ClkMux I__2930 (
            .O(N__12126),
            .I(N__11975));
    ClkMux I__2929 (
            .O(N__12125),
            .I(N__11975));
    ClkMux I__2928 (
            .O(N__12124),
            .I(N__11975));
    ClkMux I__2927 (
            .O(N__12123),
            .I(N__11975));
    ClkMux I__2926 (
            .O(N__12122),
            .I(N__11975));
    ClkMux I__2925 (
            .O(N__12121),
            .I(N__11975));
    ClkMux I__2924 (
            .O(N__12120),
            .I(N__11975));
    ClkMux I__2923 (
            .O(N__12119),
            .I(N__11975));
    ClkMux I__2922 (
            .O(N__12118),
            .I(N__11975));
    ClkMux I__2921 (
            .O(N__12117),
            .I(N__11975));
    ClkMux I__2920 (
            .O(N__12116),
            .I(N__11975));
    ClkMux I__2919 (
            .O(N__12115),
            .I(N__11975));
    ClkMux I__2918 (
            .O(N__12114),
            .I(N__11975));
    ClkMux I__2917 (
            .O(N__12113),
            .I(N__11975));
    ClkMux I__2916 (
            .O(N__12112),
            .I(N__11975));
    ClkMux I__2915 (
            .O(N__12111),
            .I(N__11975));
    ClkMux I__2914 (
            .O(N__12110),
            .I(N__11975));
    ClkMux I__2913 (
            .O(N__12109),
            .I(N__11975));
    ClkMux I__2912 (
            .O(N__12108),
            .I(N__11975));
    ClkMux I__2911 (
            .O(N__12107),
            .I(N__11975));
    ClkMux I__2910 (
            .O(N__12106),
            .I(N__11975));
    ClkMux I__2909 (
            .O(N__12105),
            .I(N__11975));
    ClkMux I__2908 (
            .O(N__12104),
            .I(N__11975));
    ClkMux I__2907 (
            .O(N__12103),
            .I(N__11975));
    ClkMux I__2906 (
            .O(N__12102),
            .I(N__11975));
    ClkMux I__2905 (
            .O(N__12101),
            .I(N__11975));
    ClkMux I__2904 (
            .O(N__12100),
            .I(N__11975));
    ClkMux I__2903 (
            .O(N__12099),
            .I(N__11975));
    ClkMux I__2902 (
            .O(N__12098),
            .I(N__11975));
    ClkMux I__2901 (
            .O(N__12097),
            .I(N__11975));
    ClkMux I__2900 (
            .O(N__12096),
            .I(N__11975));
    ClkMux I__2899 (
            .O(N__12095),
            .I(N__11975));
    ClkMux I__2898 (
            .O(N__12094),
            .I(N__11975));
    ClkMux I__2897 (
            .O(N__12093),
            .I(N__11975));
    ClkMux I__2896 (
            .O(N__12092),
            .I(N__11975));
    Glb2LocalMux I__2895 (
            .O(N__12089),
            .I(N__11975));
    ClkMux I__2894 (
            .O(N__12088),
            .I(N__11975));
    ClkMux I__2893 (
            .O(N__12087),
            .I(N__11975));
    ClkMux I__2892 (
            .O(N__12086),
            .I(N__11975));
    ClkMux I__2891 (
            .O(N__12085),
            .I(N__11975));
    ClkMux I__2890 (
            .O(N__12084),
            .I(N__11975));
    ClkMux I__2889 (
            .O(N__12083),
            .I(N__11975));
    ClkMux I__2888 (
            .O(N__12082),
            .I(N__11975));
    ClkMux I__2887 (
            .O(N__12081),
            .I(N__11975));
    ClkMux I__2886 (
            .O(N__12080),
            .I(N__11975));
    ClkMux I__2885 (
            .O(N__12079),
            .I(N__11975));
    ClkMux I__2884 (
            .O(N__12078),
            .I(N__11975));
    GlobalMux I__2883 (
            .O(N__11975),
            .I(CLK80_PLL));
    InMux I__2882 (
            .O(N__11972),
            .I(N__11968));
    InMux I__2881 (
            .O(N__11971),
            .I(N__11965));
    LocalMux I__2880 (
            .O(N__11968),
            .I(N__11962));
    LocalMux I__2879 (
            .O(N__11965),
            .I(N__11959));
    Span4Mux_v I__2878 (
            .O(N__11962),
            .I(N__11956));
    Span4Mux_v I__2877 (
            .O(N__11959),
            .I(N__11953));
    Sp12to4 I__2876 (
            .O(N__11956),
            .I(N__11948));
    Sp12to4 I__2875 (
            .O(N__11953),
            .I(N__11948));
    Span12Mux_h I__2874 (
            .O(N__11948),
            .I(N__11945));
    Span12Mux_v I__2873 (
            .O(N__11945),
            .I(N__11942));
    Odrv12 I__2872 (
            .O(N__11942),
            .I(DRA_c_0));
    CascadeMux I__2871 (
            .O(N__11939),
            .I(N__11936));
    InMux I__2870 (
            .O(N__11936),
            .I(N__11933));
    LocalMux I__2869 (
            .O(N__11933),
            .I(N__11930));
    Span4Mux_v I__2868 (
            .O(N__11930),
            .I(N__11920));
    InMux I__2867 (
            .O(N__11929),
            .I(N__11913));
    InMux I__2866 (
            .O(N__11928),
            .I(N__11913));
    InMux I__2865 (
            .O(N__11927),
            .I(N__11910));
    InMux I__2864 (
            .O(N__11926),
            .I(N__11907));
    CascadeMux I__2863 (
            .O(N__11925),
            .I(N__11904));
    InMux I__2862 (
            .O(N__11924),
            .I(N__11899));
    CascadeMux I__2861 (
            .O(N__11923),
            .I(N__11896));
    Span4Mux_h I__2860 (
            .O(N__11920),
            .I(N__11889));
    InMux I__2859 (
            .O(N__11919),
            .I(N__11886));
    InMux I__2858 (
            .O(N__11918),
            .I(N__11883));
    LocalMux I__2857 (
            .O(N__11913),
            .I(N__11876));
    LocalMux I__2856 (
            .O(N__11910),
            .I(N__11876));
    LocalMux I__2855 (
            .O(N__11907),
            .I(N__11876));
    InMux I__2854 (
            .O(N__11904),
            .I(N__11871));
    InMux I__2853 (
            .O(N__11903),
            .I(N__11871));
    InMux I__2852 (
            .O(N__11902),
            .I(N__11866));
    LocalMux I__2851 (
            .O(N__11899),
            .I(N__11863));
    InMux I__2850 (
            .O(N__11896),
            .I(N__11858));
    InMux I__2849 (
            .O(N__11895),
            .I(N__11858));
    InMux I__2848 (
            .O(N__11894),
            .I(N__11855));
    InMux I__2847 (
            .O(N__11893),
            .I(N__11852));
    InMux I__2846 (
            .O(N__11892),
            .I(N__11849));
    Span4Mux_h I__2845 (
            .O(N__11889),
            .I(N__11840));
    LocalMux I__2844 (
            .O(N__11886),
            .I(N__11840));
    LocalMux I__2843 (
            .O(N__11883),
            .I(N__11840));
    Span4Mux_v I__2842 (
            .O(N__11876),
            .I(N__11840));
    LocalMux I__2841 (
            .O(N__11871),
            .I(N__11837));
    InMux I__2840 (
            .O(N__11870),
            .I(N__11834));
    InMux I__2839 (
            .O(N__11869),
            .I(N__11831));
    LocalMux I__2838 (
            .O(N__11866),
            .I(N__11818));
    Span4Mux_h I__2837 (
            .O(N__11863),
            .I(N__11818));
    LocalMux I__2836 (
            .O(N__11858),
            .I(N__11818));
    LocalMux I__2835 (
            .O(N__11855),
            .I(N__11818));
    LocalMux I__2834 (
            .O(N__11852),
            .I(N__11818));
    LocalMux I__2833 (
            .O(N__11849),
            .I(N__11818));
    Span4Mux_h I__2832 (
            .O(N__11840),
            .I(N__11810));
    Span4Mux_v I__2831 (
            .O(N__11837),
            .I(N__11810));
    LocalMux I__2830 (
            .O(N__11834),
            .I(N__11803));
    LocalMux I__2829 (
            .O(N__11831),
            .I(N__11803));
    Span4Mux_v I__2828 (
            .O(N__11818),
            .I(N__11803));
    InMux I__2827 (
            .O(N__11817),
            .I(N__11798));
    InMux I__2826 (
            .O(N__11816),
            .I(N__11798));
    InMux I__2825 (
            .O(N__11815),
            .I(N__11795));
    Sp12to4 I__2824 (
            .O(N__11810),
            .I(N__11790));
    Sp12to4 I__2823 (
            .O(N__11803),
            .I(N__11790));
    LocalMux I__2822 (
            .O(N__11798),
            .I(N__11785));
    LocalMux I__2821 (
            .O(N__11795),
            .I(N__11785));
    Span12Mux_h I__2820 (
            .O(N__11790),
            .I(N__11782));
    Span12Mux_h I__2819 (
            .O(N__11785),
            .I(N__11779));
    Span12Mux_v I__2818 (
            .O(N__11782),
            .I(N__11776));
    Span12Mux_v I__2817 (
            .O(N__11779),
            .I(N__11773));
    Odrv12 I__2816 (
            .O(N__11776),
            .I(AGNUS_REV_c));
    Odrv12 I__2815 (
            .O(N__11773),
            .I(AGNUS_REV_c));
    InMux I__2814 (
            .O(N__11768),
            .I(N__11765));
    LocalMux I__2813 (
            .O(N__11765),
            .I(N__11760));
    InMux I__2812 (
            .O(N__11764),
            .I(N__11755));
    InMux I__2811 (
            .O(N__11763),
            .I(N__11755));
    Span4Mux_v I__2810 (
            .O(N__11760),
            .I(N__11749));
    LocalMux I__2809 (
            .O(N__11755),
            .I(N__11749));
    InMux I__2808 (
            .O(N__11754),
            .I(N__11746));
    Sp12to4 I__2807 (
            .O(N__11749),
            .I(N__11741));
    LocalMux I__2806 (
            .O(N__11746),
            .I(N__11741));
    Span12Mux_v I__2805 (
            .O(N__11741),
            .I(N__11738));
    Odrv12 I__2804 (
            .O(N__11738),
            .I(DRA_c_1));
    InMux I__2803 (
            .O(N__11735),
            .I(N__11732));
    LocalMux I__2802 (
            .O(N__11732),
            .I(N__11729));
    Span12Mux_v I__2801 (
            .O(N__11729),
            .I(N__11726));
    Odrv12 I__2800 (
            .O(N__11726),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    ClkMux I__2799 (
            .O(N__11723),
            .I(N__11702));
    ClkMux I__2798 (
            .O(N__11722),
            .I(N__11702));
    ClkMux I__2797 (
            .O(N__11721),
            .I(N__11702));
    ClkMux I__2796 (
            .O(N__11720),
            .I(N__11702));
    ClkMux I__2795 (
            .O(N__11719),
            .I(N__11702));
    ClkMux I__2794 (
            .O(N__11718),
            .I(N__11702));
    ClkMux I__2793 (
            .O(N__11717),
            .I(N__11702));
    GlobalMux I__2792 (
            .O(N__11702),
            .I(N__11699));
    gio2CtrlBuf I__2791 (
            .O(N__11699),
            .I(C3_c_g));
    CEMux I__2790 (
            .O(N__11696),
            .I(N__11651));
    CEMux I__2789 (
            .O(N__11695),
            .I(N__11651));
    CEMux I__2788 (
            .O(N__11694),
            .I(N__11651));
    CEMux I__2787 (
            .O(N__11693),
            .I(N__11651));
    CEMux I__2786 (
            .O(N__11692),
            .I(N__11651));
    CEMux I__2785 (
            .O(N__11691),
            .I(N__11651));
    CEMux I__2784 (
            .O(N__11690),
            .I(N__11651));
    CEMux I__2783 (
            .O(N__11689),
            .I(N__11651));
    CEMux I__2782 (
            .O(N__11688),
            .I(N__11651));
    CEMux I__2781 (
            .O(N__11687),
            .I(N__11651));
    CEMux I__2780 (
            .O(N__11686),
            .I(N__11651));
    CEMux I__2779 (
            .O(N__11685),
            .I(N__11651));
    CEMux I__2778 (
            .O(N__11684),
            .I(N__11651));
    CEMux I__2777 (
            .O(N__11683),
            .I(N__11651));
    CEMux I__2776 (
            .O(N__11682),
            .I(N__11651));
    GlobalMux I__2775 (
            .O(N__11651),
            .I(N__11648));
    gio2CtrlBuf I__2774 (
            .O(N__11648),
            .I(DBRn_c_i_0_g));
    InMux I__2773 (
            .O(N__11645),
            .I(N__11638));
    InMux I__2772 (
            .O(N__11644),
            .I(N__11635));
    InMux I__2771 (
            .O(N__11643),
            .I(N__11632));
    InMux I__2770 (
            .O(N__11642),
            .I(N__11629));
    InMux I__2769 (
            .O(N__11641),
            .I(N__11626));
    LocalMux I__2768 (
            .O(N__11638),
            .I(N__11612));
    LocalMux I__2767 (
            .O(N__11635),
            .I(N__11587));
    LocalMux I__2766 (
            .O(N__11632),
            .I(N__11581));
    LocalMux I__2765 (
            .O(N__11629),
            .I(N__11565));
    LocalMux I__2764 (
            .O(N__11626),
            .I(N__11559));
    SRMux I__2763 (
            .O(N__11625),
            .I(N__11435));
    SRMux I__2762 (
            .O(N__11624),
            .I(N__11435));
    SRMux I__2761 (
            .O(N__11623),
            .I(N__11435));
    SRMux I__2760 (
            .O(N__11622),
            .I(N__11435));
    SRMux I__2759 (
            .O(N__11621),
            .I(N__11435));
    SRMux I__2758 (
            .O(N__11620),
            .I(N__11435));
    SRMux I__2757 (
            .O(N__11619),
            .I(N__11435));
    SRMux I__2756 (
            .O(N__11618),
            .I(N__11435));
    SRMux I__2755 (
            .O(N__11617),
            .I(N__11435));
    SRMux I__2754 (
            .O(N__11616),
            .I(N__11435));
    SRMux I__2753 (
            .O(N__11615),
            .I(N__11435));
    Glb2LocalMux I__2752 (
            .O(N__11612),
            .I(N__11435));
    SRMux I__2751 (
            .O(N__11611),
            .I(N__11435));
    SRMux I__2750 (
            .O(N__11610),
            .I(N__11435));
    SRMux I__2749 (
            .O(N__11609),
            .I(N__11435));
    SRMux I__2748 (
            .O(N__11608),
            .I(N__11435));
    SRMux I__2747 (
            .O(N__11607),
            .I(N__11435));
    SRMux I__2746 (
            .O(N__11606),
            .I(N__11435));
    SRMux I__2745 (
            .O(N__11605),
            .I(N__11435));
    SRMux I__2744 (
            .O(N__11604),
            .I(N__11435));
    SRMux I__2743 (
            .O(N__11603),
            .I(N__11435));
    SRMux I__2742 (
            .O(N__11602),
            .I(N__11435));
    SRMux I__2741 (
            .O(N__11601),
            .I(N__11435));
    SRMux I__2740 (
            .O(N__11600),
            .I(N__11435));
    SRMux I__2739 (
            .O(N__11599),
            .I(N__11435));
    SRMux I__2738 (
            .O(N__11598),
            .I(N__11435));
    SRMux I__2737 (
            .O(N__11597),
            .I(N__11435));
    SRMux I__2736 (
            .O(N__11596),
            .I(N__11435));
    SRMux I__2735 (
            .O(N__11595),
            .I(N__11435));
    SRMux I__2734 (
            .O(N__11594),
            .I(N__11435));
    SRMux I__2733 (
            .O(N__11593),
            .I(N__11435));
    SRMux I__2732 (
            .O(N__11592),
            .I(N__11435));
    SRMux I__2731 (
            .O(N__11591),
            .I(N__11435));
    SRMux I__2730 (
            .O(N__11590),
            .I(N__11435));
    Glb2LocalMux I__2729 (
            .O(N__11587),
            .I(N__11435));
    SRMux I__2728 (
            .O(N__11586),
            .I(N__11435));
    SRMux I__2727 (
            .O(N__11585),
            .I(N__11435));
    SRMux I__2726 (
            .O(N__11584),
            .I(N__11435));
    Glb2LocalMux I__2725 (
            .O(N__11581),
            .I(N__11435));
    SRMux I__2724 (
            .O(N__11580),
            .I(N__11435));
    SRMux I__2723 (
            .O(N__11579),
            .I(N__11435));
    SRMux I__2722 (
            .O(N__11578),
            .I(N__11435));
    SRMux I__2721 (
            .O(N__11577),
            .I(N__11435));
    SRMux I__2720 (
            .O(N__11576),
            .I(N__11435));
    SRMux I__2719 (
            .O(N__11575),
            .I(N__11435));
    SRMux I__2718 (
            .O(N__11574),
            .I(N__11435));
    SRMux I__2717 (
            .O(N__11573),
            .I(N__11435));
    SRMux I__2716 (
            .O(N__11572),
            .I(N__11435));
    SRMux I__2715 (
            .O(N__11571),
            .I(N__11435));
    SRMux I__2714 (
            .O(N__11570),
            .I(N__11435));
    SRMux I__2713 (
            .O(N__11569),
            .I(N__11435));
    SRMux I__2712 (
            .O(N__11568),
            .I(N__11435));
    Glb2LocalMux I__2711 (
            .O(N__11565),
            .I(N__11435));
    SRMux I__2710 (
            .O(N__11564),
            .I(N__11435));
    SRMux I__2709 (
            .O(N__11563),
            .I(N__11435));
    SRMux I__2708 (
            .O(N__11562),
            .I(N__11435));
    Glb2LocalMux I__2707 (
            .O(N__11559),
            .I(N__11435));
    SRMux I__2706 (
            .O(N__11558),
            .I(N__11435));
    SRMux I__2705 (
            .O(N__11557),
            .I(N__11435));
    SRMux I__2704 (
            .O(N__11556),
            .I(N__11435));
    GlobalMux I__2703 (
            .O(N__11435),
            .I(N__11432));
    gio2CtrlBuf I__2702 (
            .O(N__11432),
            .I(RESETn_c_i_g));
    CascadeMux I__2701 (
            .O(N__11429),
            .I(N__11426));
    InMux I__2700 (
            .O(N__11426),
            .I(N__11421));
    InMux I__2699 (
            .O(N__11425),
            .I(N__11418));
    InMux I__2698 (
            .O(N__11424),
            .I(N__11415));
    LocalMux I__2697 (
            .O(N__11421),
            .I(N__11412));
    LocalMux I__2696 (
            .O(N__11418),
            .I(N__11408));
    LocalMux I__2695 (
            .O(N__11415),
            .I(N__11405));
    Span4Mux_v I__2694 (
            .O(N__11412),
            .I(N__11402));
    InMux I__2693 (
            .O(N__11411),
            .I(N__11399));
    Span4Mux_v I__2692 (
            .O(N__11408),
            .I(N__11395));
    Span4Mux_v I__2691 (
            .O(N__11405),
            .I(N__11392));
    Span4Mux_v I__2690 (
            .O(N__11402),
            .I(N__11389));
    LocalMux I__2689 (
            .O(N__11399),
            .I(N__11386));
    InMux I__2688 (
            .O(N__11398),
            .I(N__11383));
    Sp12to4 I__2687 (
            .O(N__11395),
            .I(N__11378));
    Sp12to4 I__2686 (
            .O(N__11392),
            .I(N__11378));
    Sp12to4 I__2685 (
            .O(N__11389),
            .I(N__11375));
    Sp12to4 I__2684 (
            .O(N__11386),
            .I(N__11370));
    LocalMux I__2683 (
            .O(N__11383),
            .I(N__11370));
    Span12Mux_h I__2682 (
            .O(N__11378),
            .I(N__11367));
    Span12Mux_h I__2681 (
            .O(N__11375),
            .I(N__11362));
    Span12Mux_v I__2680 (
            .O(N__11370),
            .I(N__11362));
    Span12Mux_v I__2679 (
            .O(N__11367),
            .I(N__11357));
    Span12Mux_h I__2678 (
            .O(N__11362),
            .I(N__11357));
    Odrv12 I__2677 (
            .O(N__11357),
            .I(RnW_c));
    InMux I__2676 (
            .O(N__11354),
            .I(N__11350));
    InMux I__2675 (
            .O(N__11353),
            .I(N__11347));
    LocalMux I__2674 (
            .O(N__11350),
            .I(N__11344));
    LocalMux I__2673 (
            .O(N__11347),
            .I(N__11341));
    Span4Mux_v I__2672 (
            .O(N__11344),
            .I(N__11338));
    Span12Mux_v I__2671 (
            .O(N__11341),
            .I(N__11335));
    Span4Mux_h I__2670 (
            .O(N__11338),
            .I(N__11332));
    Span12Mux_h I__2669 (
            .O(N__11335),
            .I(N__11328));
    Span4Mux_h I__2668 (
            .O(N__11332),
            .I(N__11325));
    InMux I__2667 (
            .O(N__11331),
            .I(N__11322));
    Odrv12 I__2666 (
            .O(N__11328),
            .I(\U712_CHIP_RAM.DMA_WRITE_CYCLEZ0 ));
    Odrv4 I__2665 (
            .O(N__11325),
            .I(\U712_CHIP_RAM.DMA_WRITE_CYCLEZ0 ));
    LocalMux I__2664 (
            .O(N__11322),
            .I(\U712_CHIP_RAM.DMA_WRITE_CYCLEZ0 ));
    IoInMux I__2663 (
            .O(N__11315),
            .I(N__11312));
    LocalMux I__2662 (
            .O(N__11312),
            .I(N__11309));
    IoSpan4Mux I__2661 (
            .O(N__11309),
            .I(N__11306));
    Span4Mux_s3_h I__2660 (
            .O(N__11306),
            .I(N__11303));
    Odrv4 I__2659 (
            .O(N__11303),
            .I(N_323_mux));
    InMux I__2658 (
            .O(N__11300),
            .I(N__11297));
    LocalMux I__2657 (
            .O(N__11297),
            .I(N__11294));
    Span4Mux_v I__2656 (
            .O(N__11294),
            .I(N__11290));
    InMux I__2655 (
            .O(N__11293),
            .I(N__11287));
    Span4Mux_v I__2654 (
            .O(N__11290),
            .I(N__11281));
    LocalMux I__2653 (
            .O(N__11287),
            .I(N__11281));
    InMux I__2652 (
            .O(N__11286),
            .I(N__11276));
    Span4Mux_v I__2651 (
            .O(N__11281),
            .I(N__11273));
    InMux I__2650 (
            .O(N__11280),
            .I(N__11268));
    InMux I__2649 (
            .O(N__11279),
            .I(N__11268));
    LocalMux I__2648 (
            .O(N__11276),
            .I(N__11265));
    Span4Mux_v I__2647 (
            .O(N__11273),
            .I(N__11262));
    LocalMux I__2646 (
            .O(N__11268),
            .I(N__11259));
    Span12Mux_h I__2645 (
            .O(N__11265),
            .I(N__11256));
    Sp12to4 I__2644 (
            .O(N__11262),
            .I(N__11253));
    Span4Mux_v I__2643 (
            .O(N__11259),
            .I(N__11250));
    Span12Mux_v I__2642 (
            .O(N__11256),
            .I(N__11247));
    Span12Mux_h I__2641 (
            .O(N__11253),
            .I(N__11244));
    Span4Mux_v I__2640 (
            .O(N__11250),
            .I(N__11241));
    Odrv12 I__2639 (
            .O(N__11247),
            .I(CASLn_c));
    Odrv12 I__2638 (
            .O(N__11244),
            .I(CASLn_c));
    Odrv4 I__2637 (
            .O(N__11241),
            .I(CASLn_c));
    InMux I__2636 (
            .O(N__11234),
            .I(N__11231));
    LocalMux I__2635 (
            .O(N__11231),
            .I(N__11228));
    Span4Mux_v I__2634 (
            .O(N__11228),
            .I(N__11225));
    Span4Mux_v I__2633 (
            .O(N__11225),
            .I(N__11220));
    InMux I__2632 (
            .O(N__11224),
            .I(N__11215));
    InMux I__2631 (
            .O(N__11223),
            .I(N__11212));
    Span4Mux_h I__2630 (
            .O(N__11220),
            .I(N__11209));
    InMux I__2629 (
            .O(N__11219),
            .I(N__11204));
    InMux I__2628 (
            .O(N__11218),
            .I(N__11204));
    LocalMux I__2627 (
            .O(N__11215),
            .I(N__11199));
    LocalMux I__2626 (
            .O(N__11212),
            .I(N__11199));
    Span4Mux_h I__2625 (
            .O(N__11209),
            .I(N__11194));
    LocalMux I__2624 (
            .O(N__11204),
            .I(N__11194));
    Span12Mux_v I__2623 (
            .O(N__11199),
            .I(N__11191));
    Span4Mux_h I__2622 (
            .O(N__11194),
            .I(N__11188));
    Span12Mux_h I__2621 (
            .O(N__11191),
            .I(N__11185));
    Span4Mux_v I__2620 (
            .O(N__11188),
            .I(N__11182));
    Odrv12 I__2619 (
            .O(N__11185),
            .I(CASUn_c));
    Odrv4 I__2618 (
            .O(N__11182),
            .I(CASUn_c));
    CascadeMux I__2617 (
            .O(N__11177),
            .I(N__11174));
    InMux I__2616 (
            .O(N__11174),
            .I(N__11171));
    LocalMux I__2615 (
            .O(N__11171),
            .I(N__11167));
    InMux I__2614 (
            .O(N__11170),
            .I(N__11164));
    Span4Mux_v I__2613 (
            .O(N__11167),
            .I(N__11161));
    LocalMux I__2612 (
            .O(N__11164),
            .I(N__11158));
    Span4Mux_v I__2611 (
            .O(N__11161),
            .I(N__11155));
    Span4Mux_v I__2610 (
            .O(N__11158),
            .I(N__11152));
    Sp12to4 I__2609 (
            .O(N__11155),
            .I(N__11147));
    Span4Mux_v I__2608 (
            .O(N__11152),
            .I(N__11144));
    InMux I__2607 (
            .O(N__11151),
            .I(N__11139));
    InMux I__2606 (
            .O(N__11150),
            .I(N__11139));
    Odrv12 I__2605 (
            .O(N__11147),
            .I(REG_CYCLEm));
    Odrv4 I__2604 (
            .O(N__11144),
            .I(REG_CYCLEm));
    LocalMux I__2603 (
            .O(N__11139),
            .I(REG_CYCLEm));
    InMux I__2602 (
            .O(N__11132),
            .I(N__11126));
    CascadeMux I__2601 (
            .O(N__11131),
            .I(N__11120));
    CascadeMux I__2600 (
            .O(N__11130),
            .I(N__11116));
    CascadeMux I__2599 (
            .O(N__11129),
            .I(N__11109));
    LocalMux I__2598 (
            .O(N__11126),
            .I(N__11105));
    CascadeMux I__2597 (
            .O(N__11125),
            .I(N__11097));
    InMux I__2596 (
            .O(N__11124),
            .I(N__11090));
    InMux I__2595 (
            .O(N__11123),
            .I(N__11085));
    InMux I__2594 (
            .O(N__11120),
            .I(N__11085));
    CascadeMux I__2593 (
            .O(N__11119),
            .I(N__11082));
    InMux I__2592 (
            .O(N__11116),
            .I(N__11077));
    InMux I__2591 (
            .O(N__11115),
            .I(N__11077));
    InMux I__2590 (
            .O(N__11114),
            .I(N__11072));
    InMux I__2589 (
            .O(N__11113),
            .I(N__11072));
    InMux I__2588 (
            .O(N__11112),
            .I(N__11067));
    InMux I__2587 (
            .O(N__11109),
            .I(N__11067));
    CascadeMux I__2586 (
            .O(N__11108),
            .I(N__11062));
    Span4Mux_v I__2585 (
            .O(N__11105),
            .I(N__11059));
    CascadeMux I__2584 (
            .O(N__11104),
            .I(N__11055));
    CascadeMux I__2583 (
            .O(N__11103),
            .I(N__11052));
    CascadeMux I__2582 (
            .O(N__11102),
            .I(N__11049));
    CascadeMux I__2581 (
            .O(N__11101),
            .I(N__11045));
    InMux I__2580 (
            .O(N__11100),
            .I(N__11041));
    InMux I__2579 (
            .O(N__11097),
            .I(N__11038));
    InMux I__2578 (
            .O(N__11096),
            .I(N__11033));
    InMux I__2577 (
            .O(N__11095),
            .I(N__11033));
    InMux I__2576 (
            .O(N__11094),
            .I(N__11028));
    InMux I__2575 (
            .O(N__11093),
            .I(N__11028));
    LocalMux I__2574 (
            .O(N__11090),
            .I(N__11025));
    LocalMux I__2573 (
            .O(N__11085),
            .I(N__11022));
    InMux I__2572 (
            .O(N__11082),
            .I(N__11019));
    LocalMux I__2571 (
            .O(N__11077),
            .I(N__11012));
    LocalMux I__2570 (
            .O(N__11072),
            .I(N__11012));
    LocalMux I__2569 (
            .O(N__11067),
            .I(N__11012));
    InMux I__2568 (
            .O(N__11066),
            .I(N__11005));
    InMux I__2567 (
            .O(N__11065),
            .I(N__11005));
    InMux I__2566 (
            .O(N__11062),
            .I(N__11005));
    Sp12to4 I__2565 (
            .O(N__11059),
            .I(N__11002));
    CascadeMux I__2564 (
            .O(N__11058),
            .I(N__10998));
    InMux I__2563 (
            .O(N__11055),
            .I(N__10989));
    InMux I__2562 (
            .O(N__11052),
            .I(N__10986));
    InMux I__2561 (
            .O(N__11049),
            .I(N__10983));
    InMux I__2560 (
            .O(N__11048),
            .I(N__10980));
    InMux I__2559 (
            .O(N__11045),
            .I(N__10977));
    InMux I__2558 (
            .O(N__11044),
            .I(N__10974));
    LocalMux I__2557 (
            .O(N__11041),
            .I(N__10970));
    LocalMux I__2556 (
            .O(N__11038),
            .I(N__10963));
    LocalMux I__2555 (
            .O(N__11033),
            .I(N__10963));
    LocalMux I__2554 (
            .O(N__11028),
            .I(N__10963));
    Span4Mux_h I__2553 (
            .O(N__11025),
            .I(N__10948));
    Span4Mux_h I__2552 (
            .O(N__11022),
            .I(N__10948));
    LocalMux I__2551 (
            .O(N__11019),
            .I(N__10948));
    Span4Mux_v I__2550 (
            .O(N__11012),
            .I(N__10948));
    LocalMux I__2549 (
            .O(N__11005),
            .I(N__10948));
    Span12Mux_s11_h I__2548 (
            .O(N__11002),
            .I(N__10945));
    InMux I__2547 (
            .O(N__11001),
            .I(N__10942));
    InMux I__2546 (
            .O(N__10998),
            .I(N__10939));
    InMux I__2545 (
            .O(N__10997),
            .I(N__10934));
    InMux I__2544 (
            .O(N__10996),
            .I(N__10934));
    InMux I__2543 (
            .O(N__10995),
            .I(N__10931));
    InMux I__2542 (
            .O(N__10994),
            .I(N__10928));
    InMux I__2541 (
            .O(N__10993),
            .I(N__10925));
    InMux I__2540 (
            .O(N__10992),
            .I(N__10922));
    LocalMux I__2539 (
            .O(N__10989),
            .I(N__10911));
    LocalMux I__2538 (
            .O(N__10986),
            .I(N__10911));
    LocalMux I__2537 (
            .O(N__10983),
            .I(N__10911));
    LocalMux I__2536 (
            .O(N__10980),
            .I(N__10911));
    LocalMux I__2535 (
            .O(N__10977),
            .I(N__10911));
    LocalMux I__2534 (
            .O(N__10974),
            .I(N__10908));
    InMux I__2533 (
            .O(N__10973),
            .I(N__10905));
    Span4Mux_v I__2532 (
            .O(N__10970),
            .I(N__10900));
    Span4Mux_v I__2531 (
            .O(N__10963),
            .I(N__10900));
    InMux I__2530 (
            .O(N__10962),
            .I(N__10891));
    InMux I__2529 (
            .O(N__10961),
            .I(N__10891));
    InMux I__2528 (
            .O(N__10960),
            .I(N__10891));
    InMux I__2527 (
            .O(N__10959),
            .I(N__10891));
    Span4Mux_h I__2526 (
            .O(N__10948),
            .I(N__10888));
    Span12Mux_v I__2525 (
            .O(N__10945),
            .I(N__10873));
    LocalMux I__2524 (
            .O(N__10942),
            .I(N__10873));
    LocalMux I__2523 (
            .O(N__10939),
            .I(N__10873));
    LocalMux I__2522 (
            .O(N__10934),
            .I(N__10873));
    LocalMux I__2521 (
            .O(N__10931),
            .I(N__10873));
    LocalMux I__2520 (
            .O(N__10928),
            .I(N__10873));
    LocalMux I__2519 (
            .O(N__10925),
            .I(N__10873));
    LocalMux I__2518 (
            .O(N__10922),
            .I(N__10868));
    Span12Mux_h I__2517 (
            .O(N__10911),
            .I(N__10868));
    Odrv4 I__2516 (
            .O(N__10908),
            .I(\U712_CHIP_RAM.CPU_CYCLEm ));
    LocalMux I__2515 (
            .O(N__10905),
            .I(\U712_CHIP_RAM.CPU_CYCLEm ));
    Odrv4 I__2514 (
            .O(N__10900),
            .I(\U712_CHIP_RAM.CPU_CYCLEm ));
    LocalMux I__2513 (
            .O(N__10891),
            .I(\U712_CHIP_RAM.CPU_CYCLEm ));
    Odrv4 I__2512 (
            .O(N__10888),
            .I(\U712_CHIP_RAM.CPU_CYCLEm ));
    Odrv12 I__2511 (
            .O(N__10873),
            .I(\U712_CHIP_RAM.CPU_CYCLEm ));
    Odrv12 I__2510 (
            .O(N__10868),
            .I(\U712_CHIP_RAM.CPU_CYCLEm ));
    IoInMux I__2509 (
            .O(N__10853),
            .I(N__10850));
    LocalMux I__2508 (
            .O(N__10850),
            .I(N__10847));
    Span4Mux_s3_v I__2507 (
            .O(N__10847),
            .I(N__10844));
    Span4Mux_v I__2506 (
            .O(N__10844),
            .I(N__10841));
    Odrv4 I__2505 (
            .O(N__10841),
            .I(N_333_mux));
    InMux I__2504 (
            .O(N__10838),
            .I(N__10834));
    InMux I__2503 (
            .O(N__10837),
            .I(N__10830));
    LocalMux I__2502 (
            .O(N__10834),
            .I(N__10826));
    InMux I__2501 (
            .O(N__10833),
            .I(N__10823));
    LocalMux I__2500 (
            .O(N__10830),
            .I(N__10820));
    InMux I__2499 (
            .O(N__10829),
            .I(N__10817));
    Span4Mux_h I__2498 (
            .O(N__10826),
            .I(N__10814));
    LocalMux I__2497 (
            .O(N__10823),
            .I(N__10811));
    Span4Mux_v I__2496 (
            .O(N__10820),
            .I(N__10806));
    LocalMux I__2495 (
            .O(N__10817),
            .I(N__10806));
    Span4Mux_v I__2494 (
            .O(N__10814),
            .I(N__10803));
    Span4Mux_v I__2493 (
            .O(N__10811),
            .I(N__10798));
    Span4Mux_h I__2492 (
            .O(N__10806),
            .I(N__10798));
    Sp12to4 I__2491 (
            .O(N__10803),
            .I(N__10793));
    Sp12to4 I__2490 (
            .O(N__10798),
            .I(N__10793));
    Span12Mux_v I__2489 (
            .O(N__10793),
            .I(N__10790));
    Odrv12 I__2488 (
            .O(N__10790),
            .I(DRA_c_9));
    InMux I__2487 (
            .O(N__10787),
            .I(N__10784));
    LocalMux I__2486 (
            .O(N__10784),
            .I(N__10781));
    Span4Mux_h I__2485 (
            .O(N__10781),
            .I(N__10778));
    Odrv4 I__2484 (
            .O(N__10778),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    InMux I__2483 (
            .O(N__10775),
            .I(N__10772));
    LocalMux I__2482 (
            .O(N__10772),
            .I(N__10769));
    Odrv4 I__2481 (
            .O(N__10769),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2480 (
            .O(N__10766),
            .I(N__10763));
    LocalMux I__2479 (
            .O(N__10763),
            .I(N__10760));
    Span4Mux_v I__2478 (
            .O(N__10760),
            .I(N__10757));
    Span4Mux_h I__2477 (
            .O(N__10757),
            .I(N__10754));
    Odrv4 I__2476 (
            .O(N__10754),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2475 (
            .O(N__10751),
            .I(N__10746));
    InMux I__2474 (
            .O(N__10750),
            .I(N__10743));
    InMux I__2473 (
            .O(N__10749),
            .I(N__10740));
    LocalMux I__2472 (
            .O(N__10746),
            .I(N__10736));
    LocalMux I__2471 (
            .O(N__10743),
            .I(N__10731));
    LocalMux I__2470 (
            .O(N__10740),
            .I(N__10731));
    InMux I__2469 (
            .O(N__10739),
            .I(N__10728));
    Span4Mux_h I__2468 (
            .O(N__10736),
            .I(N__10725));
    Span4Mux_h I__2467 (
            .O(N__10731),
            .I(N__10720));
    LocalMux I__2466 (
            .O(N__10728),
            .I(N__10720));
    Span4Mux_v I__2465 (
            .O(N__10725),
            .I(N__10717));
    Sp12to4 I__2464 (
            .O(N__10720),
            .I(N__10714));
    Sp12to4 I__2463 (
            .O(N__10717),
            .I(N__10709));
    Span12Mux_v I__2462 (
            .O(N__10714),
            .I(N__10709));
    Odrv12 I__2461 (
            .O(N__10709),
            .I(DRA_c_5));
    InMux I__2460 (
            .O(N__10706),
            .I(N__10703));
    LocalMux I__2459 (
            .O(N__10703),
            .I(N__10700));
    Span4Mux_h I__2458 (
            .O(N__10700),
            .I(N__10697));
    Odrv4 I__2457 (
            .O(N__10697),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__2456 (
            .O(N__10694),
            .I(N__10691));
    LocalMux I__2455 (
            .O(N__10691),
            .I(N__10688));
    Span4Mux_h I__2454 (
            .O(N__10688),
            .I(N__10685));
    Span4Mux_h I__2453 (
            .O(N__10685),
            .I(N__10682));
    Odrv4 I__2452 (
            .O(N__10682),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__2451 (
            .O(N__10679),
            .I(N__10676));
    LocalMux I__2450 (
            .O(N__10676),
            .I(N__10673));
    Span4Mux_h I__2449 (
            .O(N__10673),
            .I(N__10670));
    Span4Mux_h I__2448 (
            .O(N__10670),
            .I(N__10667));
    Odrv4 I__2447 (
            .O(N__10667),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__2446 (
            .O(N__10664),
            .I(N__10661));
    LocalMux I__2445 (
            .O(N__10661),
            .I(N__10658));
    Span4Mux_v I__2444 (
            .O(N__10658),
            .I(N__10654));
    InMux I__2443 (
            .O(N__10657),
            .I(N__10651));
    Span4Mux_v I__2442 (
            .O(N__10654),
            .I(N__10646));
    LocalMux I__2441 (
            .O(N__10651),
            .I(N__10646));
    Span4Mux_h I__2440 (
            .O(N__10646),
            .I(N__10640));
    CascadeMux I__2439 (
            .O(N__10645),
            .I(N__10637));
    InMux I__2438 (
            .O(N__10644),
            .I(N__10634));
    InMux I__2437 (
            .O(N__10643),
            .I(N__10631));
    Span4Mux_h I__2436 (
            .O(N__10640),
            .I(N__10628));
    InMux I__2435 (
            .O(N__10637),
            .I(N__10625));
    LocalMux I__2434 (
            .O(N__10634),
            .I(N__10622));
    LocalMux I__2433 (
            .O(N__10631),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__2432 (
            .O(N__10628),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__2431 (
            .O(N__10625),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv12 I__2430 (
            .O(N__10622),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__2429 (
            .O(N__10613),
            .I(N__10610));
    LocalMux I__2428 (
            .O(N__10610),
            .I(N__10607));
    IoSpan4Mux I__2427 (
            .O(N__10607),
            .I(N__10604));
    Span4Mux_s3_v I__2426 (
            .O(N__10604),
            .I(N__10601));
    Span4Mux_v I__2425 (
            .O(N__10601),
            .I(N__10598));
    Odrv4 I__2424 (
            .O(N__10598),
            .I(CRCSn_c));
    IoInMux I__2423 (
            .O(N__10595),
            .I(N__10592));
    LocalMux I__2422 (
            .O(N__10592),
            .I(N__10589));
    IoSpan4Mux I__2421 (
            .O(N__10589),
            .I(N__10586));
    Span4Mux_s2_v I__2420 (
            .O(N__10586),
            .I(N__10583));
    Span4Mux_v I__2419 (
            .O(N__10583),
            .I(N__10580));
    Span4Mux_v I__2418 (
            .O(N__10580),
            .I(N__10577));
    Odrv4 I__2417 (
            .O(N__10577),
            .I(CASn_c));
    CascadeMux I__2416 (
            .O(N__10574),
            .I(N__10564));
    InMux I__2415 (
            .O(N__10573),
            .I(N__10561));
    InMux I__2414 (
            .O(N__10572),
            .I(N__10558));
    CascadeMux I__2413 (
            .O(N__10571),
            .I(N__10554));
    CascadeMux I__2412 (
            .O(N__10570),
            .I(N__10550));
    InMux I__2411 (
            .O(N__10569),
            .I(N__10545));
    CascadeMux I__2410 (
            .O(N__10568),
            .I(N__10536));
    CascadeMux I__2409 (
            .O(N__10567),
            .I(N__10531));
    InMux I__2408 (
            .O(N__10564),
            .I(N__10527));
    LocalMux I__2407 (
            .O(N__10561),
            .I(N__10524));
    LocalMux I__2406 (
            .O(N__10558),
            .I(N__10521));
    InMux I__2405 (
            .O(N__10557),
            .I(N__10518));
    InMux I__2404 (
            .O(N__10554),
            .I(N__10512));
    InMux I__2403 (
            .O(N__10553),
            .I(N__10512));
    InMux I__2402 (
            .O(N__10550),
            .I(N__10505));
    InMux I__2401 (
            .O(N__10549),
            .I(N__10505));
    InMux I__2400 (
            .O(N__10548),
            .I(N__10505));
    LocalMux I__2399 (
            .O(N__10545),
            .I(N__10502));
    InMux I__2398 (
            .O(N__10544),
            .I(N__10497));
    InMux I__2397 (
            .O(N__10543),
            .I(N__10497));
    InMux I__2396 (
            .O(N__10542),
            .I(N__10492));
    InMux I__2395 (
            .O(N__10541),
            .I(N__10492));
    CascadeMux I__2394 (
            .O(N__10540),
            .I(N__10487));
    InMux I__2393 (
            .O(N__10539),
            .I(N__10484));
    InMux I__2392 (
            .O(N__10536),
            .I(N__10481));
    InMux I__2391 (
            .O(N__10535),
            .I(N__10476));
    InMux I__2390 (
            .O(N__10534),
            .I(N__10476));
    InMux I__2389 (
            .O(N__10531),
            .I(N__10471));
    InMux I__2388 (
            .O(N__10530),
            .I(N__10471));
    LocalMux I__2387 (
            .O(N__10527),
            .I(N__10462));
    Span4Mux_v I__2386 (
            .O(N__10524),
            .I(N__10462));
    Span4Mux_h I__2385 (
            .O(N__10521),
            .I(N__10462));
    LocalMux I__2384 (
            .O(N__10518),
            .I(N__10462));
    InMux I__2383 (
            .O(N__10517),
            .I(N__10457));
    LocalMux I__2382 (
            .O(N__10512),
            .I(N__10452));
    LocalMux I__2381 (
            .O(N__10505),
            .I(N__10452));
    Span4Mux_h I__2380 (
            .O(N__10502),
            .I(N__10443));
    LocalMux I__2379 (
            .O(N__10497),
            .I(N__10443));
    LocalMux I__2378 (
            .O(N__10492),
            .I(N__10443));
    InMux I__2377 (
            .O(N__10491),
            .I(N__10436));
    InMux I__2376 (
            .O(N__10490),
            .I(N__10433));
    InMux I__2375 (
            .O(N__10487),
            .I(N__10430));
    LocalMux I__2374 (
            .O(N__10484),
            .I(N__10425));
    LocalMux I__2373 (
            .O(N__10481),
            .I(N__10425));
    LocalMux I__2372 (
            .O(N__10476),
            .I(N__10418));
    LocalMux I__2371 (
            .O(N__10471),
            .I(N__10418));
    Span4Mux_h I__2370 (
            .O(N__10462),
            .I(N__10418));
    InMux I__2369 (
            .O(N__10461),
            .I(N__10415));
    InMux I__2368 (
            .O(N__10460),
            .I(N__10412));
    LocalMux I__2367 (
            .O(N__10457),
            .I(N__10409));
    Span4Mux_h I__2366 (
            .O(N__10452),
            .I(N__10406));
    InMux I__2365 (
            .O(N__10451),
            .I(N__10401));
    InMux I__2364 (
            .O(N__10450),
            .I(N__10401));
    Span4Mux_h I__2363 (
            .O(N__10443),
            .I(N__10398));
    InMux I__2362 (
            .O(N__10442),
            .I(N__10393));
    InMux I__2361 (
            .O(N__10441),
            .I(N__10393));
    InMux I__2360 (
            .O(N__10440),
            .I(N__10388));
    InMux I__2359 (
            .O(N__10439),
            .I(N__10388));
    LocalMux I__2358 (
            .O(N__10436),
            .I(N__10385));
    LocalMux I__2357 (
            .O(N__10433),
            .I(N__10374));
    LocalMux I__2356 (
            .O(N__10430),
            .I(N__10374));
    Span4Mux_v I__2355 (
            .O(N__10425),
            .I(N__10374));
    Span4Mux_v I__2354 (
            .O(N__10418),
            .I(N__10374));
    LocalMux I__2353 (
            .O(N__10415),
            .I(N__10374));
    LocalMux I__2352 (
            .O(N__10412),
            .I(N__10371));
    Odrv4 I__2351 (
            .O(N__10409),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2350 (
            .O(N__10406),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2349 (
            .O(N__10401),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2348 (
            .O(N__10398),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2347 (
            .O(N__10393),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2346 (
            .O(N__10388),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2345 (
            .O(N__10385),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2344 (
            .O(N__10374),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2343 (
            .O(N__10371),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    InMux I__2342 (
            .O(N__10352),
            .I(N__10349));
    LocalMux I__2341 (
            .O(N__10349),
            .I(\U712_CHIP_RAM.m158_xx_mm_0_2 ));
    IoInMux I__2340 (
            .O(N__10346),
            .I(N__10343));
    LocalMux I__2339 (
            .O(N__10343),
            .I(N__10340));
    Span4Mux_s2_h I__2338 (
            .O(N__10340),
            .I(N__10337));
    Sp12to4 I__2337 (
            .O(N__10337),
            .I(N__10334));
    Span12Mux_s11_v I__2336 (
            .O(N__10334),
            .I(N__10331));
    Odrv12 I__2335 (
            .O(N__10331),
            .I(CMA_c_3));
    CEMux I__2334 (
            .O(N__10328),
            .I(N__10322));
    CEMux I__2333 (
            .O(N__10327),
            .I(N__10316));
    CEMux I__2332 (
            .O(N__10326),
            .I(N__10312));
    CEMux I__2331 (
            .O(N__10325),
            .I(N__10309));
    LocalMux I__2330 (
            .O(N__10322),
            .I(N__10306));
    CEMux I__2329 (
            .O(N__10321),
            .I(N__10303));
    CEMux I__2328 (
            .O(N__10320),
            .I(N__10300));
    CEMux I__2327 (
            .O(N__10319),
            .I(N__10297));
    LocalMux I__2326 (
            .O(N__10316),
            .I(N__10294));
    CEMux I__2325 (
            .O(N__10315),
            .I(N__10290));
    LocalMux I__2324 (
            .O(N__10312),
            .I(N__10287));
    LocalMux I__2323 (
            .O(N__10309),
            .I(N__10284));
    Span4Mux_v I__2322 (
            .O(N__10306),
            .I(N__10279));
    LocalMux I__2321 (
            .O(N__10303),
            .I(N__10279));
    LocalMux I__2320 (
            .O(N__10300),
            .I(N__10272));
    LocalMux I__2319 (
            .O(N__10297),
            .I(N__10272));
    Span4Mux_h I__2318 (
            .O(N__10294),
            .I(N__10272));
    CEMux I__2317 (
            .O(N__10293),
            .I(N__10269));
    LocalMux I__2316 (
            .O(N__10290),
            .I(N__10266));
    Span4Mux_v I__2315 (
            .O(N__10287),
            .I(N__10261));
    Span4Mux_h I__2314 (
            .O(N__10284),
            .I(N__10261));
    Span4Mux_h I__2313 (
            .O(N__10279),
            .I(N__10258));
    Span4Mux_h I__2312 (
            .O(N__10272),
            .I(N__10255));
    LocalMux I__2311 (
            .O(N__10269),
            .I(\U712_CHIP_RAM.N_168_0_0 ));
    Odrv12 I__2310 (
            .O(N__10266),
            .I(\U712_CHIP_RAM.N_168_0_0 ));
    Odrv4 I__2309 (
            .O(N__10261),
            .I(\U712_CHIP_RAM.N_168_0_0 ));
    Odrv4 I__2308 (
            .O(N__10258),
            .I(\U712_CHIP_RAM.N_168_0_0 ));
    Odrv4 I__2307 (
            .O(N__10255),
            .I(\U712_CHIP_RAM.N_168_0_0 ));
    InMux I__2306 (
            .O(N__10244),
            .I(N__10238));
    InMux I__2305 (
            .O(N__10243),
            .I(N__10235));
    CascadeMux I__2304 (
            .O(N__10242),
            .I(N__10229));
    InMux I__2303 (
            .O(N__10241),
            .I(N__10221));
    LocalMux I__2302 (
            .O(N__10238),
            .I(N__10218));
    LocalMux I__2301 (
            .O(N__10235),
            .I(N__10215));
    InMux I__2300 (
            .O(N__10234),
            .I(N__10212));
    InMux I__2299 (
            .O(N__10233),
            .I(N__10205));
    InMux I__2298 (
            .O(N__10232),
            .I(N__10205));
    InMux I__2297 (
            .O(N__10229),
            .I(N__10205));
    InMux I__2296 (
            .O(N__10228),
            .I(N__10198));
    InMux I__2295 (
            .O(N__10227),
            .I(N__10198));
    InMux I__2294 (
            .O(N__10226),
            .I(N__10198));
    InMux I__2293 (
            .O(N__10225),
            .I(N__10193));
    InMux I__2292 (
            .O(N__10224),
            .I(N__10193));
    LocalMux I__2291 (
            .O(N__10221),
            .I(N__10188));
    Span4Mux_h I__2290 (
            .O(N__10218),
            .I(N__10188));
    Odrv4 I__2289 (
            .O(N__10215),
            .I(\U712_CHIP_RAM.N_3_0 ));
    LocalMux I__2288 (
            .O(N__10212),
            .I(\U712_CHIP_RAM.N_3_0 ));
    LocalMux I__2287 (
            .O(N__10205),
            .I(\U712_CHIP_RAM.N_3_0 ));
    LocalMux I__2286 (
            .O(N__10198),
            .I(\U712_CHIP_RAM.N_3_0 ));
    LocalMux I__2285 (
            .O(N__10193),
            .I(\U712_CHIP_RAM.N_3_0 ));
    Odrv4 I__2284 (
            .O(N__10188),
            .I(\U712_CHIP_RAM.N_3_0 ));
    IoInMux I__2283 (
            .O(N__10175),
            .I(N__10172));
    LocalMux I__2282 (
            .O(N__10172),
            .I(N__10169));
    Span4Mux_s2_v I__2281 (
            .O(N__10169),
            .I(N__10166));
    Span4Mux_v I__2280 (
            .O(N__10166),
            .I(N__10163));
    Span4Mux_v I__2279 (
            .O(N__10163),
            .I(N__10160));
    Span4Mux_v I__2278 (
            .O(N__10160),
            .I(N__10157));
    Odrv4 I__2277 (
            .O(N__10157),
            .I(CMA_c_10));
    InMux I__2276 (
            .O(N__10154),
            .I(N__10150));
    InMux I__2275 (
            .O(N__10153),
            .I(N__10147));
    LocalMux I__2274 (
            .O(N__10150),
            .I(N__10140));
    LocalMux I__2273 (
            .O(N__10147),
            .I(N__10140));
    InMux I__2272 (
            .O(N__10146),
            .I(N__10137));
    InMux I__2271 (
            .O(N__10145),
            .I(N__10134));
    Span4Mux_v I__2270 (
            .O(N__10140),
            .I(N__10131));
    LocalMux I__2269 (
            .O(N__10137),
            .I(N__10128));
    LocalMux I__2268 (
            .O(N__10134),
            .I(N__10125));
    Sp12to4 I__2267 (
            .O(N__10131),
            .I(N__10122));
    Span4Mux_v I__2266 (
            .O(N__10128),
            .I(N__10117));
    Span4Mux_v I__2265 (
            .O(N__10125),
            .I(N__10117));
    Span12Mux_h I__2264 (
            .O(N__10122),
            .I(N__10114));
    Sp12to4 I__2263 (
            .O(N__10117),
            .I(N__10111));
    Odrv12 I__2262 (
            .O(N__10114),
            .I(DRA_c_8));
    Odrv12 I__2261 (
            .O(N__10111),
            .I(DRA_c_8));
    InMux I__2260 (
            .O(N__10106),
            .I(N__10103));
    LocalMux I__2259 (
            .O(N__10103),
            .I(N__10100));
    Odrv12 I__2258 (
            .O(N__10100),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2257 (
            .O(N__10097),
            .I(N__10094));
    LocalMux I__2256 (
            .O(N__10094),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ));
    InMux I__2255 (
            .O(N__10091),
            .I(N__10088));
    LocalMux I__2254 (
            .O(N__10088),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_5 ));
    InMux I__2253 (
            .O(N__10085),
            .I(N__10082));
    LocalMux I__2252 (
            .O(N__10082),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ));
    InMux I__2251 (
            .O(N__10079),
            .I(N__10075));
    InMux I__2250 (
            .O(N__10078),
            .I(N__10072));
    LocalMux I__2249 (
            .O(N__10075),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ));
    LocalMux I__2248 (
            .O(N__10072),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ));
    InMux I__2247 (
            .O(N__10067),
            .I(N__10064));
    LocalMux I__2246 (
            .O(N__10064),
            .I(N__10061));
    Span4Mux_v I__2245 (
            .O(N__10061),
            .I(N__10058));
    Span4Mux_h I__2244 (
            .O(N__10058),
            .I(N__10055));
    Odrv4 I__2243 (
            .O(N__10055),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    InMux I__2242 (
            .O(N__10052),
            .I(N__10049));
    LocalMux I__2241 (
            .O(N__10049),
            .I(\U712_CHIP_RAM.m158_xx_mm_0_0 ));
    CascadeMux I__2240 (
            .O(N__10046),
            .I(N__10042));
    CascadeMux I__2239 (
            .O(N__10045),
            .I(N__10039));
    InMux I__2238 (
            .O(N__10042),
            .I(N__10035));
    InMux I__2237 (
            .O(N__10039),
            .I(N__10029));
    InMux I__2236 (
            .O(N__10038),
            .I(N__10025));
    LocalMux I__2235 (
            .O(N__10035),
            .I(N__10022));
    InMux I__2234 (
            .O(N__10034),
            .I(N__10017));
    InMux I__2233 (
            .O(N__10033),
            .I(N__10012));
    InMux I__2232 (
            .O(N__10032),
            .I(N__10012));
    LocalMux I__2231 (
            .O(N__10029),
            .I(N__10009));
    InMux I__2230 (
            .O(N__10028),
            .I(N__10006));
    LocalMux I__2229 (
            .O(N__10025),
            .I(N__10003));
    Span4Mux_h I__2228 (
            .O(N__10022),
            .I(N__10000));
    InMux I__2227 (
            .O(N__10021),
            .I(N__9997));
    InMux I__2226 (
            .O(N__10020),
            .I(N__9994));
    LocalMux I__2225 (
            .O(N__10017),
            .I(N__9987));
    LocalMux I__2224 (
            .O(N__10012),
            .I(N__9987));
    Span4Mux_h I__2223 (
            .O(N__10009),
            .I(N__9987));
    LocalMux I__2222 (
            .O(N__10006),
            .I(N__9980));
    Span4Mux_v I__2221 (
            .O(N__10003),
            .I(N__9980));
    Span4Mux_v I__2220 (
            .O(N__10000),
            .I(N__9980));
    LocalMux I__2219 (
            .O(N__9997),
            .I(\U712_CHIP_RAM.m154_a2_0 ));
    LocalMux I__2218 (
            .O(N__9994),
            .I(\U712_CHIP_RAM.m154_a2_0 ));
    Odrv4 I__2217 (
            .O(N__9987),
            .I(\U712_CHIP_RAM.m154_a2_0 ));
    Odrv4 I__2216 (
            .O(N__9980),
            .I(\U712_CHIP_RAM.m154_a2_0 ));
    InMux I__2215 (
            .O(N__9971),
            .I(N__9965));
    InMux I__2214 (
            .O(N__9970),
            .I(N__9962));
    InMux I__2213 (
            .O(N__9969),
            .I(N__9959));
    InMux I__2212 (
            .O(N__9968),
            .I(N__9956));
    LocalMux I__2211 (
            .O(N__9965),
            .I(N__9953));
    LocalMux I__2210 (
            .O(N__9962),
            .I(N__9946));
    LocalMux I__2209 (
            .O(N__9959),
            .I(N__9946));
    LocalMux I__2208 (
            .O(N__9956),
            .I(N__9946));
    Span4Mux_v I__2207 (
            .O(N__9953),
            .I(N__9943));
    Span4Mux_v I__2206 (
            .O(N__9946),
            .I(N__9940));
    Span4Mux_h I__2205 (
            .O(N__9943),
            .I(N__9937));
    Span4Mux_h I__2204 (
            .O(N__9940),
            .I(N__9934));
    Sp12to4 I__2203 (
            .O(N__9937),
            .I(N__9929));
    Sp12to4 I__2202 (
            .O(N__9934),
            .I(N__9929));
    Odrv12 I__2201 (
            .O(N__9929),
            .I(DRA_c_7));
    InMux I__2200 (
            .O(N__9926),
            .I(N__9923));
    LocalMux I__2199 (
            .O(N__9923),
            .I(N__9919));
    InMux I__2198 (
            .O(N__9922),
            .I(N__9916));
    Span4Mux_v I__2197 (
            .O(N__9919),
            .I(N__9909));
    LocalMux I__2196 (
            .O(N__9916),
            .I(N__9909));
    InMux I__2195 (
            .O(N__9915),
            .I(N__9906));
    InMux I__2194 (
            .O(N__9914),
            .I(N__9903));
    Span4Mux_h I__2193 (
            .O(N__9909),
            .I(N__9898));
    LocalMux I__2192 (
            .O(N__9906),
            .I(N__9898));
    LocalMux I__2191 (
            .O(N__9903),
            .I(N__9895));
    Span4Mux_v I__2190 (
            .O(N__9898),
            .I(N__9892));
    Sp12to4 I__2189 (
            .O(N__9895),
            .I(N__9889));
    Sp12to4 I__2188 (
            .O(N__9892),
            .I(N__9886));
    Span12Mux_v I__2187 (
            .O(N__9889),
            .I(N__9883));
    Span12Mux_h I__2186 (
            .O(N__9886),
            .I(N__9880));
    Odrv12 I__2185 (
            .O(N__9883),
            .I(DRA_c_6));
    Odrv12 I__2184 (
            .O(N__9880),
            .I(DRA_c_6));
    InMux I__2183 (
            .O(N__9875),
            .I(N__9872));
    LocalMux I__2182 (
            .O(N__9872),
            .I(N__9869));
    Span4Mux_h I__2181 (
            .O(N__9869),
            .I(N__9866));
    Odrv4 I__2180 (
            .O(N__9866),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2179 (
            .O(N__9863),
            .I(N__9860));
    LocalMux I__2178 (
            .O(N__9860),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2177 (
            .O(N__9857),
            .I(N__9854));
    LocalMux I__2176 (
            .O(N__9854),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2175 (
            .O(N__9851),
            .I(N__9848));
    LocalMux I__2174 (
            .O(N__9848),
            .I(N__9845));
    Span4Mux_h I__2173 (
            .O(N__9845),
            .I(N__9842));
    Odrv4 I__2172 (
            .O(N__9842),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2171 (
            .O(N__9839),
            .I(N__9836));
    LocalMux I__2170 (
            .O(N__9836),
            .I(N__9833));
    Span4Mux_h I__2169 (
            .O(N__9833),
            .I(N__9830));
    Span4Mux_h I__2168 (
            .O(N__9830),
            .I(N__9827));
    Odrv4 I__2167 (
            .O(N__9827),
            .I(\U712_CHIP_RAM.m228_0 ));
    InMux I__2166 (
            .O(N__9824),
            .I(N__9818));
    InMux I__2165 (
            .O(N__9823),
            .I(N__9818));
    LocalMux I__2164 (
            .O(N__9818),
            .I(\U712_CHIP_RAM.N_343 ));
    InMux I__2163 (
            .O(N__9815),
            .I(N__9810));
    InMux I__2162 (
            .O(N__9814),
            .I(N__9806));
    InMux I__2161 (
            .O(N__9813),
            .I(N__9803));
    LocalMux I__2160 (
            .O(N__9810),
            .I(N__9800));
    InMux I__2159 (
            .O(N__9809),
            .I(N__9797));
    LocalMux I__2158 (
            .O(N__9806),
            .I(N__9794));
    LocalMux I__2157 (
            .O(N__9803),
            .I(N__9791));
    Span4Mux_h I__2156 (
            .O(N__9800),
            .I(N__9787));
    LocalMux I__2155 (
            .O(N__9797),
            .I(N__9784));
    Span12Mux_h I__2154 (
            .O(N__9794),
            .I(N__9778));
    Span4Mux_h I__2153 (
            .O(N__9791),
            .I(N__9775));
    InMux I__2152 (
            .O(N__9790),
            .I(N__9772));
    Span4Mux_h I__2151 (
            .O(N__9787),
            .I(N__9767));
    Span4Mux_v I__2150 (
            .O(N__9784),
            .I(N__9767));
    InMux I__2149 (
            .O(N__9783),
            .I(N__9762));
    InMux I__2148 (
            .O(N__9782),
            .I(N__9762));
    InMux I__2147 (
            .O(N__9781),
            .I(N__9759));
    Odrv12 I__2146 (
            .O(N__9778),
            .I(\U712_CHIP_RAM.DMA_CYCLEm ));
    Odrv4 I__2145 (
            .O(N__9775),
            .I(\U712_CHIP_RAM.DMA_CYCLEm ));
    LocalMux I__2144 (
            .O(N__9772),
            .I(\U712_CHIP_RAM.DMA_CYCLEm ));
    Odrv4 I__2143 (
            .O(N__9767),
            .I(\U712_CHIP_RAM.DMA_CYCLEm ));
    LocalMux I__2142 (
            .O(N__9762),
            .I(\U712_CHIP_RAM.DMA_CYCLEm ));
    LocalMux I__2141 (
            .O(N__9759),
            .I(\U712_CHIP_RAM.DMA_CYCLEm ));
    InMux I__2140 (
            .O(N__9746),
            .I(N__9743));
    LocalMux I__2139 (
            .O(N__9743),
            .I(N__9739));
    InMux I__2138 (
            .O(N__9742),
            .I(N__9736));
    Span4Mux_v I__2137 (
            .O(N__9739),
            .I(N__9733));
    LocalMux I__2136 (
            .O(N__9736),
            .I(N__9730));
    Odrv4 I__2135 (
            .O(N__9733),
            .I(\U712_CHIP_RAM.N_342 ));
    Odrv4 I__2134 (
            .O(N__9730),
            .I(\U712_CHIP_RAM.N_342 ));
    InMux I__2133 (
            .O(N__9725),
            .I(N__9722));
    LocalMux I__2132 (
            .O(N__9722),
            .I(N__9719));
    Span4Mux_v I__2131 (
            .O(N__9719),
            .I(N__9716));
    Sp12to4 I__2130 (
            .O(N__9716),
            .I(N__9713));
    Span12Mux_h I__2129 (
            .O(N__9713),
            .I(N__9710));
    Odrv12 I__2128 (
            .O(N__9710),
            .I(A_c_12));
    CascadeMux I__2127 (
            .O(N__9707),
            .I(N__9704));
    InMux I__2126 (
            .O(N__9704),
            .I(N__9701));
    LocalMux I__2125 (
            .O(N__9701),
            .I(N__9698));
    Odrv12 I__2124 (
            .O(N__9698),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__2123 (
            .O(N__9695),
            .I(N__9692));
    LocalMux I__2122 (
            .O(N__9692),
            .I(N__9689));
    Odrv4 I__2121 (
            .O(N__9689),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__2120 (
            .O(N__9686),
            .I(N__9680));
    InMux I__2119 (
            .O(N__9685),
            .I(N__9680));
    LocalMux I__2118 (
            .O(N__9680),
            .I(N__9663));
    InMux I__2117 (
            .O(N__9679),
            .I(N__9660));
    InMux I__2116 (
            .O(N__9678),
            .I(N__9655));
    InMux I__2115 (
            .O(N__9677),
            .I(N__9655));
    InMux I__2114 (
            .O(N__9676),
            .I(N__9652));
    InMux I__2113 (
            .O(N__9675),
            .I(N__9647));
    InMux I__2112 (
            .O(N__9674),
            .I(N__9647));
    InMux I__2111 (
            .O(N__9673),
            .I(N__9642));
    InMux I__2110 (
            .O(N__9672),
            .I(N__9642));
    InMux I__2109 (
            .O(N__9671),
            .I(N__9635));
    InMux I__2108 (
            .O(N__9670),
            .I(N__9635));
    InMux I__2107 (
            .O(N__9669),
            .I(N__9635));
    InMux I__2106 (
            .O(N__9668),
            .I(N__9629));
    InMux I__2105 (
            .O(N__9667),
            .I(N__9626));
    InMux I__2104 (
            .O(N__9666),
            .I(N__9623));
    Span4Mux_v I__2103 (
            .O(N__9663),
            .I(N__9616));
    LocalMux I__2102 (
            .O(N__9660),
            .I(N__9613));
    LocalMux I__2101 (
            .O(N__9655),
            .I(N__9602));
    LocalMux I__2100 (
            .O(N__9652),
            .I(N__9602));
    LocalMux I__2099 (
            .O(N__9647),
            .I(N__9602));
    LocalMux I__2098 (
            .O(N__9642),
            .I(N__9602));
    LocalMux I__2097 (
            .O(N__9635),
            .I(N__9602));
    InMux I__2096 (
            .O(N__9634),
            .I(N__9595));
    InMux I__2095 (
            .O(N__9633),
            .I(N__9595));
    InMux I__2094 (
            .O(N__9632),
            .I(N__9595));
    LocalMux I__2093 (
            .O(N__9629),
            .I(N__9590));
    LocalMux I__2092 (
            .O(N__9626),
            .I(N__9590));
    LocalMux I__2091 (
            .O(N__9623),
            .I(N__9587));
    InMux I__2090 (
            .O(N__9622),
            .I(N__9580));
    InMux I__2089 (
            .O(N__9621),
            .I(N__9580));
    InMux I__2088 (
            .O(N__9620),
            .I(N__9580));
    InMux I__2087 (
            .O(N__9619),
            .I(N__9577));
    Span4Mux_h I__2086 (
            .O(N__9616),
            .I(N__9570));
    Span4Mux_v I__2085 (
            .O(N__9613),
            .I(N__9570));
    Span4Mux_v I__2084 (
            .O(N__9602),
            .I(N__9570));
    LocalMux I__2083 (
            .O(N__9595),
            .I(N__9567));
    Span4Mux_v I__2082 (
            .O(N__9590),
            .I(N__9560));
    Span4Mux_v I__2081 (
            .O(N__9587),
            .I(N__9553));
    LocalMux I__2080 (
            .O(N__9580),
            .I(N__9553));
    LocalMux I__2079 (
            .O(N__9577),
            .I(N__9553));
    Span4Mux_h I__2078 (
            .O(N__9570),
            .I(N__9548));
    Span4Mux_v I__2077 (
            .O(N__9567),
            .I(N__9548));
    InMux I__2076 (
            .O(N__9566),
            .I(N__9545));
    InMux I__2075 (
            .O(N__9565),
            .I(N__9540));
    InMux I__2074 (
            .O(N__9564),
            .I(N__9540));
    InMux I__2073 (
            .O(N__9563),
            .I(N__9537));
    Span4Mux_h I__2072 (
            .O(N__9560),
            .I(N__9532));
    Span4Mux_v I__2071 (
            .O(N__9553),
            .I(N__9532));
    Span4Mux_h I__2070 (
            .O(N__9548),
            .I(N__9529));
    LocalMux I__2069 (
            .O(N__9545),
            .I(N__9520));
    LocalMux I__2068 (
            .O(N__9540),
            .I(N__9520));
    LocalMux I__2067 (
            .O(N__9537),
            .I(N__9520));
    Sp12to4 I__2066 (
            .O(N__9532),
            .I(N__9520));
    Sp12to4 I__2065 (
            .O(N__9529),
            .I(N__9515));
    Span12Mux_h I__2064 (
            .O(N__9520),
            .I(N__9515));
    Odrv12 I__2063 (
            .O(N__9515),
            .I(RESETn_c));
    InMux I__2062 (
            .O(N__9512),
            .I(N__9505));
    InMux I__2061 (
            .O(N__9511),
            .I(N__9496));
    InMux I__2060 (
            .O(N__9510),
            .I(N__9496));
    InMux I__2059 (
            .O(N__9509),
            .I(N__9496));
    InMux I__2058 (
            .O(N__9508),
            .I(N__9496));
    LocalMux I__2057 (
            .O(N__9505),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__2056 (
            .O(N__9496),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__2055 (
            .O(N__9491),
            .I(N__9487));
    InMux I__2054 (
            .O(N__9490),
            .I(N__9483));
    InMux I__2053 (
            .O(N__9487),
            .I(N__9478));
    InMux I__2052 (
            .O(N__9486),
            .I(N__9478));
    LocalMux I__2051 (
            .O(N__9483),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__2050 (
            .O(N__9478),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__2049 (
            .O(N__9473),
            .I(N__9468));
    InMux I__2048 (
            .O(N__9472),
            .I(N__9463));
    InMux I__2047 (
            .O(N__9471),
            .I(N__9463));
    LocalMux I__2046 (
            .O(N__9468),
            .I(N__9457));
    LocalMux I__2045 (
            .O(N__9463),
            .I(N__9457));
    InMux I__2044 (
            .O(N__9462),
            .I(N__9454));
    Span4Mux_v I__2043 (
            .O(N__9457),
            .I(N__9451));
    LocalMux I__2042 (
            .O(N__9454),
            .I(\U712_CYCLE_TERM.TACK_STARTZ0 ));
    Odrv4 I__2041 (
            .O(N__9451),
            .I(\U712_CYCLE_TERM.TACK_STARTZ0 ));
    IoInMux I__2040 (
            .O(N__9446),
            .I(N__9442));
    IoInMux I__2039 (
            .O(N__9445),
            .I(N__9438));
    LocalMux I__2038 (
            .O(N__9442),
            .I(N__9435));
    IoInMux I__2037 (
            .O(N__9441),
            .I(N__9432));
    LocalMux I__2036 (
            .O(N__9438),
            .I(N__9429));
    IoSpan4Mux I__2035 (
            .O(N__9435),
            .I(N__9426));
    LocalMux I__2034 (
            .O(N__9432),
            .I(N__9423));
    Span4Mux_s3_v I__2033 (
            .O(N__9429),
            .I(N__9420));
    IoSpan4Mux I__2032 (
            .O(N__9426),
            .I(N__9417));
    Span12Mux_s3_v I__2031 (
            .O(N__9423),
            .I(N__9413));
    Sp12to4 I__2030 (
            .O(N__9420),
            .I(N__9410));
    Span4Mux_s2_h I__2029 (
            .O(N__9417),
            .I(N__9407));
    InMux I__2028 (
            .O(N__9416),
            .I(N__9403));
    Span12Mux_h I__2027 (
            .O(N__9413),
            .I(N__9398));
    Span12Mux_h I__2026 (
            .O(N__9410),
            .I(N__9398));
    Sp12to4 I__2025 (
            .O(N__9407),
            .I(N__9395));
    CascadeMux I__2024 (
            .O(N__9406),
            .I(N__9392));
    LocalMux I__2023 (
            .O(N__9403),
            .I(N__9389));
    Span12Mux_v I__2022 (
            .O(N__9398),
            .I(N__9386));
    Span12Mux_h I__2021 (
            .O(N__9395),
            .I(N__9383));
    InMux I__2020 (
            .O(N__9392),
            .I(N__9380));
    Span4Mux_h I__2019 (
            .O(N__9389),
            .I(N__9377));
    Odrv12 I__2018 (
            .O(N__9386),
            .I(TACK_EN));
    Odrv12 I__2017 (
            .O(N__9383),
            .I(TACK_EN));
    LocalMux I__2016 (
            .O(N__9380),
            .I(TACK_EN));
    Odrv4 I__2015 (
            .O(N__9377),
            .I(TACK_EN));
    InMux I__2014 (
            .O(N__9368),
            .I(N__9365));
    LocalMux I__2013 (
            .O(N__9365),
            .I(N__9357));
    InMux I__2012 (
            .O(N__9364),
            .I(N__9352));
    InMux I__2011 (
            .O(N__9363),
            .I(N__9342));
    InMux I__2010 (
            .O(N__9362),
            .I(N__9342));
    InMux I__2009 (
            .O(N__9361),
            .I(N__9342));
    InMux I__2008 (
            .O(N__9360),
            .I(N__9335));
    Span4Mux_v I__2007 (
            .O(N__9357),
            .I(N__9332));
    InMux I__2006 (
            .O(N__9356),
            .I(N__9329));
    InMux I__2005 (
            .O(N__9355),
            .I(N__9326));
    LocalMux I__2004 (
            .O(N__9352),
            .I(N__9323));
    InMux I__2003 (
            .O(N__9351),
            .I(N__9316));
    InMux I__2002 (
            .O(N__9350),
            .I(N__9316));
    InMux I__2001 (
            .O(N__9349),
            .I(N__9316));
    LocalMux I__2000 (
            .O(N__9342),
            .I(N__9313));
    InMux I__1999 (
            .O(N__9341),
            .I(N__9304));
    InMux I__1998 (
            .O(N__9340),
            .I(N__9304));
    InMux I__1997 (
            .O(N__9339),
            .I(N__9304));
    InMux I__1996 (
            .O(N__9338),
            .I(N__9304));
    LocalMux I__1995 (
            .O(N__9335),
            .I(U712_REG_SM_C1_SYNC_1));
    Odrv4 I__1994 (
            .O(N__9332),
            .I(U712_REG_SM_C1_SYNC_1));
    LocalMux I__1993 (
            .O(N__9329),
            .I(U712_REG_SM_C1_SYNC_1));
    LocalMux I__1992 (
            .O(N__9326),
            .I(U712_REG_SM_C1_SYNC_1));
    Odrv4 I__1991 (
            .O(N__9323),
            .I(U712_REG_SM_C1_SYNC_1));
    LocalMux I__1990 (
            .O(N__9316),
            .I(U712_REG_SM_C1_SYNC_1));
    Odrv4 I__1989 (
            .O(N__9313),
            .I(U712_REG_SM_C1_SYNC_1));
    LocalMux I__1988 (
            .O(N__9304),
            .I(U712_REG_SM_C1_SYNC_1));
    IoInMux I__1987 (
            .O(N__9287),
            .I(N__9284));
    LocalMux I__1986 (
            .O(N__9284),
            .I(N__9281));
    Span4Mux_s2_v I__1985 (
            .O(N__9281),
            .I(N__9278));
    Span4Mux_v I__1984 (
            .O(N__9278),
            .I(N__9275));
    Span4Mux_v I__1983 (
            .O(N__9275),
            .I(N__9272));
    Sp12to4 I__1982 (
            .O(N__9272),
            .I(N__9269));
    Odrv12 I__1981 (
            .O(N__9269),
            .I(ASn_c));
    CEMux I__1980 (
            .O(N__9266),
            .I(N__9263));
    LocalMux I__1979 (
            .O(N__9263),
            .I(\U712_REG_SM.N_33_0_0 ));
    IoInMux I__1978 (
            .O(N__9260),
            .I(N__9257));
    LocalMux I__1977 (
            .O(N__9257),
            .I(N__9254));
    IoSpan4Mux I__1976 (
            .O(N__9254),
            .I(N__9251));
    Span4Mux_s3_v I__1975 (
            .O(N__9251),
            .I(N__9248));
    Span4Mux_v I__1974 (
            .O(N__9248),
            .I(N__9245));
    Span4Mux_h I__1973 (
            .O(N__9245),
            .I(N__9242));
    Odrv4 I__1972 (
            .O(N__9242),
            .I(DMA_LATCH_EN_c));
    InMux I__1971 (
            .O(N__9239),
            .I(N__9236));
    LocalMux I__1970 (
            .O(N__9236),
            .I(\U712_CHIP_RAM.m160_xx_mm_0_2 ));
    IoInMux I__1969 (
            .O(N__9233),
            .I(N__9230));
    LocalMux I__1968 (
            .O(N__9230),
            .I(N__9227));
    Span12Mux_s1_h I__1967 (
            .O(N__9227),
            .I(N__9224));
    Span12Mux_h I__1966 (
            .O(N__9224),
            .I(N__9221));
    Odrv12 I__1965 (
            .O(N__9221),
            .I(CMA_c_6));
    InMux I__1964 (
            .O(N__9218),
            .I(N__9215));
    LocalMux I__1963 (
            .O(N__9215),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__1962 (
            .O(N__9212),
            .I(N__9209));
    LocalMux I__1961 (
            .O(N__9209),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1960 (
            .O(N__9206),
            .I(N__9203));
    LocalMux I__1959 (
            .O(N__9203),
            .I(N__9200));
    Span12Mux_v I__1958 (
            .O(N__9200),
            .I(N__9197));
    Span12Mux_h I__1957 (
            .O(N__9197),
            .I(N__9194));
    Odrv12 I__1956 (
            .O(N__9194),
            .I(A_c_14));
    InMux I__1955 (
            .O(N__9191),
            .I(N__9188));
    LocalMux I__1954 (
            .O(N__9188),
            .I(\U712_CHIP_RAM.m155_0_0 ));
    CascadeMux I__1953 (
            .O(N__9185),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_ ));
    InMux I__1952 (
            .O(N__9182),
            .I(N__9179));
    LocalMux I__1951 (
            .O(N__9179),
            .I(\U712_CHIP_RAM.m155_0_2 ));
    IoInMux I__1950 (
            .O(N__9176),
            .I(N__9173));
    LocalMux I__1949 (
            .O(N__9173),
            .I(N__9169));
    CascadeMux I__1948 (
            .O(N__9172),
            .I(N__9166));
    Span4Mux_s2_v I__1947 (
            .O(N__9169),
            .I(N__9163));
    InMux I__1946 (
            .O(N__9166),
            .I(N__9160));
    Span4Mux_h I__1945 (
            .O(N__9163),
            .I(N__9157));
    LocalMux I__1944 (
            .O(N__9160),
            .I(N__9154));
    Span4Mux_v I__1943 (
            .O(N__9157),
            .I(N__9151));
    Span12Mux_h I__1942 (
            .O(N__9154),
            .I(N__9148));
    Odrv4 I__1941 (
            .O(N__9151),
            .I(N_68_0));
    Odrv12 I__1940 (
            .O(N__9148),
            .I(N_68_0));
    IoInMux I__1939 (
            .O(N__9143),
            .I(N__9140));
    LocalMux I__1938 (
            .O(N__9140),
            .I(N__9137));
    Span4Mux_s2_h I__1937 (
            .O(N__9137),
            .I(N__9134));
    Sp12to4 I__1936 (
            .O(N__9134),
            .I(N__9131));
    Span12Mux_v I__1935 (
            .O(N__9131),
            .I(N__9128));
    Span12Mux_h I__1934 (
            .O(N__9128),
            .I(N__9125));
    Odrv12 I__1933 (
            .O(N__9125),
            .I(CUUBEn_c));
    InMux I__1932 (
            .O(N__9122),
            .I(N__9118));
    IoInMux I__1931 (
            .O(N__9121),
            .I(N__9115));
    LocalMux I__1930 (
            .O(N__9118),
            .I(N__9112));
    LocalMux I__1929 (
            .O(N__9115),
            .I(N__9109));
    Span4Mux_v I__1928 (
            .O(N__9112),
            .I(N__9106));
    Span12Mux_s10_v I__1927 (
            .O(N__9109),
            .I(N__9103));
    Span4Mux_v I__1926 (
            .O(N__9106),
            .I(N__9100));
    Odrv12 I__1925 (
            .O(N__9103),
            .I(N_145_0));
    Odrv4 I__1924 (
            .O(N__9100),
            .I(N_145_0));
    IoInMux I__1923 (
            .O(N__9095),
            .I(N__9092));
    LocalMux I__1922 (
            .O(N__9092),
            .I(N__9089));
    IoSpan4Mux I__1921 (
            .O(N__9089),
            .I(N__9086));
    Span4Mux_s2_v I__1920 (
            .O(N__9086),
            .I(N__9083));
    Sp12to4 I__1919 (
            .O(N__9083),
            .I(N__9080));
    Span12Mux_v I__1918 (
            .O(N__9080),
            .I(N__9077));
    Odrv12 I__1917 (
            .O(N__9077),
            .I(CLLBEn_c));
    IoInMux I__1916 (
            .O(N__9074),
            .I(N__9069));
    InMux I__1915 (
            .O(N__9073),
            .I(N__9066));
    InMux I__1914 (
            .O(N__9072),
            .I(N__9063));
    LocalMux I__1913 (
            .O(N__9069),
            .I(N__9060));
    LocalMux I__1912 (
            .O(N__9066),
            .I(N__9057));
    LocalMux I__1911 (
            .O(N__9063),
            .I(N__9054));
    Span12Mux_s4_v I__1910 (
            .O(N__9060),
            .I(N__9049));
    Span4Mux_v I__1909 (
            .O(N__9057),
            .I(N__9046));
    Span4Mux_v I__1908 (
            .O(N__9054),
            .I(N__9043));
    InMux I__1907 (
            .O(N__9053),
            .I(N__9038));
    InMux I__1906 (
            .O(N__9052),
            .I(N__9038));
    Span12Mux_v I__1905 (
            .O(N__9049),
            .I(N__9028));
    Sp12to4 I__1904 (
            .O(N__9046),
            .I(N__9028));
    Sp12to4 I__1903 (
            .O(N__9043),
            .I(N__9028));
    LocalMux I__1902 (
            .O(N__9038),
            .I(N__9028));
    InMux I__1901 (
            .O(N__9037),
            .I(N__9025));
    Odrv12 I__1900 (
            .O(N__9028),
            .I(DBENn_c));
    LocalMux I__1899 (
            .O(N__9025),
            .I(DBENn_c));
    CascadeMux I__1898 (
            .O(N__9020),
            .I(N__9017));
    InMux I__1897 (
            .O(N__9017),
            .I(N__9013));
    IoInMux I__1896 (
            .O(N__9016),
            .I(N__9010));
    LocalMux I__1895 (
            .O(N__9013),
            .I(N__9007));
    LocalMux I__1894 (
            .O(N__9010),
            .I(N__9004));
    Span4Mux_v I__1893 (
            .O(N__9007),
            .I(N__9001));
    Span12Mux_s10_v I__1892 (
            .O(N__9004),
            .I(N__8998));
    Span4Mux_v I__1891 (
            .O(N__9001),
            .I(N__8995));
    Odrv12 I__1890 (
            .O(N__8998),
            .I(N_71_0));
    Odrv4 I__1889 (
            .O(N__8995),
            .I(N_71_0));
    IoInMux I__1888 (
            .O(N__8990),
            .I(N__8987));
    LocalMux I__1887 (
            .O(N__8987),
            .I(N__8984));
    Span4Mux_s2_h I__1886 (
            .O(N__8984),
            .I(N__8981));
    Sp12to4 I__1885 (
            .O(N__8981),
            .I(N__8978));
    Span12Mux_v I__1884 (
            .O(N__8978),
            .I(N__8975));
    Span12Mux_h I__1883 (
            .O(N__8975),
            .I(N__8972));
    Odrv12 I__1882 (
            .O(N__8972),
            .I(CUMBEn_c));
    InMux I__1881 (
            .O(N__8969),
            .I(N__8966));
    LocalMux I__1880 (
            .O(N__8966),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__1879 (
            .O(N__8963),
            .I(N__8959));
    InMux I__1878 (
            .O(N__8962),
            .I(N__8953));
    LocalMux I__1877 (
            .O(N__8959),
            .I(N__8950));
    CascadeMux I__1876 (
            .O(N__8958),
            .I(N__8946));
    CascadeMux I__1875 (
            .O(N__8957),
            .I(N__8943));
    CascadeMux I__1874 (
            .O(N__8956),
            .I(N__8940));
    LocalMux I__1873 (
            .O(N__8953),
            .I(N__8935));
    Span4Mux_v I__1872 (
            .O(N__8950),
            .I(N__8935));
    InMux I__1871 (
            .O(N__8949),
            .I(N__8928));
    InMux I__1870 (
            .O(N__8946),
            .I(N__8928));
    InMux I__1869 (
            .O(N__8943),
            .I(N__8928));
    InMux I__1868 (
            .O(N__8940),
            .I(N__8925));
    Span4Mux_h I__1867 (
            .O(N__8935),
            .I(N__8922));
    LocalMux I__1866 (
            .O(N__8928),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__1865 (
            .O(N__8925),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    Odrv4 I__1864 (
            .O(N__8922),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    CascadeMux I__1863 (
            .O(N__8915),
            .I(\U712_CYCLE_TERM.N_36_0_cascade_ ));
    IoInMux I__1862 (
            .O(N__8912),
            .I(N__8908));
    IoInMux I__1861 (
            .O(N__8911),
            .I(N__8905));
    LocalMux I__1860 (
            .O(N__8908),
            .I(N__8902));
    LocalMux I__1859 (
            .O(N__8905),
            .I(N__8899));
    Span4Mux_s2_v I__1858 (
            .O(N__8902),
            .I(N__8895));
    Span4Mux_s1_h I__1857 (
            .O(N__8899),
            .I(N__8892));
    IoInMux I__1856 (
            .O(N__8898),
            .I(N__8889));
    Span4Mux_v I__1855 (
            .O(N__8895),
            .I(N__8886));
    Span4Mux_h I__1854 (
            .O(N__8892),
            .I(N__8883));
    LocalMux I__1853 (
            .O(N__8889),
            .I(N__8880));
    Sp12to4 I__1852 (
            .O(N__8886),
            .I(N__8877));
    Sp12to4 I__1851 (
            .O(N__8883),
            .I(N__8874));
    Span12Mux_s10_v I__1850 (
            .O(N__8880),
            .I(N__8871));
    Span12Mux_h I__1849 (
            .O(N__8877),
            .I(N__8868));
    Span12Mux_v I__1848 (
            .O(N__8874),
            .I(N__8865));
    Span12Mux_h I__1847 (
            .O(N__8871),
            .I(N__8861));
    Span12Mux_v I__1846 (
            .O(N__8868),
            .I(N__8856));
    Span12Mux_h I__1845 (
            .O(N__8865),
            .I(N__8856));
    InMux I__1844 (
            .O(N__8864),
            .I(N__8853));
    Odrv12 I__1843 (
            .O(N__8861),
            .I(TACK_OUT));
    Odrv12 I__1842 (
            .O(N__8856),
            .I(TACK_OUT));
    LocalMux I__1841 (
            .O(N__8853),
            .I(TACK_OUT));
    InMux I__1840 (
            .O(N__8846),
            .I(N__8842));
    InMux I__1839 (
            .O(N__8845),
            .I(N__8834));
    LocalMux I__1838 (
            .O(N__8842),
            .I(N__8831));
    InMux I__1837 (
            .O(N__8841),
            .I(N__8828));
    CascadeMux I__1836 (
            .O(N__8840),
            .I(N__8825));
    InMux I__1835 (
            .O(N__8839),
            .I(N__8817));
    InMux I__1834 (
            .O(N__8838),
            .I(N__8817));
    InMux I__1833 (
            .O(N__8837),
            .I(N__8817));
    LocalMux I__1832 (
            .O(N__8834),
            .I(N__8814));
    Span4Mux_v I__1831 (
            .O(N__8831),
            .I(N__8809));
    LocalMux I__1830 (
            .O(N__8828),
            .I(N__8809));
    InMux I__1829 (
            .O(N__8825),
            .I(N__8806));
    InMux I__1828 (
            .O(N__8824),
            .I(N__8803));
    LocalMux I__1827 (
            .O(N__8817),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__1826 (
            .O(N__8814),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__1825 (
            .O(N__8809),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1824 (
            .O(N__8806),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1823 (
            .O(N__8803),
            .I(DBR_SYNCZ0Z_1));
    InMux I__1822 (
            .O(N__8792),
            .I(N__8788));
    CascadeMux I__1821 (
            .O(N__8791),
            .I(N__8785));
    LocalMux I__1820 (
            .O(N__8788),
            .I(N__8782));
    InMux I__1819 (
            .O(N__8785),
            .I(N__8779));
    Odrv4 I__1818 (
            .O(N__8782),
            .I(DBR_SYNC_i_1));
    LocalMux I__1817 (
            .O(N__8779),
            .I(DBR_SYNC_i_1));
    InMux I__1816 (
            .O(N__8774),
            .I(N__8770));
    InMux I__1815 (
            .O(N__8773),
            .I(N__8767));
    LocalMux I__1814 (
            .O(N__8770),
            .I(N__8761));
    LocalMux I__1813 (
            .O(N__8767),
            .I(N__8761));
    InMux I__1812 (
            .O(N__8766),
            .I(N__8758));
    Span4Mux_h I__1811 (
            .O(N__8761),
            .I(N__8755));
    LocalMux I__1810 (
            .O(N__8758),
            .I(N_33_0));
    Odrv4 I__1809 (
            .O(N__8755),
            .I(N_33_0));
    InMux I__1808 (
            .O(N__8750),
            .I(N__8745));
    CascadeMux I__1807 (
            .O(N__8749),
            .I(N__8741));
    InMux I__1806 (
            .O(N__8748),
            .I(N__8738));
    LocalMux I__1805 (
            .O(N__8745),
            .I(N__8735));
    CascadeMux I__1804 (
            .O(N__8744),
            .I(N__8732));
    InMux I__1803 (
            .O(N__8741),
            .I(N__8728));
    LocalMux I__1802 (
            .O(N__8738),
            .I(N__8725));
    Span4Mux_v I__1801 (
            .O(N__8735),
            .I(N__8722));
    InMux I__1800 (
            .O(N__8732),
            .I(N__8719));
    InMux I__1799 (
            .O(N__8731),
            .I(N__8716));
    LocalMux I__1798 (
            .O(N__8728),
            .I(N__8711));
    Span4Mux_v I__1797 (
            .O(N__8725),
            .I(N__8711));
    Span4Mux_h I__1796 (
            .O(N__8722),
            .I(N__8706));
    LocalMux I__1795 (
            .O(N__8719),
            .I(N__8706));
    LocalMux I__1794 (
            .O(N__8716),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1793 (
            .O(N__8711),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1792 (
            .O(N__8706),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__1791 (
            .O(N__8699),
            .I(N__8696));
    LocalMux I__1790 (
            .O(N__8696),
            .I(N__8693));
    IoSpan4Mux I__1789 (
            .O(N__8693),
            .I(N__8690));
    Sp12to4 I__1788 (
            .O(N__8690),
            .I(N__8687));
    Span12Mux_s9_v I__1787 (
            .O(N__8687),
            .I(N__8684));
    Odrv12 I__1786 (
            .O(N__8684),
            .I(RASn_c));
    InMux I__1785 (
            .O(N__8681),
            .I(N__8678));
    LocalMux I__1784 (
            .O(N__8678),
            .I(N__8675));
    Span4Mux_v I__1783 (
            .O(N__8675),
            .I(N__8672));
    Span4Mux_v I__1782 (
            .O(N__8672),
            .I(N__8669));
    Sp12to4 I__1781 (
            .O(N__8669),
            .I(N__8666));
    Span12Mux_h I__1780 (
            .O(N__8666),
            .I(N__8663));
    Odrv12 I__1779 (
            .O(N__8663),
            .I(A_c_19));
    IoInMux I__1778 (
            .O(N__8660),
            .I(N__8657));
    LocalMux I__1777 (
            .O(N__8657),
            .I(N__8654));
    IoSpan4Mux I__1776 (
            .O(N__8654),
            .I(N__8651));
    Span4Mux_s0_h I__1775 (
            .O(N__8651),
            .I(N__8648));
    Sp12to4 I__1774 (
            .O(N__8648),
            .I(N__8645));
    Span12Mux_h I__1773 (
            .O(N__8645),
            .I(N__8642));
    Odrv12 I__1772 (
            .O(N__8642),
            .I(CMA_c_9));
    InMux I__1771 (
            .O(N__8639),
            .I(N__8636));
    LocalMux I__1770 (
            .O(N__8636),
            .I(N__8633));
    Span4Mux_h I__1769 (
            .O(N__8633),
            .I(N__8630));
    Span4Mux_h I__1768 (
            .O(N__8630),
            .I(N__8627));
    Odrv4 I__1767 (
            .O(N__8627),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    InMux I__1766 (
            .O(N__8624),
            .I(N__8621));
    LocalMux I__1765 (
            .O(N__8621),
            .I(\U712_CHIP_RAM.m160_xx_mm_0_0 ));
    InMux I__1764 (
            .O(N__8618),
            .I(N__8613));
    InMux I__1763 (
            .O(N__8617),
            .I(N__8610));
    InMux I__1762 (
            .O(N__8616),
            .I(N__8607));
    LocalMux I__1761 (
            .O(N__8613),
            .I(\U712_CHIP_RAM.m164_0 ));
    LocalMux I__1760 (
            .O(N__8610),
            .I(\U712_CHIP_RAM.m164_0 ));
    LocalMux I__1759 (
            .O(N__8607),
            .I(\U712_CHIP_RAM.m164_0 ));
    IoInMux I__1758 (
            .O(N__8600),
            .I(N__8597));
    LocalMux I__1757 (
            .O(N__8597),
            .I(N__8594));
    Span4Mux_s2_h I__1756 (
            .O(N__8594),
            .I(N__8591));
    Sp12to4 I__1755 (
            .O(N__8591),
            .I(N__8588));
    Span12Mux_s10_v I__1754 (
            .O(N__8588),
            .I(N__8585));
    Span12Mux_h I__1753 (
            .O(N__8585),
            .I(N__8582));
    Odrv12 I__1752 (
            .O(N__8582),
            .I(CMA_c_5));
    CascadeMux I__1751 (
            .O(N__8579),
            .I(N__8576));
    InMux I__1750 (
            .O(N__8576),
            .I(N__8573));
    LocalMux I__1749 (
            .O(N__8573),
            .I(\U712_CHIP_RAM.m159_xx_mm_0_2 ));
    IoInMux I__1748 (
            .O(N__8570),
            .I(N__8567));
    LocalMux I__1747 (
            .O(N__8567),
            .I(N__8564));
    Span4Mux_s3_h I__1746 (
            .O(N__8564),
            .I(N__8561));
    Sp12to4 I__1745 (
            .O(N__8561),
            .I(N__8558));
    Span12Mux_v I__1744 (
            .O(N__8558),
            .I(N__8555));
    Odrv12 I__1743 (
            .O(N__8555),
            .I(CMA_c_4));
    CascadeMux I__1742 (
            .O(N__8552),
            .I(N__8549));
    InMux I__1741 (
            .O(N__8549),
            .I(N__8546));
    LocalMux I__1740 (
            .O(N__8546),
            .I(\U712_CHIP_RAM.m161_xx_mm_0_2 ));
    IoInMux I__1739 (
            .O(N__8543),
            .I(N__8540));
    LocalMux I__1738 (
            .O(N__8540),
            .I(N__8537));
    IoSpan4Mux I__1737 (
            .O(N__8537),
            .I(N__8534));
    Span4Mux_s3_h I__1736 (
            .O(N__8534),
            .I(N__8531));
    Sp12to4 I__1735 (
            .O(N__8531),
            .I(N__8528));
    Span12Mux_h I__1734 (
            .O(N__8528),
            .I(N__8525));
    Odrv12 I__1733 (
            .O(N__8525),
            .I(CMA_c_7));
    InMux I__1732 (
            .O(N__8522),
            .I(N__8518));
    InMux I__1731 (
            .O(N__8521),
            .I(N__8515));
    LocalMux I__1730 (
            .O(N__8518),
            .I(N__8510));
    LocalMux I__1729 (
            .O(N__8515),
            .I(N__8510));
    Odrv12 I__1728 (
            .O(N__8510),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ));
    InMux I__1727 (
            .O(N__8507),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ));
    InMux I__1726 (
            .O(N__8504),
            .I(N__8501));
    LocalMux I__1725 (
            .O(N__8501),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ));
    InMux I__1724 (
            .O(N__8498),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ));
    InMux I__1723 (
            .O(N__8495),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ));
    InMux I__1722 (
            .O(N__8492),
            .I(N__8486));
    InMux I__1721 (
            .O(N__8491),
            .I(N__8486));
    LocalMux I__1720 (
            .O(N__8486),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ));
    InMux I__1719 (
            .O(N__8483),
            .I(N__8480));
    LocalMux I__1718 (
            .O(N__8480),
            .I(N__8477));
    Odrv4 I__1717 (
            .O(N__8477),
            .I(\U712_CHIP_RAM.N_325 ));
    InMux I__1716 (
            .O(N__8474),
            .I(N__8471));
    LocalMux I__1715 (
            .O(N__8471),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ));
    CascadeMux I__1714 (
            .O(N__8468),
            .I(N__8465));
    InMux I__1713 (
            .O(N__8465),
            .I(N__8459));
    InMux I__1712 (
            .O(N__8464),
            .I(N__8459));
    LocalMux I__1711 (
            .O(N__8459),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_1 ));
    CascadeMux I__1710 (
            .O(N__8456),
            .I(N__8453));
    InMux I__1709 (
            .O(N__8453),
            .I(N__8450));
    LocalMux I__1708 (
            .O(N__8450),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3 ));
    InMux I__1707 (
            .O(N__8447),
            .I(N__8441));
    InMux I__1706 (
            .O(N__8446),
            .I(N__8441));
    LocalMux I__1705 (
            .O(N__8441),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ));
    InMux I__1704 (
            .O(N__8438),
            .I(N__8435));
    LocalMux I__1703 (
            .O(N__8435),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ));
    InMux I__1702 (
            .O(N__8432),
            .I(N__8426));
    InMux I__1701 (
            .O(N__8431),
            .I(N__8426));
    LocalMux I__1700 (
            .O(N__8426),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ));
    InMux I__1699 (
            .O(N__8423),
            .I(N__8420));
    LocalMux I__1698 (
            .O(N__8420),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    CascadeMux I__1697 (
            .O(N__8417),
            .I(\U712_CHIP_RAM.m159_xx_mm_0_0_cascade_ ));
    InMux I__1696 (
            .O(N__8414),
            .I(N__8411));
    LocalMux I__1695 (
            .O(N__8411),
            .I(N__8408));
    Span4Mux_v I__1694 (
            .O(N__8408),
            .I(N__8405));
    Span4Mux_v I__1693 (
            .O(N__8405),
            .I(N__8402));
    Sp12to4 I__1692 (
            .O(N__8402),
            .I(N__8399));
    Span12Mux_h I__1691 (
            .O(N__8399),
            .I(N__8396));
    Odrv12 I__1690 (
            .O(N__8396),
            .I(A_c_15));
    CascadeMux I__1689 (
            .O(N__8393),
            .I(N__8390));
    InMux I__1688 (
            .O(N__8390),
            .I(N__8387));
    LocalMux I__1687 (
            .O(N__8387),
            .I(\U712_CHIP_RAM.m156_xx_mm_0_2 ));
    IoInMux I__1686 (
            .O(N__8384),
            .I(N__8381));
    LocalMux I__1685 (
            .O(N__8381),
            .I(N__8378));
    Span4Mux_s2_v I__1684 (
            .O(N__8378),
            .I(N__8375));
    Sp12to4 I__1683 (
            .O(N__8375),
            .I(N__8372));
    Span12Mux_h I__1682 (
            .O(N__8372),
            .I(N__8369));
    Odrv12 I__1681 (
            .O(N__8369),
            .I(CMA_c_0));
    InMux I__1680 (
            .O(N__8366),
            .I(N__8363));
    LocalMux I__1679 (
            .O(N__8363),
            .I(N__8358));
    InMux I__1678 (
            .O(N__8362),
            .I(N__8355));
    CascadeMux I__1677 (
            .O(N__8361),
            .I(N__8351));
    Span4Mux_v I__1676 (
            .O(N__8358),
            .I(N__8345));
    LocalMux I__1675 (
            .O(N__8355),
            .I(N__8345));
    InMux I__1674 (
            .O(N__8354),
            .I(N__8342));
    InMux I__1673 (
            .O(N__8351),
            .I(N__8339));
    InMux I__1672 (
            .O(N__8350),
            .I(N__8336));
    Span4Mux_h I__1671 (
            .O(N__8345),
            .I(N__8333));
    LocalMux I__1670 (
            .O(N__8342),
            .I(N__8330));
    LocalMux I__1669 (
            .O(N__8339),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1668 (
            .O(N__8336),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1667 (
            .O(N__8333),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1666 (
            .O(N__8330),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1665 (
            .O(N__8321),
            .I(N__8317));
    InMux I__1664 (
            .O(N__8320),
            .I(N__8314));
    LocalMux I__1663 (
            .O(N__8317),
            .I(N__8311));
    LocalMux I__1662 (
            .O(N__8314),
            .I(N__8308));
    Span12Mux_s4_v I__1661 (
            .O(N__8311),
            .I(N__8305));
    Span4Mux_v I__1660 (
            .O(N__8308),
            .I(N__8302));
    Span12Mux_v I__1659 (
            .O(N__8305),
            .I(N__8299));
    Sp12to4 I__1658 (
            .O(N__8302),
            .I(N__8296));
    Span12Mux_h I__1657 (
            .O(N__8299),
            .I(N__8293));
    Span12Mux_h I__1656 (
            .O(N__8296),
            .I(N__8290));
    Odrv12 I__1655 (
            .O(N__8293),
            .I(A_c_9));
    Odrv12 I__1654 (
            .O(N__8290),
            .I(A_c_9));
    CascadeMux I__1653 (
            .O(N__8285),
            .I(\U712_CHIP_RAM.N_3_0_cascade_ ));
    CascadeMux I__1652 (
            .O(N__8282),
            .I(N__8279));
    InMux I__1651 (
            .O(N__8279),
            .I(N__8276));
    LocalMux I__1650 (
            .O(N__8276),
            .I(\U712_CHIP_RAM.m156_xx_mm_0_0 ));
    IoInMux I__1649 (
            .O(N__8273),
            .I(N__8270));
    LocalMux I__1648 (
            .O(N__8270),
            .I(N__8267));
    IoSpan4Mux I__1647 (
            .O(N__8267),
            .I(N__8263));
    InMux I__1646 (
            .O(N__8266),
            .I(N__8260));
    Span4Mux_s2_v I__1645 (
            .O(N__8263),
            .I(N__8257));
    LocalMux I__1644 (
            .O(N__8260),
            .I(N__8254));
    Span4Mux_v I__1643 (
            .O(N__8257),
            .I(N__8251));
    Span4Mux_v I__1642 (
            .O(N__8254),
            .I(N__8248));
    Span4Mux_v I__1641 (
            .O(N__8251),
            .I(N__8243));
    Span4Mux_v I__1640 (
            .O(N__8248),
            .I(N__8243));
    Odrv4 I__1639 (
            .O(N__8243),
            .I(N_144_0));
    IoInMux I__1638 (
            .O(N__8240),
            .I(N__8237));
    LocalMux I__1637 (
            .O(N__8237),
            .I(N__8234));
    Span4Mux_s3_h I__1636 (
            .O(N__8234),
            .I(N__8231));
    Sp12to4 I__1635 (
            .O(N__8231),
            .I(N__8228));
    Span12Mux_v I__1634 (
            .O(N__8228),
            .I(N__8225));
    Span12Mux_h I__1633 (
            .O(N__8225),
            .I(N__8222));
    Odrv12 I__1632 (
            .O(N__8222),
            .I(CLMBEn_c));
    CascadeMux I__1631 (
            .O(N__8219),
            .I(N__8216));
    InMux I__1630 (
            .O(N__8216),
            .I(N__8212));
    InMux I__1629 (
            .O(N__8215),
            .I(N__8209));
    LocalMux I__1628 (
            .O(N__8212),
            .I(N__8206));
    LocalMux I__1627 (
            .O(N__8209),
            .I(N__8203));
    Span12Mux_h I__1626 (
            .O(N__8206),
            .I(N__8200));
    Span4Mux_v I__1625 (
            .O(N__8203),
            .I(N__8197));
    Odrv12 I__1624 (
            .O(N__8200),
            .I(DBRn_c_i));
    Odrv4 I__1623 (
            .O(N__8197),
            .I(DBRn_c_i));
    InMux I__1622 (
            .O(N__8192),
            .I(N__8188));
    InMux I__1621 (
            .O(N__8191),
            .I(N__8185));
    LocalMux I__1620 (
            .O(N__8188),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    LocalMux I__1619 (
            .O(N__8185),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    InMux I__1618 (
            .O(N__8180),
            .I(N__8172));
    InMux I__1617 (
            .O(N__8179),
            .I(N__8172));
    InMux I__1616 (
            .O(N__8178),
            .I(N__8169));
    InMux I__1615 (
            .O(N__8177),
            .I(N__8166));
    LocalMux I__1614 (
            .O(N__8172),
            .I(U712_REG_SM_WRITE_CYCLE));
    LocalMux I__1613 (
            .O(N__8169),
            .I(U712_REG_SM_WRITE_CYCLE));
    LocalMux I__1612 (
            .O(N__8166),
            .I(U712_REG_SM_WRITE_CYCLE));
    CascadeMux I__1611 (
            .O(N__8159),
            .I(N__8156));
    InMux I__1610 (
            .O(N__8156),
            .I(N__8153));
    LocalMux I__1609 (
            .O(N__8153),
            .I(N_20_0));
    IoInMux I__1608 (
            .O(N__8150),
            .I(N__8147));
    LocalMux I__1607 (
            .O(N__8147),
            .I(N__8144));
    IoSpan4Mux I__1606 (
            .O(N__8144),
            .I(N__8141));
    Sp12to4 I__1605 (
            .O(N__8141),
            .I(N__8138));
    Span12Mux_v I__1604 (
            .O(N__8138),
            .I(N__8134));
    InMux I__1603 (
            .O(N__8137),
            .I(N__8131));
    Odrv12 I__1602 (
            .O(N__8134),
            .I(PRnW_c));
    LocalMux I__1601 (
            .O(N__8131),
            .I(PRnW_c));
    InMux I__1600 (
            .O(N__8126),
            .I(N__8120));
    InMux I__1599 (
            .O(N__8125),
            .I(N__8117));
    CascadeMux I__1598 (
            .O(N__8124),
            .I(N__8114));
    CascadeMux I__1597 (
            .O(N__8123),
            .I(N__8110));
    LocalMux I__1596 (
            .O(N__8120),
            .I(N__8101));
    LocalMux I__1595 (
            .O(N__8117),
            .I(N__8101));
    InMux I__1594 (
            .O(N__8114),
            .I(N__8098));
    CascadeMux I__1593 (
            .O(N__8113),
            .I(N__8091));
    InMux I__1592 (
            .O(N__8110),
            .I(N__8088));
    InMux I__1591 (
            .O(N__8109),
            .I(N__8085));
    InMux I__1590 (
            .O(N__8108),
            .I(N__8078));
    InMux I__1589 (
            .O(N__8107),
            .I(N__8078));
    InMux I__1588 (
            .O(N__8106),
            .I(N__8078));
    Span4Mux_v I__1587 (
            .O(N__8101),
            .I(N__8073));
    LocalMux I__1586 (
            .O(N__8098),
            .I(N__8073));
    InMux I__1585 (
            .O(N__8097),
            .I(N__8068));
    InMux I__1584 (
            .O(N__8096),
            .I(N__8068));
    InMux I__1583 (
            .O(N__8095),
            .I(N__8061));
    InMux I__1582 (
            .O(N__8094),
            .I(N__8061));
    InMux I__1581 (
            .O(N__8091),
            .I(N__8061));
    LocalMux I__1580 (
            .O(N__8088),
            .I(U712_REG_SM_C3_SYNC_1));
    LocalMux I__1579 (
            .O(N__8085),
            .I(U712_REG_SM_C3_SYNC_1));
    LocalMux I__1578 (
            .O(N__8078),
            .I(U712_REG_SM_C3_SYNC_1));
    Odrv4 I__1577 (
            .O(N__8073),
            .I(U712_REG_SM_C3_SYNC_1));
    LocalMux I__1576 (
            .O(N__8068),
            .I(U712_REG_SM_C3_SYNC_1));
    LocalMux I__1575 (
            .O(N__8061),
            .I(U712_REG_SM_C3_SYNC_1));
    IoInMux I__1574 (
            .O(N__8048),
            .I(N__8045));
    LocalMux I__1573 (
            .O(N__8045),
            .I(N__8041));
    IoInMux I__1572 (
            .O(N__8044),
            .I(N__8038));
    Span4Mux_s1_v I__1571 (
            .O(N__8041),
            .I(N__8035));
    LocalMux I__1570 (
            .O(N__8038),
            .I(N__8032));
    Span4Mux_v I__1569 (
            .O(N__8035),
            .I(N__8029));
    Span12Mux_s11_v I__1568 (
            .O(N__8032),
            .I(N__8026));
    Sp12to4 I__1567 (
            .O(N__8029),
            .I(N__8023));
    Span12Mux_h I__1566 (
            .O(N__8026),
            .I(N__8020));
    Span12Mux_h I__1565 (
            .O(N__8023),
            .I(N__8017));
    Odrv12 I__1564 (
            .O(N__8020),
            .I(BLSn_c));
    Odrv12 I__1563 (
            .O(N__8017),
            .I(BLSn_c));
    CEMux I__1562 (
            .O(N__8012),
            .I(N__8009));
    LocalMux I__1561 (
            .O(N__8009),
            .I(N__8006));
    Span4Mux_v I__1560 (
            .O(N__8006),
            .I(N__8003));
    Odrv4 I__1559 (
            .O(N__8003),
            .I(\U712_REG_SM.N_20_0_0 ));
    InMux I__1558 (
            .O(N__8000),
            .I(N__7997));
    LocalMux I__1557 (
            .O(N__7997),
            .I(N_172_0));
    IoInMux I__1556 (
            .O(N__7994),
            .I(N__7991));
    LocalMux I__1555 (
            .O(N__7991),
            .I(N__7988));
    Span12Mux_s1_v I__1554 (
            .O(N__7988),
            .I(N__7985));
    Span12Mux_h I__1553 (
            .O(N__7985),
            .I(N__7981));
    InMux I__1552 (
            .O(N__7984),
            .I(N__7978));
    Odrv12 I__1551 (
            .O(N__7981),
            .I(LDSn_c));
    LocalMux I__1550 (
            .O(N__7978),
            .I(LDSn_c));
    IoInMux I__1549 (
            .O(N__7973),
            .I(N__7970));
    LocalMux I__1548 (
            .O(N__7970),
            .I(N__7967));
    Span12Mux_s3_v I__1547 (
            .O(N__7967),
            .I(N__7964));
    Odrv12 I__1546 (
            .O(N__7964),
            .I(RESETn_c_i));
    IoInMux I__1545 (
            .O(N__7961),
            .I(N__7958));
    LocalMux I__1544 (
            .O(N__7958),
            .I(N__7955));
    IoSpan4Mux I__1543 (
            .O(N__7955),
            .I(N__7952));
    IoSpan4Mux I__1542 (
            .O(N__7952),
            .I(N__7949));
    Span4Mux_s2_h I__1541 (
            .O(N__7949),
            .I(N__7946));
    Sp12to4 I__1540 (
            .O(N__7946),
            .I(N__7943));
    Span12Mux_h I__1539 (
            .O(N__7943),
            .I(N__7940));
    Odrv12 I__1538 (
            .O(N__7940),
            .I(WEn_c));
    InMux I__1537 (
            .O(N__7937),
            .I(N__7934));
    LocalMux I__1536 (
            .O(N__7934),
            .I(N__7931));
    Sp12to4 I__1535 (
            .O(N__7931),
            .I(N__7928));
    Span12Mux_v I__1534 (
            .O(N__7928),
            .I(N__7925));
    Span12Mux_h I__1533 (
            .O(N__7925),
            .I(N__7922));
    Odrv12 I__1532 (
            .O(N__7922),
            .I(A_c_16));
    InMux I__1531 (
            .O(N__7919),
            .I(N__7916));
    LocalMux I__1530 (
            .O(N__7916),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    CascadeMux I__1529 (
            .O(N__7913),
            .I(\U712_CHIP_RAM.m161_xx_mm_0_0_cascade_ ));
    InMux I__1528 (
            .O(N__7910),
            .I(N__7907));
    LocalMux I__1527 (
            .O(N__7907),
            .I(N__7904));
    Span4Mux_v I__1526 (
            .O(N__7904),
            .I(N__7901));
    Sp12to4 I__1525 (
            .O(N__7901),
            .I(N__7898));
    Span12Mux_h I__1524 (
            .O(N__7898),
            .I(N__7895));
    Odrv12 I__1523 (
            .O(N__7895),
            .I(A_c_13));
    InMux I__1522 (
            .O(N__7892),
            .I(N__7889));
    LocalMux I__1521 (
            .O(N__7889),
            .I(N__7886));
    Span12Mux_v I__1520 (
            .O(N__7886),
            .I(N__7883));
    Span12Mux_h I__1519 (
            .O(N__7883),
            .I(N__7880));
    Odrv12 I__1518 (
            .O(N__7880),
            .I(A_c_17));
    InMux I__1517 (
            .O(N__7877),
            .I(N__7874));
    LocalMux I__1516 (
            .O(N__7874),
            .I(N__7871));
    Span4Mux_h I__1515 (
            .O(N__7871),
            .I(N__7868));
    Odrv4 I__1514 (
            .O(N__7868),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8 ));
    CascadeMux I__1513 (
            .O(N__7865),
            .I(\U712_CHIP_RAM.m162_xx_mm_0_0_cascade_ ));
    CascadeMux I__1512 (
            .O(N__7862),
            .I(\U712_CHIP_RAM.m162_xx_mm_0_2_cascade_ ));
    IoInMux I__1511 (
            .O(N__7859),
            .I(N__7856));
    LocalMux I__1510 (
            .O(N__7856),
            .I(N__7853));
    IoSpan4Mux I__1509 (
            .O(N__7853),
            .I(N__7850));
    Span4Mux_s3_h I__1508 (
            .O(N__7850),
            .I(N__7847));
    Span4Mux_v I__1507 (
            .O(N__7847),
            .I(N__7844));
    Span4Mux_v I__1506 (
            .O(N__7844),
            .I(N__7841));
    Sp12to4 I__1505 (
            .O(N__7841),
            .I(N__7838));
    Odrv12 I__1504 (
            .O(N__7838),
            .I(CMA_c_8));
    InMux I__1503 (
            .O(N__7835),
            .I(N__7832));
    LocalMux I__1502 (
            .O(N__7832),
            .I(U712_CHIP_RAM_m45_0));
    InMux I__1501 (
            .O(N__7829),
            .I(N__7826));
    LocalMux I__1500 (
            .O(N__7826),
            .I(N__7822));
    InMux I__1499 (
            .O(N__7825),
            .I(N__7819));
    Odrv4 I__1498 (
            .O(N__7822),
            .I(REG_TACK));
    LocalMux I__1497 (
            .O(N__7819),
            .I(REG_TACK));
    InMux I__1496 (
            .O(N__7814),
            .I(N__7811));
    LocalMux I__1495 (
            .O(N__7811),
            .I(U712_REG_SM_REG_TACK_7_0));
    CascadeMux I__1494 (
            .O(N__7808),
            .I(N__7805));
    InMux I__1493 (
            .O(N__7805),
            .I(N__7797));
    InMux I__1492 (
            .O(N__7804),
            .I(N__7792));
    InMux I__1491 (
            .O(N__7803),
            .I(N__7792));
    InMux I__1490 (
            .O(N__7802),
            .I(N__7785));
    InMux I__1489 (
            .O(N__7801),
            .I(N__7785));
    InMux I__1488 (
            .O(N__7800),
            .I(N__7785));
    LocalMux I__1487 (
            .O(N__7797),
            .I(U712_REG_SM_STATE_COUNT_8));
    LocalMux I__1486 (
            .O(N__7792),
            .I(U712_REG_SM_STATE_COUNT_8));
    LocalMux I__1485 (
            .O(N__7785),
            .I(U712_REG_SM_STATE_COUNT_8));
    InMux I__1484 (
            .O(N__7778),
            .I(N__7770));
    InMux I__1483 (
            .O(N__7777),
            .I(N__7770));
    InMux I__1482 (
            .O(N__7776),
            .I(N__7765));
    InMux I__1481 (
            .O(N__7775),
            .I(N__7765));
    LocalMux I__1480 (
            .O(N__7770),
            .I(U712_REG_SM_STATE_COUNT_3));
    LocalMux I__1479 (
            .O(N__7765),
            .I(U712_REG_SM_STATE_COUNT_3));
    CascadeMux I__1478 (
            .O(N__7760),
            .I(N__7757));
    InMux I__1477 (
            .O(N__7757),
            .I(N__7754));
    LocalMux I__1476 (
            .O(N__7754),
            .I(N_44_0));
    InMux I__1475 (
            .O(N__7751),
            .I(N__7747));
    InMux I__1474 (
            .O(N__7750),
            .I(N__7743));
    LocalMux I__1473 (
            .O(N__7747),
            .I(N__7740));
    InMux I__1472 (
            .O(N__7746),
            .I(N__7737));
    LocalMux I__1471 (
            .O(N__7743),
            .I(N_175_0));
    Odrv4 I__1470 (
            .O(N__7740),
            .I(N_175_0));
    LocalMux I__1469 (
            .O(N__7737),
            .I(N_175_0));
    InMux I__1468 (
            .O(N__7730),
            .I(N__7726));
    InMux I__1467 (
            .O(N__7729),
            .I(N__7723));
    LocalMux I__1466 (
            .O(N__7726),
            .I(N__7720));
    LocalMux I__1465 (
            .O(N__7723),
            .I(N__7717));
    Span4Mux_v I__1464 (
            .O(N__7720),
            .I(N__7714));
    Span4Mux_v I__1463 (
            .O(N__7717),
            .I(N__7711));
    Sp12to4 I__1462 (
            .O(N__7714),
            .I(N__7706));
    Sp12to4 I__1461 (
            .O(N__7711),
            .I(N__7706));
    Span12Mux_h I__1460 (
            .O(N__7706),
            .I(N__7703));
    Odrv12 I__1459 (
            .O(N__7703),
            .I(DBRn_c));
    InMux I__1458 (
            .O(N__7700),
            .I(N__7697));
    LocalMux I__1457 (
            .O(N__7697),
            .I(DBR_SYNCZ0Z_0));
    IoInMux I__1456 (
            .O(N__7694),
            .I(N__7691));
    LocalMux I__1455 (
            .O(N__7691),
            .I(N__7688));
    Span12Mux_s8_v I__1454 (
            .O(N__7688),
            .I(N__7685));
    Odrv12 I__1453 (
            .O(N__7685),
            .I(CMA_c_1));
    InMux I__1452 (
            .O(N__7682),
            .I(N__7679));
    LocalMux I__1451 (
            .O(N__7679),
            .I(\U712_CHIP_RAM.m154_0_2 ));
    InMux I__1450 (
            .O(N__7676),
            .I(N__7673));
    LocalMux I__1449 (
            .O(N__7673),
            .I(N__7669));
    InMux I__1448 (
            .O(N__7672),
            .I(N__7666));
    Span4Mux_h I__1447 (
            .O(N__7669),
            .I(N__7663));
    LocalMux I__1446 (
            .O(N__7666),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ));
    Odrv4 I__1445 (
            .O(N__7663),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ));
    InMux I__1444 (
            .O(N__7658),
            .I(N__7655));
    LocalMux I__1443 (
            .O(N__7655),
            .I(\U712_CHIP_RAM.m154_0_0 ));
    IoInMux I__1442 (
            .O(N__7652),
            .I(N__7649));
    LocalMux I__1441 (
            .O(N__7649),
            .I(N__7646));
    Span4Mux_s0_v I__1440 (
            .O(N__7646),
            .I(N__7643));
    Span4Mux_v I__1439 (
            .O(N__7643),
            .I(N__7639));
    InMux I__1438 (
            .O(N__7642),
            .I(N__7636));
    Span4Mux_v I__1437 (
            .O(N__7639),
            .I(N__7633));
    LocalMux I__1436 (
            .O(N__7636),
            .I(N__7630));
    Sp12to4 I__1435 (
            .O(N__7633),
            .I(N__7627));
    Span4Mux_v I__1434 (
            .O(N__7630),
            .I(N__7624));
    Span12Mux_h I__1433 (
            .O(N__7627),
            .I(N__7621));
    Sp12to4 I__1432 (
            .O(N__7624),
            .I(N__7618));
    Span12Mux_v I__1431 (
            .O(N__7621),
            .I(N__7613));
    Span12Mux_h I__1430 (
            .O(N__7618),
            .I(N__7613));
    Odrv12 I__1429 (
            .O(N__7613),
            .I(A_c_10));
    InMux I__1428 (
            .O(N__7610),
            .I(N__7607));
    LocalMux I__1427 (
            .O(N__7607),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    IoInMux I__1426 (
            .O(N__7604),
            .I(N__7601));
    LocalMux I__1425 (
            .O(N__7601),
            .I(N__7598));
    IoSpan4Mux I__1424 (
            .O(N__7598),
            .I(N__7595));
    Span4Mux_s2_v I__1423 (
            .O(N__7595),
            .I(N__7592));
    Sp12to4 I__1422 (
            .O(N__7592),
            .I(N__7588));
    InMux I__1421 (
            .O(N__7591),
            .I(N__7585));
    Span12Mux_s8_v I__1420 (
            .O(N__7588),
            .I(N__7582));
    LocalMux I__1419 (
            .O(N__7585),
            .I(N__7579));
    Span12Mux_v I__1418 (
            .O(N__7582),
            .I(N__7576));
    Span12Mux_v I__1417 (
            .O(N__7579),
            .I(N__7573));
    Span12Mux_h I__1416 (
            .O(N__7576),
            .I(N__7570));
    Span12Mux_h I__1415 (
            .O(N__7573),
            .I(N__7567));
    Odrv12 I__1414 (
            .O(N__7570),
            .I(A_c_11));
    Odrv12 I__1413 (
            .O(N__7567),
            .I(A_c_11));
    InMux I__1412 (
            .O(N__7562),
            .I(N__7559));
    LocalMux I__1411 (
            .O(N__7559),
            .I(N__7556));
    Span4Mux_v I__1410 (
            .O(N__7556),
            .I(N__7553));
    Odrv4 I__1409 (
            .O(N__7553),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    CascadeMux I__1408 (
            .O(N__7550),
            .I(\U712_CHIP_RAM.m157_xx_mm_0_0_cascade_ ));
    InMux I__1407 (
            .O(N__7547),
            .I(N__7544));
    LocalMux I__1406 (
            .O(N__7544),
            .I(\U712_CHIP_RAM.m157_xx_mm_0_2 ));
    InMux I__1405 (
            .O(N__7541),
            .I(N__7538));
    LocalMux I__1404 (
            .O(N__7538),
            .I(N__7535));
    Odrv4 I__1403 (
            .O(N__7535),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    InMux I__1402 (
            .O(N__7532),
            .I(N__7528));
    InMux I__1401 (
            .O(N__7531),
            .I(N__7525));
    LocalMux I__1400 (
            .O(N__7528),
            .I(N__7522));
    LocalMux I__1399 (
            .O(N__7525),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ));
    Odrv12 I__1398 (
            .O(N__7522),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ));
    InMux I__1397 (
            .O(N__7517),
            .I(N__7513));
    InMux I__1396 (
            .O(N__7516),
            .I(N__7510));
    LocalMux I__1395 (
            .O(N__7513),
            .I(N__7507));
    LocalMux I__1394 (
            .O(N__7510),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ));
    Odrv12 I__1393 (
            .O(N__7507),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ));
    InMux I__1392 (
            .O(N__7502),
            .I(N__7498));
    InMux I__1391 (
            .O(N__7501),
            .I(N__7495));
    LocalMux I__1390 (
            .O(N__7498),
            .I(U712_REG_SM_STATE_COUNT_2));
    LocalMux I__1389 (
            .O(N__7495),
            .I(U712_REG_SM_STATE_COUNT_2));
    InMux I__1388 (
            .O(N__7490),
            .I(N__7484));
    InMux I__1387 (
            .O(N__7489),
            .I(N__7484));
    LocalMux I__1386 (
            .O(N__7484),
            .I(\U712_CHIP_RAM.N_37_0 ));
    InMux I__1385 (
            .O(N__7481),
            .I(N__7478));
    LocalMux I__1384 (
            .O(N__7478),
            .I(N_174_0));
    IoInMux I__1383 (
            .O(N__7475),
            .I(N__7472));
    LocalMux I__1382 (
            .O(N__7472),
            .I(N__7469));
    Span12Mux_s5_v I__1381 (
            .O(N__7469),
            .I(N__7466));
    Span12Mux_h I__1380 (
            .O(N__7466),
            .I(N__7462));
    InMux I__1379 (
            .O(N__7465),
            .I(N__7459));
    Odrv12 I__1378 (
            .O(N__7462),
            .I(UDSn_c));
    LocalMux I__1377 (
            .O(N__7459),
            .I(UDSn_c));
    InMux I__1376 (
            .O(N__7454),
            .I(N__7449));
    InMux I__1375 (
            .O(N__7453),
            .I(N__7446));
    InMux I__1374 (
            .O(N__7452),
            .I(N__7443));
    LocalMux I__1373 (
            .O(N__7449),
            .I(N__7437));
    LocalMux I__1372 (
            .O(N__7446),
            .I(N__7432));
    LocalMux I__1371 (
            .O(N__7443),
            .I(N__7432));
    InMux I__1370 (
            .O(N__7442),
            .I(N__7429));
    InMux I__1369 (
            .O(N__7441),
            .I(N__7426));
    CascadeMux I__1368 (
            .O(N__7440),
            .I(N__7423));
    Span4Mux_v I__1367 (
            .O(N__7437),
            .I(N__7414));
    Span4Mux_h I__1366 (
            .O(N__7432),
            .I(N__7414));
    LocalMux I__1365 (
            .O(N__7429),
            .I(N__7414));
    LocalMux I__1364 (
            .O(N__7426),
            .I(N__7414));
    InMux I__1363 (
            .O(N__7423),
            .I(N__7411));
    Span4Mux_h I__1362 (
            .O(N__7414),
            .I(N__7406));
    LocalMux I__1361 (
            .O(N__7411),
            .I(N__7406));
    Span4Mux_v I__1360 (
            .O(N__7406),
            .I(N__7403));
    Span4Mux_v I__1359 (
            .O(N__7403),
            .I(N__7400));
    Sp12to4 I__1358 (
            .O(N__7400),
            .I(N__7397));
    Span12Mux_h I__1357 (
            .O(N__7397),
            .I(N__7394));
    Odrv12 I__1356 (
            .O(N__7394),
            .I(SIZ_c_0));
    CascadeMux I__1355 (
            .O(N__7391),
            .I(N__7386));
    CascadeMux I__1354 (
            .O(N__7390),
            .I(N__7383));
    InMux I__1353 (
            .O(N__7389),
            .I(N__7376));
    InMux I__1352 (
            .O(N__7386),
            .I(N__7376));
    InMux I__1351 (
            .O(N__7383),
            .I(N__7376));
    LocalMux I__1350 (
            .O(N__7376),
            .I(N__7373));
    Odrv12 I__1349 (
            .O(N__7373),
            .I(\U712_CHIP_RAM.N_326_mux ));
    CascadeMux I__1348 (
            .O(N__7370),
            .I(N__7367));
    InMux I__1347 (
            .O(N__7367),
            .I(N__7359));
    InMux I__1346 (
            .O(N__7366),
            .I(N__7359));
    InMux I__1345 (
            .O(N__7365),
            .I(N__7356));
    InMux I__1344 (
            .O(N__7364),
            .I(N__7353));
    LocalMux I__1343 (
            .O(N__7359),
            .I(N__7346));
    LocalMux I__1342 (
            .O(N__7356),
            .I(N__7346));
    LocalMux I__1341 (
            .O(N__7353),
            .I(N__7346));
    Span4Mux_v I__1340 (
            .O(N__7346),
            .I(N__7343));
    Sp12to4 I__1339 (
            .O(N__7343),
            .I(N__7340));
    Span12Mux_h I__1338 (
            .O(N__7340),
            .I(N__7337));
    Odrv12 I__1337 (
            .O(N__7337),
            .I(A_c_1));
    InMux I__1336 (
            .O(N__7334),
            .I(N__7330));
    InMux I__1335 (
            .O(N__7333),
            .I(N__7327));
    LocalMux I__1334 (
            .O(N__7330),
            .I(N__7324));
    LocalMux I__1333 (
            .O(N__7327),
            .I(N__7321));
    Span4Mux_h I__1332 (
            .O(N__7324),
            .I(N__7313));
    Span4Mux_h I__1331 (
            .O(N__7321),
            .I(N__7313));
    InMux I__1330 (
            .O(N__7320),
            .I(N__7310));
    InMux I__1329 (
            .O(N__7319),
            .I(N__7307));
    InMux I__1328 (
            .O(N__7318),
            .I(N__7304));
    Span4Mux_v I__1327 (
            .O(N__7313),
            .I(N__7300));
    LocalMux I__1326 (
            .O(N__7310),
            .I(N__7293));
    LocalMux I__1325 (
            .O(N__7307),
            .I(N__7293));
    LocalMux I__1324 (
            .O(N__7304),
            .I(N__7293));
    InMux I__1323 (
            .O(N__7303),
            .I(N__7290));
    Span4Mux_v I__1322 (
            .O(N__7300),
            .I(N__7287));
    Sp12to4 I__1321 (
            .O(N__7293),
            .I(N__7282));
    LocalMux I__1320 (
            .O(N__7290),
            .I(N__7282));
    Sp12to4 I__1319 (
            .O(N__7287),
            .I(N__7277));
    Span12Mux_v I__1318 (
            .O(N__7282),
            .I(N__7277));
    Span12Mux_h I__1317 (
            .O(N__7277),
            .I(N__7274));
    Odrv12 I__1316 (
            .O(N__7274),
            .I(SIZ_c_1));
    IoInMux I__1315 (
            .O(N__7271),
            .I(N__7268));
    LocalMux I__1314 (
            .O(N__7268),
            .I(N__7264));
    InMux I__1313 (
            .O(N__7267),
            .I(N__7261));
    IoSpan4Mux I__1312 (
            .O(N__7264),
            .I(N__7258));
    LocalMux I__1311 (
            .O(N__7261),
            .I(N__7255));
    IoSpan4Mux I__1310 (
            .O(N__7258),
            .I(N__7252));
    Span12Mux_h I__1309 (
            .O(N__7255),
            .I(N__7249));
    IoSpan4Mux I__1308 (
            .O(N__7252),
            .I(N__7246));
    Odrv12 I__1307 (
            .O(N__7249),
            .I(C1_c));
    Odrv4 I__1306 (
            .O(N__7246),
            .I(C1_c));
    InMux I__1305 (
            .O(N__7241),
            .I(N__7238));
    LocalMux I__1304 (
            .O(N__7238),
            .I(N__7235));
    Odrv4 I__1303 (
            .O(N__7235),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    ClkMux I__1302 (
            .O(N__7232),
            .I(N__7228));
    ClkMux I__1301 (
            .O(N__7231),
            .I(N__7225));
    LocalMux I__1300 (
            .O(N__7228),
            .I(N__7222));
    LocalMux I__1299 (
            .O(N__7225),
            .I(N__7219));
    Span4Mux_h I__1298 (
            .O(N__7222),
            .I(N__7216));
    Span4Mux_v I__1297 (
            .O(N__7219),
            .I(N__7213));
    Span4Mux_v I__1296 (
            .O(N__7216),
            .I(N__7210));
    Sp12to4 I__1295 (
            .O(N__7213),
            .I(N__7206));
    Span4Mux_v I__1294 (
            .O(N__7210),
            .I(N__7203));
    InMux I__1293 (
            .O(N__7209),
            .I(N__7200));
    Span12Mux_h I__1292 (
            .O(N__7206),
            .I(N__7197));
    Span4Mux_v I__1291 (
            .O(N__7203),
            .I(N__7192));
    LocalMux I__1290 (
            .O(N__7200),
            .I(N__7192));
    Span12Mux_v I__1289 (
            .O(N__7197),
            .I(N__7189));
    Span4Mux_v I__1288 (
            .O(N__7192),
            .I(N__7186));
    Odrv12 I__1287 (
            .O(N__7189),
            .I(CLK40_PLL));
    Odrv4 I__1286 (
            .O(N__7186),
            .I(CLK40_PLL));
    IoInMux I__1285 (
            .O(N__7181),
            .I(N__7177));
    IoInMux I__1284 (
            .O(N__7180),
            .I(N__7173));
    LocalMux I__1283 (
            .O(N__7177),
            .I(N__7170));
    IoInMux I__1282 (
            .O(N__7176),
            .I(N__7167));
    LocalMux I__1281 (
            .O(N__7173),
            .I(N__7164));
    Span4Mux_s1_v I__1280 (
            .O(N__7170),
            .I(N__7161));
    LocalMux I__1279 (
            .O(N__7167),
            .I(N__7158));
    Span12Mux_s1_v I__1278 (
            .O(N__7164),
            .I(N__7155));
    Sp12to4 I__1277 (
            .O(N__7161),
            .I(N__7152));
    Span4Mux_s2_h I__1276 (
            .O(N__7158),
            .I(N__7149));
    Span12Mux_h I__1275 (
            .O(N__7155),
            .I(N__7146));
    Span12Mux_h I__1274 (
            .O(N__7152),
            .I(N__7143));
    Sp12to4 I__1273 (
            .O(N__7149),
            .I(N__7140));
    Span12Mux_v I__1272 (
            .O(N__7146),
            .I(N__7137));
    Span12Mux_v I__1271 (
            .O(N__7143),
            .I(N__7134));
    Span12Mux_v I__1270 (
            .O(N__7140),
            .I(N__7131));
    Span12Mux_v I__1269 (
            .O(N__7137),
            .I(N__7128));
    Span12Mux_v I__1268 (
            .O(N__7134),
            .I(N__7123));
    Span12Mux_h I__1267 (
            .O(N__7131),
            .I(N__7123));
    Odrv12 I__1266 (
            .O(N__7128),
            .I(CLK40_PLL_iso_i));
    Odrv12 I__1265 (
            .O(N__7123),
            .I(CLK40_PLL_iso_i));
    CascadeMux I__1264 (
            .O(N__7118),
            .I(i66_mux_cascade_));
    InMux I__1263 (
            .O(N__7115),
            .I(N__7112));
    LocalMux I__1262 (
            .O(N__7112),
            .I(\U712_CHIP_RAM.m40_nsZ0Z_1 ));
    InMux I__1261 (
            .O(N__7109),
            .I(N__7106));
    LocalMux I__1260 (
            .O(N__7106),
            .I(N_10_0));
    InMux I__1259 (
            .O(N__7103),
            .I(N__7100));
    LocalMux I__1258 (
            .O(N__7100),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    CascadeMux I__1257 (
            .O(N__7097),
            .I(N__7094));
    InMux I__1256 (
            .O(N__7094),
            .I(N__7091));
    LocalMux I__1255 (
            .O(N__7091),
            .I(N__7088));
    Odrv4 I__1254 (
            .O(N__7088),
            .I(U712_REG_SM_STATE_COUNT_7));
    InMux I__1253 (
            .O(N__7085),
            .I(N__7082));
    LocalMux I__1252 (
            .O(N__7082),
            .I(\U712_CHIP_RAM.N_21_0 ));
    CascadeMux I__1251 (
            .O(N__7079),
            .I(\U712_CHIP_RAM.N_21_0_cascade_ ));
    InMux I__1250 (
            .O(N__7076),
            .I(N__7073));
    LocalMux I__1249 (
            .O(N__7073),
            .I(\U712_CHIP_RAM.N_31_0 ));
    InMux I__1248 (
            .O(N__7070),
            .I(N__7067));
    LocalMux I__1247 (
            .O(N__7067),
            .I(\U712_CHIP_RAM.N_329 ));
    CascadeMux I__1246 (
            .O(N__7064),
            .I(N__7058));
    InMux I__1245 (
            .O(N__7063),
            .I(N__7052));
    InMux I__1244 (
            .O(N__7062),
            .I(N__7052));
    InMux I__1243 (
            .O(N__7061),
            .I(N__7049));
    InMux I__1242 (
            .O(N__7058),
            .I(N__7044));
    InMux I__1241 (
            .O(N__7057),
            .I(N__7044));
    LocalMux I__1240 (
            .O(N__7052),
            .I(U712_REG_SM_STATE_COUNT_1));
    LocalMux I__1239 (
            .O(N__7049),
            .I(U712_REG_SM_STATE_COUNT_1));
    LocalMux I__1238 (
            .O(N__7044),
            .I(U712_REG_SM_STATE_COUNT_1));
    CascadeMux I__1237 (
            .O(N__7037),
            .I(N_20_0_cascade_));
    SRMux I__1236 (
            .O(N__7034),
            .I(N__7031));
    LocalMux I__1235 (
            .O(N__7031),
            .I(\U712_CYCLE_TERM.TACK_RST_0_i ));
    CascadeMux I__1234 (
            .O(N__7028),
            .I(N__7025));
    InMux I__1233 (
            .O(N__7025),
            .I(N__7019));
    InMux I__1232 (
            .O(N__7024),
            .I(N__7019));
    LocalMux I__1231 (
            .O(N__7019),
            .I(U712_REG_SM_STATE_COUNT_5));
    InMux I__1230 (
            .O(N__7016),
            .I(N__7013));
    LocalMux I__1229 (
            .O(N__7013),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    CascadeMux I__1228 (
            .O(N__7010),
            .I(N_10_0_cascade_));
    InMux I__1227 (
            .O(N__7007),
            .I(N__7004));
    LocalMux I__1226 (
            .O(N__7004),
            .I(N__6999));
    CascadeMux I__1225 (
            .O(N__7003),
            .I(N__6996));
    InMux I__1224 (
            .O(N__7002),
            .I(N__6992));
    Span4Mux_h I__1223 (
            .O(N__6999),
            .I(N__6989));
    InMux I__1222 (
            .O(N__6996),
            .I(N__6984));
    InMux I__1221 (
            .O(N__6995),
            .I(N__6984));
    LocalMux I__1220 (
            .O(N__6992),
            .I(U712_REG_SM_REG_CYCLE_START));
    Odrv4 I__1219 (
            .O(N__6989),
            .I(U712_REG_SM_REG_CYCLE_START));
    LocalMux I__1218 (
            .O(N__6984),
            .I(U712_REG_SM_REG_CYCLE_START));
    CascadeMux I__1217 (
            .O(N__6977),
            .I(\U712_CHIP_RAM.N_84_0_cascade_ ));
    InMux I__1216 (
            .O(N__6974),
            .I(N__6968));
    InMux I__1215 (
            .O(N__6973),
            .I(N__6965));
    InMux I__1214 (
            .O(N__6972),
            .I(N__6960));
    InMux I__1213 (
            .O(N__6971),
            .I(N__6960));
    LocalMux I__1212 (
            .O(N__6968),
            .I(U712_REG_SM_STATE_COUNT_0));
    LocalMux I__1211 (
            .O(N__6965),
            .I(U712_REG_SM_STATE_COUNT_0));
    LocalMux I__1210 (
            .O(N__6960),
            .I(U712_REG_SM_STATE_COUNT_0));
    InMux I__1209 (
            .O(N__6953),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__1208 (
            .O(N__6950),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__1207 (
            .O(N__6947),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__1206 (
            .O(N__6944),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__1205 (
            .O(N__6941),
            .I(N__6911));
    ClkMux I__1204 (
            .O(N__6940),
            .I(N__6911));
    ClkMux I__1203 (
            .O(N__6939),
            .I(N__6911));
    ClkMux I__1202 (
            .O(N__6938),
            .I(N__6911));
    ClkMux I__1201 (
            .O(N__6937),
            .I(N__6911));
    ClkMux I__1200 (
            .O(N__6936),
            .I(N__6911));
    ClkMux I__1199 (
            .O(N__6935),
            .I(N__6911));
    ClkMux I__1198 (
            .O(N__6934),
            .I(N__6911));
    ClkMux I__1197 (
            .O(N__6933),
            .I(N__6911));
    ClkMux I__1196 (
            .O(N__6932),
            .I(N__6911));
    GlobalMux I__1195 (
            .O(N__6911),
            .I(N__6908));
    gio2CtrlBuf I__1194 (
            .O(N__6908),
            .I(C1_c_g));
    SRMux I__1193 (
            .O(N__6905),
            .I(N__6902));
    LocalMux I__1192 (
            .O(N__6902),
            .I(N__6899));
    Span4Mux_h I__1191 (
            .O(N__6899),
            .I(N__6896));
    Odrv4 I__1190 (
            .O(N__6896),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__1189 (
            .O(N__6893),
            .I(N__6889));
    InMux I__1188 (
            .O(N__6892),
            .I(N__6886));
    LocalMux I__1187 (
            .O(N__6889),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__1186 (
            .O(N__6886),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__1185 (
            .O(N__6881),
            .I(N__6877));
    InMux I__1184 (
            .O(N__6880),
            .I(N__6874));
    LocalMux I__1183 (
            .O(N__6877),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__1182 (
            .O(N__6874),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    CascadeMux I__1181 (
            .O(N__6869),
            .I(N__6865));
    InMux I__1180 (
            .O(N__6868),
            .I(N__6862));
    InMux I__1179 (
            .O(N__6865),
            .I(N__6859));
    LocalMux I__1178 (
            .O(N__6862),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__1177 (
            .O(N__6859),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__1176 (
            .O(N__6854),
            .I(N__6850));
    InMux I__1175 (
            .O(N__6853),
            .I(N__6847));
    LocalMux I__1174 (
            .O(N__6850),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__1173 (
            .O(N__6847),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__1172 (
            .O(N__6842),
            .I(N__6838));
    InMux I__1171 (
            .O(N__6841),
            .I(N__6835));
    LocalMux I__1170 (
            .O(N__6838),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__1169 (
            .O(N__6835),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__1168 (
            .O(N__6830),
            .I(N__6826));
    InMux I__1167 (
            .O(N__6829),
            .I(N__6823));
    LocalMux I__1166 (
            .O(N__6826),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__1165 (
            .O(N__6823),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    CascadeMux I__1164 (
            .O(N__6818),
            .I(\U712_CHIP_RAM.REFRESH5lt7_cascade_ ));
    InMux I__1163 (
            .O(N__6815),
            .I(N__6811));
    InMux I__1162 (
            .O(N__6814),
            .I(N__6808));
    LocalMux I__1161 (
            .O(N__6811),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__1160 (
            .O(N__6808),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    CascadeMux I__1159 (
            .O(N__6803),
            .I(N__6799));
    CascadeMux I__1158 (
            .O(N__6802),
            .I(N__6795));
    InMux I__1157 (
            .O(N__6799),
            .I(N__6791));
    InMux I__1156 (
            .O(N__6798),
            .I(N__6788));
    InMux I__1155 (
            .O(N__6795),
            .I(N__6785));
    InMux I__1154 (
            .O(N__6794),
            .I(N__6782));
    LocalMux I__1153 (
            .O(N__6791),
            .I(N__6778));
    LocalMux I__1152 (
            .O(N__6788),
            .I(N__6771));
    LocalMux I__1151 (
            .O(N__6785),
            .I(N__6771));
    LocalMux I__1150 (
            .O(N__6782),
            .I(N__6771));
    InMux I__1149 (
            .O(N__6781),
            .I(N__6768));
    Span4Mux_h I__1148 (
            .O(N__6778),
            .I(N__6765));
    Span4Mux_v I__1147 (
            .O(N__6771),
            .I(N__6762));
    LocalMux I__1146 (
            .O(N__6768),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__1145 (
            .O(N__6765),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__1144 (
            .O(N__6762),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__1143 (
            .O(N__6755),
            .I(N__6752));
    LocalMux I__1142 (
            .O(N__6752),
            .I(\U712_CHIP_RAM.N_168_0 ));
    InMux I__1141 (
            .O(N__6749),
            .I(N__6746));
    LocalMux I__1140 (
            .O(N__6746),
            .I(N__6742));
    InMux I__1139 (
            .O(N__6745),
            .I(N__6739));
    Odrv4 I__1138 (
            .O(N__6742),
            .I(CPU_TACKm));
    LocalMux I__1137 (
            .O(N__6739),
            .I(CPU_TACKm));
    CascadeMux I__1136 (
            .O(N__6734),
            .I(\U712_CHIP_RAM.N_66_0_cascade_ ));
    InMux I__1135 (
            .O(N__6731),
            .I(N__6727));
    InMux I__1134 (
            .O(N__6730),
            .I(N__6724));
    LocalMux I__1133 (
            .O(N__6727),
            .I(N__6721));
    LocalMux I__1132 (
            .O(N__6724),
            .I(N__6718));
    Span4Mux_v I__1131 (
            .O(N__6721),
            .I(N__6712));
    Span4Mux_v I__1130 (
            .O(N__6718),
            .I(N__6712));
    CascadeMux I__1129 (
            .O(N__6717),
            .I(N__6709));
    Span4Mux_h I__1128 (
            .O(N__6712),
            .I(N__6705));
    InMux I__1127 (
            .O(N__6709),
            .I(N__6702));
    InMux I__1126 (
            .O(N__6708),
            .I(N__6699));
    Sp12to4 I__1125 (
            .O(N__6705),
            .I(N__6692));
    LocalMux I__1124 (
            .O(N__6702),
            .I(N__6692));
    LocalMux I__1123 (
            .O(N__6699),
            .I(N__6692));
    Span12Mux_h I__1122 (
            .O(N__6692),
            .I(N__6689));
    Odrv12 I__1121 (
            .O(N__6689),
            .I(A_c_0));
    IoInMux I__1120 (
            .O(N__6686),
            .I(N__6683));
    LocalMux I__1119 (
            .O(N__6683),
            .I(N__6680));
    Span12Mux_s5_v I__1118 (
            .O(N__6680),
            .I(N__6677));
    Odrv12 I__1117 (
            .O(N__6677),
            .I(CMA_c_2));
    InMux I__1116 (
            .O(N__6674),
            .I(N__6671));
    LocalMux I__1115 (
            .O(N__6671),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__1114 (
            .O(N__6668),
            .I(bfn_11_8_0_));
    InMux I__1113 (
            .O(N__6665),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__1112 (
            .O(N__6662),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__1111 (
            .O(N__6659),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__1110 (
            .O(N__6656),
            .I(N__6652));
    InMux I__1109 (
            .O(N__6655),
            .I(N__6644));
    LocalMux I__1108 (
            .O(N__6652),
            .I(N__6640));
    InMux I__1107 (
            .O(N__6651),
            .I(N__6635));
    InMux I__1106 (
            .O(N__6650),
            .I(N__6635));
    InMux I__1105 (
            .O(N__6649),
            .I(N__6632));
    CascadeMux I__1104 (
            .O(N__6648),
            .I(N__6629));
    InMux I__1103 (
            .O(N__6647),
            .I(N__6626));
    LocalMux I__1102 (
            .O(N__6644),
            .I(N__6623));
    InMux I__1101 (
            .O(N__6643),
            .I(N__6620));
    Span4Mux_v I__1100 (
            .O(N__6640),
            .I(N__6612));
    LocalMux I__1099 (
            .O(N__6635),
            .I(N__6612));
    LocalMux I__1098 (
            .O(N__6632),
            .I(N__6612));
    InMux I__1097 (
            .O(N__6629),
            .I(N__6609));
    LocalMux I__1096 (
            .O(N__6626),
            .I(N__6606));
    Span4Mux_v I__1095 (
            .O(N__6623),
            .I(N__6601));
    LocalMux I__1094 (
            .O(N__6620),
            .I(N__6601));
    InMux I__1093 (
            .O(N__6619),
            .I(N__6598));
    Span4Mux_h I__1092 (
            .O(N__6612),
            .I(N__6595));
    LocalMux I__1091 (
            .O(N__6609),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1090 (
            .O(N__6606),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1089 (
            .O(N__6601),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1088 (
            .O(N__6598),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1087 (
            .O(N__6595),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1086 (
            .O(N__6584),
            .I(N__6581));
    LocalMux I__1085 (
            .O(N__6581),
            .I(N__6578));
    Span4Mux_v I__1084 (
            .O(N__6578),
            .I(N__6573));
    InMux I__1083 (
            .O(N__6577),
            .I(N__6568));
    InMux I__1082 (
            .O(N__6576),
            .I(N__6568));
    Odrv4 I__1081 (
            .O(N__6573),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    LocalMux I__1080 (
            .O(N__6568),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    IoInMux I__1079 (
            .O(N__6563),
            .I(N__6560));
    LocalMux I__1078 (
            .O(N__6560),
            .I(N__6557));
    IoSpan4Mux I__1077 (
            .O(N__6557),
            .I(N__6554));
    IoSpan4Mux I__1076 (
            .O(N__6554),
            .I(N__6551));
    Span4Mux_s3_h I__1075 (
            .O(N__6551),
            .I(N__6547));
    InMux I__1074 (
            .O(N__6550),
            .I(N__6544));
    Span4Mux_h I__1073 (
            .O(N__6547),
            .I(N__6541));
    LocalMux I__1072 (
            .O(N__6544),
            .I(N__6538));
    Sp12to4 I__1071 (
            .O(N__6541),
            .I(N__6535));
    Span4Mux_v I__1070 (
            .O(N__6538),
            .I(N__6532));
    Span12Mux_h I__1069 (
            .O(N__6535),
            .I(N__6527));
    Sp12to4 I__1068 (
            .O(N__6532),
            .I(N__6527));
    Span12Mux_h I__1067 (
            .O(N__6527),
            .I(N__6524));
    Odrv12 I__1066 (
            .O(N__6524),
            .I(C3_c));
    InMux I__1065 (
            .O(N__6521),
            .I(N__6518));
    LocalMux I__1064 (
            .O(N__6518),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    CascadeMux I__1063 (
            .O(N__6515),
            .I(\U712_CHIP_RAM.N_28_0_cascade_ ));
    InMux I__1062 (
            .O(N__6512),
            .I(N__6509));
    LocalMux I__1061 (
            .O(N__6509),
            .I(\U712_CHIP_RAM.N_16_0 ));
    CascadeMux I__1060 (
            .O(N__6506),
            .I(\U712_CHIP_RAM.N_16_0_cascade_ ));
    CascadeMux I__1059 (
            .O(N__6503),
            .I(N__6489));
    InMux I__1058 (
            .O(N__6502),
            .I(N__6485));
    CascadeMux I__1057 (
            .O(N__6501),
            .I(N__6482));
    CascadeMux I__1056 (
            .O(N__6500),
            .I(N__6478));
    InMux I__1055 (
            .O(N__6499),
            .I(N__6471));
    InMux I__1054 (
            .O(N__6498),
            .I(N__6471));
    InMux I__1053 (
            .O(N__6497),
            .I(N__6471));
    InMux I__1052 (
            .O(N__6496),
            .I(N__6466));
    InMux I__1051 (
            .O(N__6495),
            .I(N__6463));
    InMux I__1050 (
            .O(N__6494),
            .I(N__6459));
    InMux I__1049 (
            .O(N__6493),
            .I(N__6450));
    InMux I__1048 (
            .O(N__6492),
            .I(N__6450));
    InMux I__1047 (
            .O(N__6489),
            .I(N__6450));
    InMux I__1046 (
            .O(N__6488),
            .I(N__6450));
    LocalMux I__1045 (
            .O(N__6485),
            .I(N__6439));
    InMux I__1044 (
            .O(N__6482),
            .I(N__6434));
    InMux I__1043 (
            .O(N__6481),
            .I(N__6434));
    InMux I__1042 (
            .O(N__6478),
            .I(N__6431));
    LocalMux I__1041 (
            .O(N__6471),
            .I(N__6428));
    InMux I__1040 (
            .O(N__6470),
            .I(N__6425));
    InMux I__1039 (
            .O(N__6469),
            .I(N__6422));
    LocalMux I__1038 (
            .O(N__6466),
            .I(N__6417));
    LocalMux I__1037 (
            .O(N__6463),
            .I(N__6417));
    InMux I__1036 (
            .O(N__6462),
            .I(N__6414));
    LocalMux I__1035 (
            .O(N__6459),
            .I(N__6409));
    LocalMux I__1034 (
            .O(N__6450),
            .I(N__6409));
    InMux I__1033 (
            .O(N__6449),
            .I(N__6404));
    InMux I__1032 (
            .O(N__6448),
            .I(N__6404));
    InMux I__1031 (
            .O(N__6447),
            .I(N__6397));
    InMux I__1030 (
            .O(N__6446),
            .I(N__6397));
    InMux I__1029 (
            .O(N__6445),
            .I(N__6397));
    InMux I__1028 (
            .O(N__6444),
            .I(N__6390));
    InMux I__1027 (
            .O(N__6443),
            .I(N__6390));
    InMux I__1026 (
            .O(N__6442),
            .I(N__6390));
    Span4Mux_v I__1025 (
            .O(N__6439),
            .I(N__6381));
    LocalMux I__1024 (
            .O(N__6434),
            .I(N__6381));
    LocalMux I__1023 (
            .O(N__6431),
            .I(N__6381));
    Span4Mux_v I__1022 (
            .O(N__6428),
            .I(N__6381));
    LocalMux I__1021 (
            .O(N__6425),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1020 (
            .O(N__6422),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1019 (
            .O(N__6417),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1018 (
            .O(N__6414),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1017 (
            .O(N__6409),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1016 (
            .O(N__6404),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1015 (
            .O(N__6397),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1014 (
            .O(N__6390),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1013 (
            .O(N__6381),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1012 (
            .O(N__6362),
            .I(N__6357));
    CascadeMux I__1011 (
            .O(N__6361),
            .I(N__6353));
    InMux I__1010 (
            .O(N__6360),
            .I(N__6350));
    LocalMux I__1009 (
            .O(N__6357),
            .I(N__6347));
    InMux I__1008 (
            .O(N__6356),
            .I(N__6344));
    InMux I__1007 (
            .O(N__6353),
            .I(N__6341));
    LocalMux I__1006 (
            .O(N__6350),
            .I(N__6338));
    Odrv4 I__1005 (
            .O(N__6347),
            .I(\U712_CHIP_RAM.N_111_0 ));
    LocalMux I__1004 (
            .O(N__6344),
            .I(\U712_CHIP_RAM.N_111_0 ));
    LocalMux I__1003 (
            .O(N__6341),
            .I(\U712_CHIP_RAM.N_111_0 ));
    Odrv12 I__1002 (
            .O(N__6338),
            .I(\U712_CHIP_RAM.N_111_0 ));
    InMux I__1001 (
            .O(N__6329),
            .I(N__6319));
    CascadeMux I__1000 (
            .O(N__6328),
            .I(N__6313));
    InMux I__999 (
            .O(N__6327),
            .I(N__6304));
    InMux I__998 (
            .O(N__6326),
            .I(N__6304));
    InMux I__997 (
            .O(N__6325),
            .I(N__6304));
    InMux I__996 (
            .O(N__6324),
            .I(N__6301));
    InMux I__995 (
            .O(N__6323),
            .I(N__6296));
    InMux I__994 (
            .O(N__6322),
            .I(N__6296));
    LocalMux I__993 (
            .O(N__6319),
            .I(N__6292));
    InMux I__992 (
            .O(N__6318),
            .I(N__6280));
    InMux I__991 (
            .O(N__6317),
            .I(N__6280));
    InMux I__990 (
            .O(N__6316),
            .I(N__6280));
    InMux I__989 (
            .O(N__6313),
            .I(N__6270));
    InMux I__988 (
            .O(N__6312),
            .I(N__6270));
    InMux I__987 (
            .O(N__6311),
            .I(N__6270));
    LocalMux I__986 (
            .O(N__6304),
            .I(N__6264));
    LocalMux I__985 (
            .O(N__6301),
            .I(N__6259));
    LocalMux I__984 (
            .O(N__6296),
            .I(N__6259));
    InMux I__983 (
            .O(N__6295),
            .I(N__6255));
    Span4Mux_h I__982 (
            .O(N__6292),
            .I(N__6252));
    InMux I__981 (
            .O(N__6291),
            .I(N__6247));
    InMux I__980 (
            .O(N__6290),
            .I(N__6247));
    InMux I__979 (
            .O(N__6289),
            .I(N__6240));
    InMux I__978 (
            .O(N__6288),
            .I(N__6240));
    InMux I__977 (
            .O(N__6287),
            .I(N__6240));
    LocalMux I__976 (
            .O(N__6280),
            .I(N__6237));
    InMux I__975 (
            .O(N__6279),
            .I(N__6230));
    InMux I__974 (
            .O(N__6278),
            .I(N__6230));
    InMux I__973 (
            .O(N__6277),
            .I(N__6230));
    LocalMux I__972 (
            .O(N__6270),
            .I(N__6227));
    InMux I__971 (
            .O(N__6269),
            .I(N__6220));
    InMux I__970 (
            .O(N__6268),
            .I(N__6220));
    InMux I__969 (
            .O(N__6267),
            .I(N__6220));
    Span4Mux_h I__968 (
            .O(N__6264),
            .I(N__6217));
    Span4Mux_h I__967 (
            .O(N__6259),
            .I(N__6214));
    InMux I__966 (
            .O(N__6258),
            .I(N__6211));
    LocalMux I__965 (
            .O(N__6255),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__964 (
            .O(N__6252),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__963 (
            .O(N__6247),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__962 (
            .O(N__6240),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__961 (
            .O(N__6237),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__960 (
            .O(N__6230),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__959 (
            .O(N__6227),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__958 (
            .O(N__6220),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__957 (
            .O(N__6217),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__956 (
            .O(N__6214),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__955 (
            .O(N__6211),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    CascadeMux I__954 (
            .O(N__6188),
            .I(\U712_CHIP_RAM.N_359_cascade_ ));
    InMux I__953 (
            .O(N__6185),
            .I(N__6182));
    LocalMux I__952 (
            .O(N__6182),
            .I(N__6177));
    InMux I__951 (
            .O(N__6181),
            .I(N__6173));
    InMux I__950 (
            .O(N__6180),
            .I(N__6170));
    Span4Mux_h I__949 (
            .O(N__6177),
            .I(N__6167));
    InMux I__948 (
            .O(N__6176),
            .I(N__6164));
    LocalMux I__947 (
            .O(N__6173),
            .I(\U712_CHIP_RAM.N_130_0 ));
    LocalMux I__946 (
            .O(N__6170),
            .I(\U712_CHIP_RAM.N_130_0 ));
    Odrv4 I__945 (
            .O(N__6167),
            .I(\U712_CHIP_RAM.N_130_0 ));
    LocalMux I__944 (
            .O(N__6164),
            .I(\U712_CHIP_RAM.N_130_0 ));
    CascadeMux I__943 (
            .O(N__6155),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_1_cascade_ ));
    InMux I__942 (
            .O(N__6152),
            .I(N__6149));
    LocalMux I__941 (
            .O(N__6149),
            .I(N__6146));
    Odrv4 I__940 (
            .O(N__6146),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1 ));
    CascadeMux I__939 (
            .O(N__6143),
            .I(\U712_CHIP_RAM.N_135_0_cascade_ ));
    InMux I__938 (
            .O(N__6140),
            .I(N__6137));
    LocalMux I__937 (
            .O(N__6137),
            .I(\U712_CHIP_RAM.N_125_0 ));
    CascadeMux I__936 (
            .O(N__6134),
            .I(N__6125));
    InMux I__935 (
            .O(N__6133),
            .I(N__6120));
    InMux I__934 (
            .O(N__6132),
            .I(N__6117));
    InMux I__933 (
            .O(N__6131),
            .I(N__6114));
    InMux I__932 (
            .O(N__6130),
            .I(N__6111));
    InMux I__931 (
            .O(N__6129),
            .I(N__6105));
    InMux I__930 (
            .O(N__6128),
            .I(N__6105));
    InMux I__929 (
            .O(N__6125),
            .I(N__6102));
    InMux I__928 (
            .O(N__6124),
            .I(N__6098));
    InMux I__927 (
            .O(N__6123),
            .I(N__6093));
    LocalMux I__926 (
            .O(N__6120),
            .I(N__6086));
    LocalMux I__925 (
            .O(N__6117),
            .I(N__6086));
    LocalMux I__924 (
            .O(N__6114),
            .I(N__6086));
    LocalMux I__923 (
            .O(N__6111),
            .I(N__6083));
    InMux I__922 (
            .O(N__6110),
            .I(N__6077));
    LocalMux I__921 (
            .O(N__6105),
            .I(N__6073));
    LocalMux I__920 (
            .O(N__6102),
            .I(N__6070));
    InMux I__919 (
            .O(N__6101),
            .I(N__6067));
    LocalMux I__918 (
            .O(N__6098),
            .I(N__6064));
    InMux I__917 (
            .O(N__6097),
            .I(N__6059));
    InMux I__916 (
            .O(N__6096),
            .I(N__6059));
    LocalMux I__915 (
            .O(N__6093),
            .I(N__6052));
    Span4Mux_v I__914 (
            .O(N__6086),
            .I(N__6052));
    Span4Mux_v I__913 (
            .O(N__6083),
            .I(N__6052));
    InMux I__912 (
            .O(N__6082),
            .I(N__6045));
    InMux I__911 (
            .O(N__6081),
            .I(N__6045));
    InMux I__910 (
            .O(N__6080),
            .I(N__6045));
    LocalMux I__909 (
            .O(N__6077),
            .I(N__6042));
    InMux I__908 (
            .O(N__6076),
            .I(N__6039));
    Odrv4 I__907 (
            .O(N__6073),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__906 (
            .O(N__6070),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__905 (
            .O(N__6067),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__904 (
            .O(N__6064),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__903 (
            .O(N__6059),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__902 (
            .O(N__6052),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__901 (
            .O(N__6045),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__900 (
            .O(N__6042),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__899 (
            .O(N__6039),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__898 (
            .O(N__6020),
            .I(N__6017));
    LocalMux I__897 (
            .O(N__6017),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_3 ));
    InMux I__896 (
            .O(N__6014),
            .I(N__6011));
    LocalMux I__895 (
            .O(N__6011),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_3 ));
    InMux I__894 (
            .O(N__6008),
            .I(N__6002));
    InMux I__893 (
            .O(N__6007),
            .I(N__5999));
    InMux I__892 (
            .O(N__6006),
            .I(N__5996));
    InMux I__891 (
            .O(N__6005),
            .I(N__5993));
    LocalMux I__890 (
            .O(N__6002),
            .I(N__5990));
    LocalMux I__889 (
            .O(N__5999),
            .I(\U712_CHIP_RAM.N_204_0 ));
    LocalMux I__888 (
            .O(N__5996),
            .I(\U712_CHIP_RAM.N_204_0 ));
    LocalMux I__887 (
            .O(N__5993),
            .I(\U712_CHIP_RAM.N_204_0 ));
    Odrv4 I__886 (
            .O(N__5990),
            .I(\U712_CHIP_RAM.N_204_0 ));
    CascadeMux I__885 (
            .O(N__5981),
            .I(\U712_CHIP_RAM.N_120_0_cascade_ ));
    InMux I__884 (
            .O(N__5978),
            .I(N__5975));
    LocalMux I__883 (
            .O(N__5975),
            .I(\U712_CHIP_RAM.N_363 ));
    InMux I__882 (
            .O(N__5972),
            .I(N__5969));
    LocalMux I__881 (
            .O(N__5969),
            .I(\U712_CHIP_RAM.m225_0 ));
    CascadeMux I__880 (
            .O(N__5966),
            .I(N__5962));
    CascadeMux I__879 (
            .O(N__5965),
            .I(N__5959));
    InMux I__878 (
            .O(N__5962),
            .I(N__5949));
    InMux I__877 (
            .O(N__5959),
            .I(N__5949));
    CascadeMux I__876 (
            .O(N__5958),
            .I(N__5944));
    CascadeMux I__875 (
            .O(N__5957),
            .I(N__5941));
    InMux I__874 (
            .O(N__5956),
            .I(N__5936));
    InMux I__873 (
            .O(N__5955),
            .I(N__5931));
    InMux I__872 (
            .O(N__5954),
            .I(N__5931));
    LocalMux I__871 (
            .O(N__5949),
            .I(N__5928));
    InMux I__870 (
            .O(N__5948),
            .I(N__5925));
    InMux I__869 (
            .O(N__5947),
            .I(N__5920));
    InMux I__868 (
            .O(N__5944),
            .I(N__5917));
    InMux I__867 (
            .O(N__5941),
            .I(N__5910));
    InMux I__866 (
            .O(N__5940),
            .I(N__5910));
    InMux I__865 (
            .O(N__5939),
            .I(N__5910));
    LocalMux I__864 (
            .O(N__5936),
            .I(N__5905));
    LocalMux I__863 (
            .O(N__5931),
            .I(N__5905));
    Span4Mux_v I__862 (
            .O(N__5928),
            .I(N__5900));
    LocalMux I__861 (
            .O(N__5925),
            .I(N__5900));
    InMux I__860 (
            .O(N__5924),
            .I(N__5895));
    InMux I__859 (
            .O(N__5923),
            .I(N__5895));
    LocalMux I__858 (
            .O(N__5920),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__857 (
            .O(N__5917),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__856 (
            .O(N__5910),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__855 (
            .O(N__5905),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__854 (
            .O(N__5900),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__853 (
            .O(N__5895),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__852 (
            .O(N__5882),
            .I(N__5876));
    CascadeMux I__851 (
            .O(N__5881),
            .I(N__5870));
    InMux I__850 (
            .O(N__5880),
            .I(N__5864));
    InMux I__849 (
            .O(N__5879),
            .I(N__5864));
    InMux I__848 (
            .O(N__5876),
            .I(N__5858));
    InMux I__847 (
            .O(N__5875),
            .I(N__5858));
    InMux I__846 (
            .O(N__5874),
            .I(N__5852));
    InMux I__845 (
            .O(N__5873),
            .I(N__5852));
    InMux I__844 (
            .O(N__5870),
            .I(N__5849));
    InMux I__843 (
            .O(N__5869),
            .I(N__5846));
    LocalMux I__842 (
            .O(N__5864),
            .I(N__5843));
    InMux I__841 (
            .O(N__5863),
            .I(N__5840));
    LocalMux I__840 (
            .O(N__5858),
            .I(N__5837));
    InMux I__839 (
            .O(N__5857),
            .I(N__5834));
    LocalMux I__838 (
            .O(N__5852),
            .I(\U712_CHIP_RAM.N_110_0 ));
    LocalMux I__837 (
            .O(N__5849),
            .I(\U712_CHIP_RAM.N_110_0 ));
    LocalMux I__836 (
            .O(N__5846),
            .I(\U712_CHIP_RAM.N_110_0 ));
    Odrv4 I__835 (
            .O(N__5843),
            .I(\U712_CHIP_RAM.N_110_0 ));
    LocalMux I__834 (
            .O(N__5840),
            .I(\U712_CHIP_RAM.N_110_0 ));
    Odrv4 I__833 (
            .O(N__5837),
            .I(\U712_CHIP_RAM.N_110_0 ));
    LocalMux I__832 (
            .O(N__5834),
            .I(\U712_CHIP_RAM.N_110_0 ));
    InMux I__831 (
            .O(N__5819),
            .I(N__5816));
    LocalMux I__830 (
            .O(N__5816),
            .I(\U712_CHIP_RAM.N_112_0 ));
    CascadeMux I__829 (
            .O(N__5813),
            .I(\U712_CHIP_RAM.N_112_0_cascade_ ));
    CascadeMux I__828 (
            .O(N__5810),
            .I(N__5806));
    InMux I__827 (
            .O(N__5809),
            .I(N__5802));
    InMux I__826 (
            .O(N__5806),
            .I(N__5793));
    InMux I__825 (
            .O(N__5805),
            .I(N__5790));
    LocalMux I__824 (
            .O(N__5802),
            .I(N__5787));
    InMux I__823 (
            .O(N__5801),
            .I(N__5780));
    InMux I__822 (
            .O(N__5800),
            .I(N__5780));
    InMux I__821 (
            .O(N__5799),
            .I(N__5780));
    InMux I__820 (
            .O(N__5798),
            .I(N__5775));
    InMux I__819 (
            .O(N__5797),
            .I(N__5775));
    InMux I__818 (
            .O(N__5796),
            .I(N__5772));
    LocalMux I__817 (
            .O(N__5793),
            .I(\U712_CHIP_RAM.N_94_0 ));
    LocalMux I__816 (
            .O(N__5790),
            .I(\U712_CHIP_RAM.N_94_0 ));
    Odrv4 I__815 (
            .O(N__5787),
            .I(\U712_CHIP_RAM.N_94_0 ));
    LocalMux I__814 (
            .O(N__5780),
            .I(\U712_CHIP_RAM.N_94_0 ));
    LocalMux I__813 (
            .O(N__5775),
            .I(\U712_CHIP_RAM.N_94_0 ));
    LocalMux I__812 (
            .O(N__5772),
            .I(\U712_CHIP_RAM.N_94_0 ));
    CascadeMux I__811 (
            .O(N__5759),
            .I(N__5756));
    InMux I__810 (
            .O(N__5756),
            .I(N__5753));
    LocalMux I__809 (
            .O(N__5753),
            .I(N__5749));
    IoInMux I__808 (
            .O(N__5752),
            .I(N__5746));
    Span12Mux_h I__807 (
            .O(N__5749),
            .I(N__5743));
    LocalMux I__806 (
            .O(N__5746),
            .I(N__5740));
    Span12Mux_v I__805 (
            .O(N__5743),
            .I(N__5737));
    IoSpan4Mux I__804 (
            .O(N__5740),
            .I(N__5734));
    Odrv12 I__803 (
            .O(N__5737),
            .I(RAMENn_c));
    Odrv4 I__802 (
            .O(N__5734),
            .I(RAMENn_c));
    InMux I__801 (
            .O(N__5729),
            .I(N__5723));
    InMux I__800 (
            .O(N__5728),
            .I(N__5720));
    InMux I__799 (
            .O(N__5727),
            .I(N__5715));
    InMux I__798 (
            .O(N__5726),
            .I(N__5715));
    LocalMux I__797 (
            .O(N__5723),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__796 (
            .O(N__5720),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__795 (
            .O(N__5715),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__794 (
            .O(N__5708),
            .I(N__5705));
    LocalMux I__793 (
            .O(N__5705),
            .I(N__5702));
    Span4Mux_v I__792 (
            .O(N__5702),
            .I(N__5699));
    Sp12to4 I__791 (
            .O(N__5699),
            .I(N__5696));
    Span12Mux_h I__790 (
            .O(N__5696),
            .I(N__5693));
    Span12Mux_v I__789 (
            .O(N__5693),
            .I(N__5690));
    Odrv12 I__788 (
            .O(N__5690),
            .I(REGSPACEn_c));
    InMux I__787 (
            .O(N__5687),
            .I(N__5684));
    LocalMux I__786 (
            .O(N__5684),
            .I(N__5680));
    InMux I__785 (
            .O(N__5683),
            .I(N__5677));
    Span4Mux_h I__784 (
            .O(N__5680),
            .I(N__5672));
    LocalMux I__783 (
            .O(N__5677),
            .I(N__5672));
    Span4Mux_v I__782 (
            .O(N__5672),
            .I(N__5669));
    Span4Mux_v I__781 (
            .O(N__5669),
            .I(N__5666));
    Sp12to4 I__780 (
            .O(N__5666),
            .I(N__5663));
    Span12Mux_h I__779 (
            .O(N__5663),
            .I(N__5660));
    Odrv12 I__778 (
            .O(N__5660),
            .I(TSn_c));
    CascadeMux I__777 (
            .O(N__5657),
            .I(N__5654));
    InMux I__776 (
            .O(N__5654),
            .I(N__5648));
    InMux I__775 (
            .O(N__5653),
            .I(N__5648));
    LocalMux I__774 (
            .O(N__5648),
            .I(U712_REG_SM_START_RST));
    InMux I__773 (
            .O(N__5645),
            .I(N__5636));
    InMux I__772 (
            .O(N__5644),
            .I(N__5636));
    InMux I__771 (
            .O(N__5643),
            .I(N__5636));
    LocalMux I__770 (
            .O(N__5636),
            .I(N__5629));
    InMux I__769 (
            .O(N__5635),
            .I(N__5626));
    InMux I__768 (
            .O(N__5634),
            .I(N__5623));
    InMux I__767 (
            .O(N__5633),
            .I(N__5620));
    InMux I__766 (
            .O(N__5632),
            .I(N__5617));
    Odrv4 I__765 (
            .O(N__5629),
            .I(\U712_CHIP_RAM.N_96_0 ));
    LocalMux I__764 (
            .O(N__5626),
            .I(\U712_CHIP_RAM.N_96_0 ));
    LocalMux I__763 (
            .O(N__5623),
            .I(\U712_CHIP_RAM.N_96_0 ));
    LocalMux I__762 (
            .O(N__5620),
            .I(\U712_CHIP_RAM.N_96_0 ));
    LocalMux I__761 (
            .O(N__5617),
            .I(\U712_CHIP_RAM.N_96_0 ));
    CascadeMux I__760 (
            .O(N__5606),
            .I(\U712_CHIP_RAM.m123_0_cascade_ ));
    InMux I__759 (
            .O(N__5603),
            .I(N__5600));
    LocalMux I__758 (
            .O(N__5600),
            .I(\U712_CHIP_RAM.N_117_0 ));
    InMux I__757 (
            .O(N__5597),
            .I(N__5593));
    InMux I__756 (
            .O(N__5596),
            .I(N__5587));
    LocalMux I__755 (
            .O(N__5593),
            .I(N__5584));
    InMux I__754 (
            .O(N__5592),
            .I(N__5577));
    InMux I__753 (
            .O(N__5591),
            .I(N__5577));
    InMux I__752 (
            .O(N__5590),
            .I(N__5577));
    LocalMux I__751 (
            .O(N__5587),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    Odrv12 I__750 (
            .O(N__5584),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__749 (
            .O(N__5577),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__748 (
            .O(N__5570),
            .I(N__5566));
    InMux I__747 (
            .O(N__5569),
            .I(N__5563));
    InMux I__746 (
            .O(N__5566),
            .I(N__5560));
    LocalMux I__745 (
            .O(N__5563),
            .I(N__5552));
    LocalMux I__744 (
            .O(N__5560),
            .I(N__5552));
    InMux I__743 (
            .O(N__5559),
            .I(N__5545));
    InMux I__742 (
            .O(N__5558),
            .I(N__5545));
    InMux I__741 (
            .O(N__5557),
            .I(N__5545));
    Odrv4 I__740 (
            .O(N__5552),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__739 (
            .O(N__5545),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    CascadeMux I__738 (
            .O(N__5540),
            .I(N__5536));
    InMux I__737 (
            .O(N__5539),
            .I(N__5530));
    InMux I__736 (
            .O(N__5536),
            .I(N__5530));
    InMux I__735 (
            .O(N__5535),
            .I(N__5527));
    LocalMux I__734 (
            .O(N__5530),
            .I(N__5524));
    LocalMux I__733 (
            .O(N__5527),
            .I(\U712_CHIP_RAM.m92_0 ));
    Odrv4 I__732 (
            .O(N__5524),
            .I(\U712_CHIP_RAM.m92_0 ));
    CascadeMux I__731 (
            .O(N__5519),
            .I(\U712_CHIP_RAM.N_130_0_cascade_ ));
    CascadeMux I__730 (
            .O(N__5516),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5Z0Z_3_cascade_ ));
    InMux I__729 (
            .O(N__5513),
            .I(N__5510));
    LocalMux I__728 (
            .O(N__5510),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIG3845Z0Z_0 ));
    InMux I__727 (
            .O(N__5507),
            .I(N__5504));
    LocalMux I__726 (
            .O(N__5504),
            .I(\U712_CHIP_RAM.m203_ns_1 ));
    CascadeMux I__725 (
            .O(N__5501),
            .I(\U712_CHIP_RAM.N_363_mux_cascade_ ));
    CascadeMux I__724 (
            .O(N__5498),
            .I(N__5495));
    InMux I__723 (
            .O(N__5495),
            .I(N__5492));
    LocalMux I__722 (
            .O(N__5492),
            .I(N__5489));
    Span4Mux_v I__721 (
            .O(N__5489),
            .I(N__5485));
    InMux I__720 (
            .O(N__5488),
            .I(N__5482));
    Odrv4 I__719 (
            .O(N__5485),
            .I(\U712_CHIP_RAM.m186_0 ));
    LocalMux I__718 (
            .O(N__5482),
            .I(\U712_CHIP_RAM.m186_0 ));
    InMux I__717 (
            .O(N__5477),
            .I(N__5474));
    LocalMux I__716 (
            .O(N__5474),
            .I(\U712_CHIP_RAM.m141_ns_1 ));
    InMux I__715 (
            .O(N__5471),
            .I(N__5465));
    InMux I__714 (
            .O(N__5470),
            .I(N__5465));
    LocalMux I__713 (
            .O(N__5465),
            .I(\U712_CHIP_RAM.N_140_0 ));
    CascadeMux I__712 (
            .O(N__5462),
            .I(\U712_CHIP_RAM.N_140_0_cascade_ ));
    InMux I__711 (
            .O(N__5459),
            .I(N__5454));
    InMux I__710 (
            .O(N__5458),
            .I(N__5451));
    InMux I__709 (
            .O(N__5457),
            .I(N__5446));
    LocalMux I__708 (
            .O(N__5454),
            .I(N__5443));
    LocalMux I__707 (
            .O(N__5451),
            .I(N__5440));
    InMux I__706 (
            .O(N__5450),
            .I(N__5435));
    InMux I__705 (
            .O(N__5449),
            .I(N__5435));
    LocalMux I__704 (
            .O(N__5446),
            .I(\U712_CHIP_RAM.N_103_0 ));
    Odrv4 I__703 (
            .O(N__5443),
            .I(\U712_CHIP_RAM.N_103_0 ));
    Odrv4 I__702 (
            .O(N__5440),
            .I(\U712_CHIP_RAM.N_103_0 ));
    LocalMux I__701 (
            .O(N__5435),
            .I(\U712_CHIP_RAM.N_103_0 ));
    InMux I__700 (
            .O(N__5426),
            .I(N__5422));
    InMux I__699 (
            .O(N__5425),
            .I(N__5419));
    LocalMux I__698 (
            .O(N__5422),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ));
    LocalMux I__697 (
            .O(N__5419),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ));
    InMux I__696 (
            .O(N__5414),
            .I(N__5410));
    InMux I__695 (
            .O(N__5413),
            .I(N__5407));
    LocalMux I__694 (
            .O(N__5410),
            .I(N__5404));
    LocalMux I__693 (
            .O(N__5407),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    Odrv4 I__692 (
            .O(N__5404),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    InMux I__691 (
            .O(N__5399),
            .I(N__5395));
    InMux I__690 (
            .O(N__5398),
            .I(N__5392));
    LocalMux I__689 (
            .O(N__5395),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ));
    LocalMux I__688 (
            .O(N__5392),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ));
    InMux I__687 (
            .O(N__5387),
            .I(N__5383));
    InMux I__686 (
            .O(N__5386),
            .I(N__5380));
    LocalMux I__685 (
            .O(N__5383),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ));
    LocalMux I__684 (
            .O(N__5380),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ));
    InMux I__683 (
            .O(N__5375),
            .I(N__5367));
    InMux I__682 (
            .O(N__5374),
            .I(N__5367));
    InMux I__681 (
            .O(N__5373),
            .I(N__5364));
    InMux I__680 (
            .O(N__5372),
            .I(N__5361));
    LocalMux I__679 (
            .O(N__5367),
            .I(N__5358));
    LocalMux I__678 (
            .O(N__5364),
            .I(N__5355));
    LocalMux I__677 (
            .O(N__5361),
            .I(N__5352));
    Span4Mux_h I__676 (
            .O(N__5358),
            .I(N__5349));
    Odrv4 I__675 (
            .O(N__5355),
            .I(\U712_CHIP_RAM.N_358 ));
    Odrv4 I__674 (
            .O(N__5352),
            .I(\U712_CHIP_RAM.N_358 ));
    Odrv4 I__673 (
            .O(N__5349),
            .I(\U712_CHIP_RAM.N_358 ));
    InMux I__672 (
            .O(N__5342),
            .I(N__5337));
    InMux I__671 (
            .O(N__5341),
            .I(N__5334));
    InMux I__670 (
            .O(N__5340),
            .I(N__5331));
    LocalMux I__669 (
            .O(N__5337),
            .I(\U712_CHIP_RAM.N_188_0 ));
    LocalMux I__668 (
            .O(N__5334),
            .I(\U712_CHIP_RAM.N_188_0 ));
    LocalMux I__667 (
            .O(N__5331),
            .I(\U712_CHIP_RAM.N_188_0 ));
    CEMux I__666 (
            .O(N__5324),
            .I(N__5321));
    LocalMux I__665 (
            .O(N__5321),
            .I(N__5318));
    Span4Mux_v I__664 (
            .O(N__5318),
            .I(N__5315));
    Odrv4 I__663 (
            .O(N__5315),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0 ));
    InMux I__662 (
            .O(N__5312),
            .I(N__5309));
    LocalMux I__661 (
            .O(N__5309),
            .I(N__5305));
    InMux I__660 (
            .O(N__5308),
            .I(N__5302));
    Odrv4 I__659 (
            .O(N__5305),
            .I(\U712_CHIP_RAM.N_344 ));
    LocalMux I__658 (
            .O(N__5302),
            .I(\U712_CHIP_RAM.N_344 ));
    CascadeMux I__657 (
            .O(N__5297),
            .I(\U712_CHIP_RAM.N_358_cascade_ ));
    InMux I__656 (
            .O(N__5294),
            .I(N__5291));
    LocalMux I__655 (
            .O(N__5291),
            .I(\U712_CHIP_RAM.m219_0 ));
    CascadeMux I__654 (
            .O(N__5288),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_2_cascade_ ));
    InMux I__653 (
            .O(N__5285),
            .I(N__5282));
    LocalMux I__652 (
            .O(N__5282),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2 ));
    CascadeMux I__651 (
            .O(N__5279),
            .I(N__5276));
    InMux I__650 (
            .O(N__5276),
            .I(N__5273));
    LocalMux I__649 (
            .O(N__5273),
            .I(N__5269));
    InMux I__648 (
            .O(N__5272),
            .I(N__5266));
    Odrv4 I__647 (
            .O(N__5269),
            .I(\U712_CHIP_RAM.N_137_0 ));
    LocalMux I__646 (
            .O(N__5266),
            .I(\U712_CHIP_RAM.N_137_0 ));
    CascadeMux I__645 (
            .O(N__5261),
            .I(\U712_CHIP_RAM.N_142_0_cascade_ ));
    IoInMux I__644 (
            .O(N__5258),
            .I(N__5255));
    LocalMux I__643 (
            .O(N__5255),
            .I(N__5252));
    Span4Mux_s1_h I__642 (
            .O(N__5252),
            .I(N__5249));
    Sp12to4 I__641 (
            .O(N__5249),
            .I(N__5246));
    Span12Mux_v I__640 (
            .O(N__5246),
            .I(N__5243));
    Span12Mux_h I__639 (
            .O(N__5243),
            .I(N__5239));
    InMux I__638 (
            .O(N__5242),
            .I(N__5236));
    Odrv12 I__637 (
            .O(N__5239),
            .I(CLK_EN_c));
    LocalMux I__636 (
            .O(N__5236),
            .I(CLK_EN_c));
    InMux I__635 (
            .O(N__5231),
            .I(N__5228));
    LocalMux I__634 (
            .O(N__5228),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER43 ));
    CascadeMux I__633 (
            .O(N__5225),
            .I(\U712_CHIP_RAM.m207_ns_1_cascade_ ));
    InMux I__632 (
            .O(N__5222),
            .I(N__5219));
    LocalMux I__631 (
            .O(N__5219),
            .I(\U712_CHIP_RAM.N_206_0 ));
    CascadeMux I__630 (
            .O(N__5216),
            .I(N__5213));
    InMux I__629 (
            .O(N__5213),
            .I(N__5210));
    LocalMux I__628 (
            .O(N__5210),
            .I(N__5207));
    Span4Mux_v I__627 (
            .O(N__5207),
            .I(N__5204));
    Odrv4 I__626 (
            .O(N__5204),
            .I(\U712_CHIP_RAM.N_208_0 ));
    InMux I__625 (
            .O(N__5201),
            .I(N__5197));
    InMux I__624 (
            .O(N__5200),
            .I(N__5194));
    LocalMux I__623 (
            .O(N__5197),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__622 (
            .O(N__5194),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__621 (
            .O(N__5189),
            .I(N__5185));
    InMux I__620 (
            .O(N__5188),
            .I(N__5182));
    LocalMux I__619 (
            .O(N__5185),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__618 (
            .O(N__5182),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__617 (
            .O(N__5177),
            .I(\U712_CHIP_RAM.m92_0_cascade_ ));
    InMux I__616 (
            .O(N__5174),
            .I(N__5171));
    LocalMux I__615 (
            .O(N__5171),
            .I(\U712_CHIP_RAM.N_190_0 ));
    CascadeMux I__614 (
            .O(N__5168),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_ ));
    CascadeMux I__613 (
            .O(N__5165),
            .I(N__5161));
    InMux I__612 (
            .O(N__5164),
            .I(N__5157));
    InMux I__611 (
            .O(N__5161),
            .I(N__5152));
    InMux I__610 (
            .O(N__5160),
            .I(N__5152));
    LocalMux I__609 (
            .O(N__5157),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__608 (
            .O(N__5152),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    CascadeMux I__607 (
            .O(N__5147),
            .I(\U712_CHIP_RAM.N_222_0_cascade_ ));
    CEMux I__606 (
            .O(N__5144),
            .I(N__5141));
    LocalMux I__605 (
            .O(N__5141),
            .I(N__5138));
    Span4Mux_v I__604 (
            .O(N__5138),
            .I(N__5134));
    CEMux I__603 (
            .O(N__5137),
            .I(N__5131));
    Span4Mux_v I__602 (
            .O(N__5134),
            .I(N__5126));
    LocalMux I__601 (
            .O(N__5131),
            .I(N__5126));
    Odrv4 I__600 (
            .O(N__5126),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__599 (
            .O(N__5123),
            .I(N__5119));
    InMux I__598 (
            .O(N__5122),
            .I(N__5116));
    LocalMux I__597 (
            .O(N__5119),
            .I(N__5111));
    LocalMux I__596 (
            .O(N__5116),
            .I(N__5108));
    InMux I__595 (
            .O(N__5115),
            .I(N__5102));
    InMux I__594 (
            .O(N__5114),
            .I(N__5102));
    Span4Mux_h I__593 (
            .O(N__5111),
            .I(N__5099));
    Span4Mux_h I__592 (
            .O(N__5108),
            .I(N__5096));
    InMux I__591 (
            .O(N__5107),
            .I(N__5093));
    LocalMux I__590 (
            .O(N__5102),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__589 (
            .O(N__5099),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__588 (
            .O(N__5096),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__587 (
            .O(N__5093),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    CascadeMux I__586 (
            .O(N__5084),
            .I(\U712_CHIP_RAM.N_111_0_cascade_ ));
    InMux I__585 (
            .O(N__5081),
            .I(N__5078));
    LocalMux I__584 (
            .O(N__5078),
            .I(\U712_CHIP_RAM.N_50 ));
    InMux I__583 (
            .O(N__5075),
            .I(N__5072));
    LocalMux I__582 (
            .O(N__5072),
            .I(N__5069));
    Odrv4 I__581 (
            .O(N__5069),
            .I(\U712_CHIP_RAM.m138_0 ));
    CascadeMux I__580 (
            .O(N__5066),
            .I(\U712_CHIP_RAM.N_352_mux_cascade_ ));
    InMux I__579 (
            .O(N__5063),
            .I(N__5060));
    LocalMux I__578 (
            .O(N__5060),
            .I(\U712_CHIP_RAM.N_183_0 ));
    CascadeMux I__577 (
            .O(N__5057),
            .I(\U712_CHIP_RAM.N_137_0_cascade_ ));
    InMux I__576 (
            .O(N__5054),
            .I(N__5051));
    LocalMux I__575 (
            .O(N__5051),
            .I(\U712_CHIP_RAM.N_178_0 ));
    CascadeMux I__574 (
            .O(N__5048),
            .I(\U712_CHIP_RAM.N_94_0_cascade_ ));
    CascadeMux I__573 (
            .O(N__5045),
            .I(\U712_CHIP_RAM.N_96_0_cascade_ ));
    IoInMux I__572 (
            .O(N__5042),
            .I(N__5039));
    LocalMux I__571 (
            .O(N__5039),
            .I(N__5036));
    Span12Mux_s7_v I__570 (
            .O(N__5036),
            .I(N__5033));
    Odrv12 I__569 (
            .O(N__5033),
            .I(VBENn_c));
    InMux I__568 (
            .O(N__5030),
            .I(N__5027));
    LocalMux I__567 (
            .O(N__5027),
            .I(N__5024));
    Span12Mux_h I__566 (
            .O(N__5024),
            .I(N__5021));
    Span12Mux_v I__565 (
            .O(N__5021),
            .I(N__5018));
    Odrv12 I__564 (
            .O(N__5018),
            .I(A_c_2));
    InMux I__563 (
            .O(N__5015),
            .I(N__5012));
    LocalMux I__562 (
            .O(N__5012),
            .I(N__5009));
    Span4Mux_v I__561 (
            .O(N__5009),
            .I(N__5006));
    Span4Mux_v I__560 (
            .O(N__5006),
            .I(N__5003));
    Sp12to4 I__559 (
            .O(N__5003),
            .I(N__5000));
    Odrv12 I__558 (
            .O(N__5000),
            .I(A_c_5));
    InMux I__557 (
            .O(N__4997),
            .I(N__4994));
    LocalMux I__556 (
            .O(N__4994),
            .I(N__4991));
    Span4Mux_v I__555 (
            .O(N__4991),
            .I(N__4988));
    Span4Mux_h I__554 (
            .O(N__4988),
            .I(N__4985));
    Span4Mux_h I__553 (
            .O(N__4985),
            .I(N__4982));
    Odrv4 I__552 (
            .O(N__4982),
            .I(A_c_6));
    InMux I__551 (
            .O(N__4979),
            .I(N__4976));
    LocalMux I__550 (
            .O(N__4976),
            .I(N__4973));
    Span4Mux_h I__549 (
            .O(N__4973),
            .I(N__4970));
    Sp12to4 I__548 (
            .O(N__4970),
            .I(N__4967));
    Span12Mux_v I__547 (
            .O(N__4967),
            .I(N__4964));
    Odrv12 I__546 (
            .O(N__4964),
            .I(A_c_3));
    InMux I__545 (
            .O(N__4961),
            .I(N__4958));
    LocalMux I__544 (
            .O(N__4958),
            .I(N__4955));
    Span12Mux_v I__543 (
            .O(N__4955),
            .I(N__4952));
    Odrv12 I__542 (
            .O(N__4952),
            .I(A_c_7));
    InMux I__541 (
            .O(N__4949),
            .I(N__4946));
    LocalMux I__540 (
            .O(N__4946),
            .I(N__4943));
    Span4Mux_v I__539 (
            .O(N__4943),
            .I(N__4940));
    Span4Mux_v I__538 (
            .O(N__4940),
            .I(N__4937));
    Span4Mux_h I__537 (
            .O(N__4937),
            .I(N__4934));
    Span4Mux_h I__536 (
            .O(N__4934),
            .I(N__4931));
    Odrv4 I__535 (
            .O(N__4931),
            .I(A_c_4));
    InMux I__534 (
            .O(N__4928),
            .I(N__4907));
    InMux I__533 (
            .O(N__4927),
            .I(N__4907));
    InMux I__532 (
            .O(N__4926),
            .I(N__4907));
    InMux I__531 (
            .O(N__4925),
            .I(N__4907));
    InMux I__530 (
            .O(N__4924),
            .I(N__4907));
    InMux I__529 (
            .O(N__4923),
            .I(N__4907));
    InMux I__528 (
            .O(N__4922),
            .I(N__4902));
    InMux I__527 (
            .O(N__4921),
            .I(N__4902));
    InMux I__526 (
            .O(N__4920),
            .I(N__4899));
    LocalMux I__525 (
            .O(N__4907),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    LocalMux I__524 (
            .O(N__4902),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    LocalMux I__523 (
            .O(N__4899),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    CascadeMux I__522 (
            .O(N__4892),
            .I(\U712_CHIP_RAM.N_206_0_cascade_ ));
    CascadeMux I__521 (
            .O(N__4889),
            .I(\U712_CHIP_RAM.N_214_0_cascade_ ));
    InMux I__520 (
            .O(N__4886),
            .I(N__4883));
    LocalMux I__519 (
            .O(N__4883),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    CascadeMux I__518 (
            .O(N__4880),
            .I(\U712_CHIP_RAM.N_216_0_i_cascade_ ));
    CascadeMux I__517 (
            .O(N__4877),
            .I(N__4873));
    InMux I__516 (
            .O(N__4876),
            .I(N__4870));
    InMux I__515 (
            .O(N__4873),
            .I(N__4867));
    LocalMux I__514 (
            .O(N__4870),
            .I(N__4864));
    LocalMux I__513 (
            .O(N__4867),
            .I(\U712_CHIP_RAM.N_217_0 ));
    Odrv12 I__512 (
            .O(N__4864),
            .I(\U712_CHIP_RAM.N_217_0 ));
    InMux I__511 (
            .O(N__4859),
            .I(N__4850));
    InMux I__510 (
            .O(N__4858),
            .I(N__4841));
    InMux I__509 (
            .O(N__4857),
            .I(N__4841));
    InMux I__508 (
            .O(N__4856),
            .I(N__4841));
    InMux I__507 (
            .O(N__4855),
            .I(N__4841));
    InMux I__506 (
            .O(N__4854),
            .I(N__4836));
    InMux I__505 (
            .O(N__4853),
            .I(N__4836));
    LocalMux I__504 (
            .O(N__4850),
            .I(\U712_CHIP_RAM.N_216_0_i ));
    LocalMux I__503 (
            .O(N__4841),
            .I(\U712_CHIP_RAM.N_216_0_i ));
    LocalMux I__502 (
            .O(N__4836),
            .I(\U712_CHIP_RAM.N_216_0_i ));
    InMux I__501 (
            .O(N__4829),
            .I(N__4826));
    LocalMux I__500 (
            .O(N__4826),
            .I(N__4823));
    Odrv4 I__499 (
            .O(N__4823),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    CascadeMux I__498 (
            .O(N__4820),
            .I(\U712_CHIP_RAM.N_195_0_cascade_ ));
    InMux I__497 (
            .O(N__4817),
            .I(N__4814));
    LocalMux I__496 (
            .O(N__4814),
            .I(\U712_CHIP_RAM.N_213_0 ));
    CascadeMux I__495 (
            .O(N__4811),
            .I(N__4808));
    InMux I__494 (
            .O(N__4808),
            .I(N__4805));
    LocalMux I__493 (
            .O(N__4805),
            .I(N__4801));
    InMux I__492 (
            .O(N__4804),
            .I(N__4798));
    Odrv4 I__491 (
            .O(N__4801),
            .I(\U712_CHIP_RAM.N_189_0 ));
    LocalMux I__490 (
            .O(N__4798),
            .I(\U712_CHIP_RAM.N_189_0 ));
    InMux I__489 (
            .O(N__4793),
            .I(N__4790));
    LocalMux I__488 (
            .O(N__4790),
            .I(\U712_CHIP_RAM.N_195_0 ));
    InMux I__487 (
            .O(N__4787),
            .I(N__4783));
    InMux I__486 (
            .O(N__4786),
            .I(N__4780));
    LocalMux I__485 (
            .O(N__4783),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ));
    LocalMux I__484 (
            .O(N__4780),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ));
    InMux I__483 (
            .O(N__4775),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__482 (
            .O(N__4772),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__481 (
            .O(N__4769),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__480 (
            .O(N__4766),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__479 (
            .O(N__4763),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__478 (
            .O(N__4760),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__477 (
            .O(N__4757),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    InMux I__476 (
            .O(N__4754),
            .I(N__4751));
    LocalMux I__475 (
            .O(N__4751),
            .I(\U712_CHIP_RAM.N_233 ));
    IoInMux I__474 (
            .O(N__4748),
            .I(N__4745));
    LocalMux I__473 (
            .O(N__4745),
            .I(N__4742));
    Span4Mux_s3_v I__472 (
            .O(N__4742),
            .I(N__4739));
    Span4Mux_v I__471 (
            .O(N__4739),
            .I(N__4736));
    Span4Mux_v I__470 (
            .O(N__4736),
            .I(N__4733));
    Span4Mux_v I__469 (
            .O(N__4733),
            .I(N__4729));
    InMux I__468 (
            .O(N__4732),
            .I(N__4726));
    Odrv4 I__467 (
            .O(N__4729),
            .I(DBDIR_c));
    LocalMux I__466 (
            .O(N__4726),
            .I(DBDIR_c));
    InMux I__465 (
            .O(N__4721),
            .I(N__4715));
    InMux I__464 (
            .O(N__4720),
            .I(N__4715));
    LocalMux I__463 (
            .O(N__4715),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    InMux I__462 (
            .O(N__4712),
            .I(N__4709));
    LocalMux I__461 (
            .O(N__4709),
            .I(N__4704));
    InMux I__460 (
            .O(N__4708),
            .I(N__4699));
    InMux I__459 (
            .O(N__4707),
            .I(N__4699));
    Span4Mux_v I__458 (
            .O(N__4704),
            .I(N__4694));
    LocalMux I__457 (
            .O(N__4699),
            .I(N__4694));
    Span4Mux_v I__456 (
            .O(N__4694),
            .I(N__4691));
    Span4Mux_v I__455 (
            .O(N__4691),
            .I(N__4688));
    Span4Mux_v I__454 (
            .O(N__4688),
            .I(N__4685));
    IoSpan4Mux I__453 (
            .O(N__4685),
            .I(N__4682));
    Odrv4 I__452 (
            .O(N__4682),
            .I(AWEn_c));
    InMux I__451 (
            .O(N__4679),
            .I(N__4676));
    LocalMux I__450 (
            .O(N__4676),
            .I(N__4673));
    Span4Mux_v I__449 (
            .O(N__4673),
            .I(N__4670));
    Sp12to4 I__448 (
            .O(N__4670),
            .I(N__4667));
    Span12Mux_h I__447 (
            .O(N__4667),
            .I(N__4664));
    Span12Mux_v I__446 (
            .O(N__4664),
            .I(N__4661));
    Odrv12 I__445 (
            .O(N__4661),
            .I(A_c_18));
    InMux I__444 (
            .O(N__4658),
            .I(N__4655));
    LocalMux I__443 (
            .O(N__4655),
            .I(N__4652));
    Span4Mux_v I__442 (
            .O(N__4652),
            .I(N__4649));
    Span4Mux_v I__441 (
            .O(N__4649),
            .I(N__4646));
    Sp12to4 I__440 (
            .O(N__4646),
            .I(N__4643));
    Odrv12 I__439 (
            .O(N__4643),
            .I(A_c_20));
    InMux I__438 (
            .O(N__4640),
            .I(N__4637));
    LocalMux I__437 (
            .O(N__4637),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0 ));
    IoInMux I__436 (
            .O(N__4634),
            .I(N__4631));
    LocalMux I__435 (
            .O(N__4631),
            .I(N__4628));
    Span4Mux_s3_v I__434 (
            .O(N__4628),
            .I(N__4625));
    Sp12to4 I__433 (
            .O(N__4625),
            .I(N__4622));
    Span12Mux_h I__432 (
            .O(N__4622),
            .I(N__4619));
    Span12Mux_v I__431 (
            .O(N__4619),
            .I(N__4615));
    InMux I__430 (
            .O(N__4618),
            .I(N__4612));
    Odrv12 I__429 (
            .O(N__4615),
            .I(CONSTANT_ONE_NET));
    LocalMux I__428 (
            .O(N__4612),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__427 (
            .O(N__4607),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ));
    CascadeMux I__426 (
            .O(N__4604),
            .I(\U712_CHIP_RAM.m104_ns_1_cascade_ ));
    CascadeMux I__425 (
            .O(N__4601),
            .I(\U712_CHIP_RAM.N_105_0_cascade_ ));
    InMux I__424 (
            .O(N__4598),
            .I(N__4595));
    LocalMux I__423 (
            .O(N__4595),
            .I(\U712_CHIP_RAM.N_106_0 ));
    CascadeMux I__422 (
            .O(N__4592),
            .I(\U712_CHIP_RAM.N_106_0_cascade_ ));
    InMux I__421 (
            .O(N__4589),
            .I(N__4586));
    LocalMux I__420 (
            .O(N__4586),
            .I(\U712_CHIP_RAM.DBENn_8_0 ));
    IoInMux I__419 (
            .O(N__4583),
            .I(N__4580));
    LocalMux I__418 (
            .O(N__4580),
            .I(N__4577));
    Span4Mux_s2_v I__417 (
            .O(N__4577),
            .I(N__4574));
    Span4Mux_v I__416 (
            .O(N__4574),
            .I(N__4571));
    Odrv4 I__415 (
            .O(N__4571),
            .I(CLK80_PLL_i_i));
    IoInMux I__414 (
            .O(N__4568),
            .I(N__4565));
    LocalMux I__413 (
            .O(N__4565),
            .I(N__4562));
    Odrv12 I__412 (
            .O(N__4562),
            .I(DBRn_c_i_0));
    InMux I__411 (
            .O(N__4559),
            .I(N__4556));
    LocalMux I__410 (
            .O(N__4556),
            .I(N__4553));
    Sp12to4 I__409 (
            .O(N__4553),
            .I(N__4550));
    Span12Mux_v I__408 (
            .O(N__4550),
            .I(N__4547));
    Odrv12 I__407 (
            .O(N__4547),
            .I(A_c_8));
    IoInMux I__406 (
            .O(N__4544),
            .I(N__4541));
    LocalMux I__405 (
            .O(N__4541),
            .I(N__4538));
    IoSpan4Mux I__404 (
            .O(N__4538),
            .I(N__4535));
    Span4Mux_s2_v I__403 (
            .O(N__4535),
            .I(N__4532));
    Span4Mux_v I__402 (
            .O(N__4532),
            .I(N__4529));
    Sp12to4 I__401 (
            .O(N__4529),
            .I(N__4525));
    InMux I__400 (
            .O(N__4528),
            .I(N__4522));
    Odrv12 I__399 (
            .O(N__4525),
            .I(LATCH_CLK_c));
    LocalMux I__398 (
            .O(N__4522),
            .I(LATCH_CLK_c));
    IoInMux I__397 (
            .O(N__4517),
            .I(N__4514));
    LocalMux I__396 (
            .O(N__4514),
            .I(N__4511));
    IoSpan4Mux I__395 (
            .O(N__4511),
            .I(N__4508));
    Span4Mux_s2_v I__394 (
            .O(N__4508),
            .I(N__4505));
    Sp12to4 I__393 (
            .O(N__4505),
            .I(N__4502));
    Span12Mux_v I__392 (
            .O(N__4502),
            .I(N__4499));
    Odrv12 I__391 (
            .O(N__4499),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__6935));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .I(N__6937));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__6940));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__6939));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .I(N__6941));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__6933));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__6934));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .I(N__6938));
    INV \INVU712_CYCLE_TERM.TACK_ENC  (
            .O(\INVU712_CYCLE_TERM.TACK_ENC_net ),
            .I(N__7231));
    INV \INVU712_CYCLE_TERM.TACK_OUTC  (
            .O(\INVU712_CYCLE_TERM.TACK_OUTC_net ),
            .I(N__7232));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .I(N__6932));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_13_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__7271),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7973),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4568),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__6563),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_2_1_0.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_2_1_0.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_2_1_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_2_1_0 (
            .in0(N__12134),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_11_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_11_7  (
            .in0(N__8215),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11645),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_6_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_6_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_6_LC_6_10_2  (
            .in0(N__4559),
            .in1(N__4787),
            .in2(_gnd_net_),
            .in3(N__4920),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12117),
            .ce(),
            .sr(N__11605));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_6_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_6_10_3 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_6_10_3  (
            .in0(N__4528),
            .in1(N__9790),
            .in2(N__6328),
            .in3(N__4640),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12117),
            .ce(),
            .sr(N__11605));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_6_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_6_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_6_10_5  (
            .in0(N__6312),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4618),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_6_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_6_10_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_6_10_6  (
            .in0(N__10995),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6311),
            .lcout(\U712_CHIP_RAM.m138_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_6_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_6_10_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_6_10_7  (
            .in0(N__4712),
            .in1(N__11424),
            .in2(_gnd_net_),
            .in3(N__6656),
            .lcout(\U712_CHIP_RAM.N_233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_6_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_6_11_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_6_11_0  (
            .in0(N__5645),
            .in1(N__5374),
            .in2(_gnd_net_),
            .in3(N__6650),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_6_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_6_11_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_LC_6_11_1  (
            .in0(N__6128),
            .in1(N__9783),
            .in2(N__4607),
            .in3(N__4598),
            .lcout(\U712_CHIP_RAM.DMA_CYCLEm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12123),
            .ce(),
            .sr(N__11598));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_6_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_6_11_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_6_11_2  (
            .in0(N__5644),
            .in1(N__6469),
            .in2(_gnd_net_),
            .in3(N__10679),
            .lcout(\U712_CHIP_RAM.DBENn_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIMF791_LC_6_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIMF791_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIMF791_LC_6_11_3 .LUT_INIT=16'b0001010110111111;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIMF791_LC_6_11_3  (
            .in0(N__6290),
            .in1(N__5114),
            .in2(N__5958),
            .in3(N__9782),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m104_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JFD6_0_LC_6_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JFD6_0_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JFD6_0_LC_6_11_4 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JFD6_0_LC_6_11_4  (
            .in0(N__5809),
            .in1(N__6291),
            .in2(N__4604),
            .in3(N__5458),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_105_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNINNJKA_LC_6_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNINNJKA_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNINNJKA_LC_6_11_5 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNINNJKA_LC_6_11_5  (
            .in0(N__6651),
            .in1(N__6495),
            .in2(N__4601),
            .in3(N__5643),
            .lcout(\U712_CHIP_RAM.N_106_0 ),
            .ltout(\U712_CHIP_RAM.N_106_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_6_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_6_11_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_6_11_6 .LUT_INIT=16'b0010101011101010;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_6_11_6  (
            .in0(N__9037),
            .in1(N__6129),
            .in2(N__4592),
            .in3(N__4589),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12123),
            .ce(),
            .sr(N__11598));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_6_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_6_11_7 .LUT_INIT=16'b0111111100100000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_6_11_7  (
            .in0(N__5375),
            .in1(N__4754),
            .in2(N__4877),
            .in3(N__5115),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12123),
            .ce(),
            .sr(N__11598));
    defparam \U712_CHIP_RAM.DBDIR_LC_6_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_6_12_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_6_12_1 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_6_12_1  (
            .in0(N__4707),
            .in1(N__4720),
            .in2(_gnd_net_),
            .in3(N__4732),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12127),
            .ce(),
            .sr(N__11591));
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_6_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_6_12_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_6_12_2 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_6_12_2  (
            .in0(N__4721),
            .in1(N__4708),
            .in2(_gnd_net_),
            .in3(N__11331),
            .lcout(\U712_CHIP_RAM.DMA_WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12127),
            .ce(),
            .sr(N__11591));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_7_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_7_9_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_7_LC_7_9_0  (
            .in0(N__4679),
            .in1(N__4921),
            .in2(_gnd_net_),
            .in3(N__7531),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12104),
            .ce(),
            .sr(N__11606));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_7_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_7_9_5 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_7_9_5  (
            .in0(N__4922),
            .in1(N__4658),
            .in2(N__11939),
            .in3(N__5413),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12104),
            .ce(),
            .sr(N__11606));
    defparam \U712_CHIP_RAM.REFRESH_RNIU7TF5_LC_7_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIU7TF5_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIU7TF5_LC_7_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIU7TF5_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__5372),
            .in2(_gnd_net_),
            .in3(N__5341),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNI50JL4_LC_7_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNI50JL4_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNI50JL4_LC_7_10_2 .LUT_INIT=16'b1011101000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNI50JL4_LC_7_10_2  (
            .in0(N__6655),
            .in1(N__6798),
            .in2(N__5498),
            .in3(N__5635),
            .lcout(\U712_CHIP_RAM.N_217_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_7_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_7_10_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_7_10_3  (
            .in0(N__6124),
            .in1(N__6470),
            .in2(_gnd_net_),
            .in3(N__5054),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_10_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_10_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_10_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_7_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_7_10_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_7_10_6  (
            .in0(N__10994),
            .in1(N__4786),
            .in2(_gnd_net_),
            .in3(N__10491),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_7_11_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_7_11_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__6324),
            .in2(_gnd_net_),
            .in3(N__4804),
            .lcout(\U712_CHIP_RAM.N_190_0 ),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_11_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_11_1  (
            .in0(N__4855),
            .in1(N__6462),
            .in2(_gnd_net_),
            .in3(N__4775),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__12118),
            .ce(N__5144),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_11_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__5164),
            .in2(_gnd_net_),
            .in3(N__4772),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_11_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_11_3  (
            .in0(N__4856),
            .in1(N__5947),
            .in2(_gnd_net_),
            .in3(N__4769),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__12118),
            .ce(N__5144),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_11_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_11_4  (
            .in0(N__4853),
            .in1(N__5189),
            .in2(_gnd_net_),
            .in3(N__4766),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__12118),
            .ce(N__5144),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_11_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_11_5  (
            .in0(N__4857),
            .in1(N__5596),
            .in2(_gnd_net_),
            .in3(N__4763),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__12118),
            .ce(N__5144),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_11_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_11_6  (
            .in0(N__4854),
            .in1(N__5569),
            .in2(_gnd_net_),
            .in3(N__4760),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__12118),
            .ce(N__5144),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_11_7  (
            .in0(N__4858),
            .in1(N__5201),
            .in2(_gnd_net_),
            .in3(N__4757),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12118),
            .ce(N__5144),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIJB9Q7_LC_7_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIJB9Q7_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIJB9Q7_LC_7_12_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_RNIJB9Q7_LC_7_12_0  (
            .in0(N__5450),
            .in1(N__9781),
            .in2(N__4811),
            .in3(N__6278),
            .lcout(\U712_CHIP_RAM.N_206_0 ),
            .ltout(\U712_CHIP_RAM.N_206_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOVP2B_1_LC_7_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOVP2B_1_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOVP2B_1_LC_7_12_1 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOVP2B_1_LC_7_12_1  (
            .in0(N__6279),
            .in1(N__6449),
            .in2(N__4892),
            .in3(N__6185),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_214_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIJR1UI_LC_7_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIJR1UI_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIJR1UI_LC_7_12_2 .LUT_INIT=16'b1111011111010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIJR1UI_LC_7_12_2  (
            .in0(N__9685),
            .in1(N__6101),
            .in2(N__4889),
            .in3(N__4817),
            .lcout(\U712_CHIP_RAM.N_216_0_i ),
            .ltout(\U712_CHIP_RAM.N_216_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_7_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_7_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_7_12_3 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_7_12_3  (
            .in0(N__4886),
            .in1(N__5294),
            .in2(N__4880),
            .in3(N__4876),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12124),
            .ce(N__5137),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_7_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_7_12_4 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_7_12_4  (
            .in0(N__9686),
            .in1(N__4859),
            .in2(N__5216),
            .in3(N__4829),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12124),
            .ce(N__5137),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_7_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_7_12_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_3_LC_7_12_5  (
            .in0(N__6277),
            .in1(N__5956),
            .in2(_gnd_net_),
            .in3(N__5869),
            .lcout(\U712_CHIP_RAM.N_195_0 ),
            .ltout(\U712_CHIP_RAM.N_195_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA1VV6_1_LC_7_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA1VV6_1_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA1VV6_1_LC_7_12_6 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIA1VV6_1_LC_7_12_6  (
            .in0(N__6448),
            .in1(N__5632),
            .in2(N__4820),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_213_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNICSPO4_LC_7_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNICSPO4_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNICSPO4_LC_7_12_7 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNICSPO4_LC_7_12_7  (
            .in0(N__5857),
            .in1(N__5449),
            .in2(_gnd_net_),
            .in3(N__5107),
            .lcout(\U712_CHIP_RAM.N_189_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_13_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_13_0 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_13_0  (
            .in0(N__6123),
            .in1(N__6496),
            .in2(_gnd_net_),
            .in3(N__4793),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12128),
            .ce(),
            .sr(N__11578));
    defparam DBRn_ibuf_RNIBAB_LC_7_14_1.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_7_14_1.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_7_14_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_7_14_1 (
            .in0(N__7729),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNI59L8_LC_8_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNI59L8_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNI59L8_LC_8_8_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNI59L8_LC_8_8_6  (
            .in0(N__11170),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11044),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_8_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_0_LC_8_9_0  (
            .in0(N__5030),
            .in1(N__5399),
            .in2(_gnd_net_),
            .in3(N__4923),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12097),
            .ce(),
            .sr(N__11599));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_8_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_8_9_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_3_LC_8_9_2  (
            .in0(N__5015),
            .in1(N__5387),
            .in2(_gnd_net_),
            .in3(N__4926),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12097),
            .ce(),
            .sr(N__11599));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_8_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_8_9_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_4_LC_8_9_3  (
            .in0(N__4927),
            .in1(N__4997),
            .in2(_gnd_net_),
            .in3(N__7516),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12097),
            .ce(),
            .sr(N__11599));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_8_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_8_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_1_LC_8_9_4  (
            .in0(N__4979),
            .in1(N__7672),
            .in2(_gnd_net_),
            .in3(N__4924),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12097),
            .ce(),
            .sr(N__11599));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_8_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_8_9_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_5_LC_8_9_5  (
            .in0(N__4928),
            .in1(N__4961),
            .in2(_gnd_net_),
            .in3(N__8522),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12097),
            .ce(),
            .sr(N__11599));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_8_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_8_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_2_LC_8_9_6  (
            .in0(N__4949),
            .in1(N__5426),
            .in2(_gnd_net_),
            .in3(N__4925),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12097),
            .ce(),
            .sr(N__11599));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_10_0 .LUT_INIT=16'b0100000011111111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_10_0  (
            .in0(N__6318),
            .in1(N__10973),
            .in2(N__6361),
            .in3(N__6447),
            .lcout(\U712_CHIP_RAM.N_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_0_3_LC_8_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_0_3_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_0_3_LC_8_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_0_3_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__5939),
            .in2(_gnd_net_),
            .in3(N__5863),
            .lcout(\U712_CHIP_RAM.N_111_0 ),
            .ltout(\U712_CHIP_RAM.N_111_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_10_2 .LUT_INIT=16'b0110010000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_10_2  (
            .in0(N__6317),
            .in1(N__6445),
            .in2(N__5084),
            .in3(N__5800),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_10_3 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_8_10_3  (
            .in0(N__6745),
            .in1(N__5081),
            .in2(N__6134),
            .in3(N__5063),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12105),
            .ce(),
            .sr(N__11592));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_10_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_10_4  (
            .in0(N__5312),
            .in1(N__6356),
            .in2(N__5957),
            .in3(N__5801),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_352_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_5 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_10_5  (
            .in0(N__6446),
            .in1(N__5075),
            .in2(N__5066),
            .in3(N__5272),
            .lcout(\U712_CHIP_RAM.N_183_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI2E2T2_LC_8_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI2E2T2_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI2E2T2_LC_8_10_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNI2E2T2_LC_8_10_6  (
            .in0(N__5940),
            .in1(N__5123),
            .in2(_gnd_net_),
            .in3(N__5799),
            .lcout(\U712_CHIP_RAM.N_137_0 ),
            .ltout(\U712_CHIP_RAM.N_137_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_10_7 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_8_10_7  (
            .in0(N__9809),
            .in1(N__6316),
            .in2(N__5057),
            .in3(N__5457),
            .lcout(\U712_CHIP_RAM.N_178_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_0_2_LC_8_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_0_2_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_0_2_LC_8_11_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_0_2_LC_8_11_0  (
            .in0(N__5559),
            .in1(N__5539),
            .in2(N__5165),
            .in3(N__5592),
            .lcout(\U712_CHIP_RAM.N_94_0 ),
            .ltout(\U712_CHIP_RAM.N_94_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_0_3_LC_8_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_0_3_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_0_3_LC_8_11_1 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_0_3_LC_8_11_1  (
            .in0(N__5924),
            .in1(_gnd_net_),
            .in2(N__5048),
            .in3(N__6258),
            .lcout(\U712_CHIP_RAM.N_96_0 ),
            .ltout(\U712_CHIP_RAM.N_96_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNI50JL4_0_LC_8_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNI50JL4_0_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNI50JL4_0_LC_8_11_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNI50JL4_0_LC_8_11_2  (
            .in0(N__6794),
            .in1(N__6649),
            .in2(N__5045),
            .in3(N__5488),
            .lcout(\U712_CHIP_RAM.N_188_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5NRT_7_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5NRT_7_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5NRT_7_LC_8_11_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5NRT_7_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__5200),
            .in2(_gnd_net_),
            .in3(N__5188),
            .lcout(\U712_CHIP_RAM.m92_0 ),
            .ltout(\U712_CHIP_RAM.m92_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_5_LC_8_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_5_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_5_LC_8_11_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_5_LC_8_11_4  (
            .in0(N__5557),
            .in1(N__5591),
            .in2(N__5177),
            .in3(N__5923),
            .lcout(\U712_CHIP_RAM.N_103_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_11_5 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_11_5  (
            .in0(N__6110),
            .in1(N__5174),
            .in2(N__6500),
            .in3(N__5340),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_11_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5168),
            .in3(N__11644),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_2_LC_8_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_2_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_2_LC_8_11_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI96LA2_2_LC_8_11_7  (
            .in0(N__5590),
            .in1(N__5160),
            .in2(N__5540),
            .in3(N__5558),
            .lcout(\U712_CHIP_RAM.N_110_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIO7T54_LC_8_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIO7T54_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIO7T54_LC_8_12_0 .LUT_INIT=16'b1000100010001100;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIO7T54_LC_8_12_0  (
            .in0(N__6584),
            .in1(N__5633),
            .in2(N__6802),
            .in3(N__5728),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_222_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_12_1 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_8_12_1  (
            .in0(N__6643),
            .in1(N__5972),
            .in2(N__5147),
            .in3(N__6096),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_8_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_8_12_2 .LUT_INIT=16'b1010000001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_8_12_2  (
            .in0(N__6268),
            .in1(N__6176),
            .in2(N__5881),
            .in3(N__6443),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_8_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_8_12_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__6267),
            .in2(_gnd_net_),
            .in3(N__5122),
            .lcout(\U712_CHIP_RAM.N_344 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_8_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_8_12_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIP7AQ_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__6442),
            .in2(_gnd_net_),
            .in3(N__6076),
            .lcout(\U712_CHIP_RAM.N_358 ),
            .ltout(\U712_CHIP_RAM.N_358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_8_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_8_12_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5297),
            .in3(N__9668),
            .lcout(\U712_CHIP_RAM.m219_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_8_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_8_12_6 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_8_12_6  (
            .in0(N__6269),
            .in1(N__5819),
            .in2(N__5810),
            .in3(N__6444),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_12_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__6097),
            .in2(N__5288),
            .in3(N__5285),
            .lcout(\U712_CHIP_RAM.N_117_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_13_0 .LUT_INIT=16'b1000100001010000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_13_0  (
            .in0(N__5477),
            .in1(N__5955),
            .in2(N__5279),
            .in3(N__6493),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_142_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_8_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_8_13_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_8_13_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_8_13_1  (
            .in0(N__6082),
            .in1(N__5242),
            .in2(N__5261),
            .in3(N__5231),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12125),
            .ce(),
            .sr(N__11577));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_8_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_8_13_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_8_13_2  (
            .in0(N__5471),
            .in1(N__6492),
            .in2(_gnd_net_),
            .in3(N__6295),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_8_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_8_13_3 .LUT_INIT=16'b0011000011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_8_13_3  (
            .in0(N__6360),
            .in1(N__5470),
            .in2(N__6503),
            .in3(N__6288),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m207_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_13_4 .LUT_INIT=16'b1100101001000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_13_4  (
            .in0(N__6494),
            .in1(N__6081),
            .in2(N__5225),
            .in3(N__5222),
            .lcout(\U712_CHIP_RAM.N_208_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_8_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_8_13_5 .LUT_INIT=16'b0001000111110101;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_2_LC_8_13_5  (
            .in0(N__6488),
            .in1(N__11100),
            .in2(N__5882),
            .in3(N__6289),
            .lcout(\U712_CHIP_RAM.m141_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_8_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_8_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__5954),
            .in2(_gnd_net_),
            .in3(N__5875),
            .lcout(\U712_CHIP_RAM.N_140_0 ),
            .ltout(\U712_CHIP_RAM.N_140_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIBDIU5_LC_8_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIBDIU5_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIBDIU5_LC_8_13_7 .LUT_INIT=16'b0001010110111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIBDIU5_LC_8_13_7  (
            .in0(N__6080),
            .in1(N__6287),
            .in2(N__5462),
            .in3(N__5459),
            .lcout(\U712_CHIP_RAM.m203_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_9_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_9_1  (
            .in0(N__5425),
            .in1(N__10960),
            .in2(_gnd_net_),
            .in3(N__10450),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_9_9_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_9_9_2  (
            .in0(N__10962),
            .in1(N__10440),
            .in2(_gnd_net_),
            .in3(N__5414),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_9_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_9_3  (
            .in0(N__5398),
            .in1(N__10961),
            .in2(_gnd_net_),
            .in3(N__10451),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_9_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_9_4  (
            .in0(N__10959),
            .in1(N__10439),
            .in2(_gnd_net_),
            .in3(N__5386),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__5373),
            .in2(_gnd_net_),
            .in3(N__5342),
            .lcout(\U712_CHIP_RAM.CPU_CYCLEm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12098),
            .ce(N__5324),
            .sr(N__11584));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_11_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__6481),
            .in2(_gnd_net_),
            .in3(N__5308),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m123_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_11_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_11_1  (
            .in0(N__6131),
            .in1(N__5634),
            .in2(N__5606),
            .in3(N__5874),
            .lcout(\U712_CHIP_RAM.N_125_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_11_2 .LUT_INIT=16'b1011000111111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_11_2  (
            .in0(N__6005),
            .in1(N__5603),
            .in2(N__8749),
            .in3(N__9566),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12106),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_0_5_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_0_5_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_0_5_LC_9_11_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIA7LA2_0_5_LC_9_11_3  (
            .in0(N__5597),
            .in1(N__5948),
            .in2(N__5570),
            .in3(N__5535),
            .lcout(\U712_CHIP_RAM.N_130_0 ),
            .ltout(\U712_CHIP_RAM.N_130_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG3845_0_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG3845_0_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG3845_0_LC_9_11_4 .LUT_INIT=16'b0011110000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIG3845_0_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__6322),
            .in2(N__5519),
            .in3(N__5796),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_RNIG3845Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_11_7 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_11_7  (
            .in0(N__6323),
            .in1(N__6180),
            .in2(N__6501),
            .in3(N__5873),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5_3_LC_9_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5_3_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5_3_LC_9_12_0 .LUT_INIT=16'b1000010110000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5_3_LC_9_12_0  (
            .in0(N__6326),
            .in1(N__5798),
            .in2(N__5966),
            .in3(N__5880),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIU9G4C_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIU9G4C_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIU9G4C_LC_9_12_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIU9G4C_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__5978),
            .in2(N__5516),
            .in3(N__5513),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_363_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2VCTI_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2VCTI_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2VCTI_LC_9_12_2 .LUT_INIT=16'b0101010111000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2VCTI_LC_9_12_2  (
            .in0(N__5507),
            .in1(N__6130),
            .in2(N__5501),
            .in3(N__6499),
            .lcout(\U712_CHIP_RAM.N_204_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNI4OCE_LC_9_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNI4OCE_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNI4OCE_LC_9_12_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNI4OCE_LC_9_12_3  (
            .in0(N__6576),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5726),
            .lcout(\U712_CHIP_RAM.m186_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_12_4 .LUT_INIT=16'b0011001100000001;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_12_4  (
            .in0(N__5727),
            .in1(N__6619),
            .in2(N__6803),
            .in3(N__6577),
            .lcout(\U712_CHIP_RAM.N_363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIK0QU_1_LC_9_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIK0QU_1_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIK0QU_1_LC_9_12_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIK0QU_1_LC_9_12_5  (
            .in0(N__6497),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9667),
            .lcout(\U712_CHIP_RAM.m225_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5_0_3_LC_9_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5_0_3_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5_0_3_LC_9_12_6 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIFR5J5_0_3_LC_9_12_6  (
            .in0(N__6325),
            .in1(N__5797),
            .in2(N__5965),
            .in3(N__5879),
            .lcout(\U712_CHIP_RAM.N_112_0 ),
            .ltout(\U712_CHIP_RAM.N_112_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_12_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_12_7  (
            .in0(N__6498),
            .in1(N__6327),
            .in2(N__5813),
            .in3(N__5805),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_13_2 .LUT_INIT=16'b0011011100000101;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_13_2  (
            .in0(N__5687),
            .in1(N__10992),
            .in2(N__5759),
            .in3(N__5729),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12119),
            .ce(),
            .sr(N__11573));
    defparam \U712_REG_SM.START_RST_LC_9_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.START_RST_LC_9_14_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_REG_SM.START_RST_LC_9_14_1  (
            .in0(N__5653),
            .in1(N__7746),
            .in2(_gnd_net_),
            .in3(N__7061),
            .lcout(U712_REG_SM_START_RST),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12126),
            .ce(),
            .sr(N__11570));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_14_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_14_3 .LUT_INIT=16'b0001111100010001;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_9_14_3  (
            .in0(N__5708),
            .in1(N__5683),
            .in2(N__5657),
            .in3(N__7002),
            .lcout(U712_REG_SM_REG_CYCLE_START),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12126),
            .ce(),
            .sr(N__11570));
    defparam \U712_CHIP_RAM.m69_LC_9_16_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m69_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m69_LC_9_16_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.m69_LC_9_16_5  (
            .in0(N__7441),
            .in1(N__6708),
            .in2(_gnd_net_),
            .in3(N__7318),
            .lcout(\U712_CHIP_RAM.N_326_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_0_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_0_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_0_LC_10_8_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_0_LC_10_8_3  (
            .in0(N__8354),
            .in1(N__10460),
            .in2(N__8744),
            .in3(N__10644),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_10_10_0 .LUT_INIT=16'b0000010100001011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_10_10_0  (
            .in0(N__8731),
            .in1(N__8350),
            .in2(N__10645),
            .in3(N__10441),
            .lcout(\U712_CHIP_RAM.N_168_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_10_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_10_10_2  (
            .in0(N__6502),
            .in1(N__6781),
            .in2(_gnd_net_),
            .in3(N__6647),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_359_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_10_10_3 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_10_10_3  (
            .in0(N__6362),
            .in1(N__6329),
            .in2(N__6188),
            .in3(N__6181),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_RNO_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(N__6132),
            .in2(N__6155),
            .in3(N__6152),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_135_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_5 .LUT_INIT=16'b1011101100111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_5  (
            .in0(N__10442),
            .in1(N__9679),
            .in2(N__6143),
            .in3(N__6008),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12095),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_11_1 .LUT_INIT=16'b1101000111111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_11_1  (
            .in0(N__6140),
            .in1(N__6007),
            .in2(N__8361),
            .in3(N__9564),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12099),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_5  (
            .in0(N__6133),
            .in1(N__6020),
            .in2(_gnd_net_),
            .in3(N__6014),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_120_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_6 .LUT_INIT=16'b1101111101010111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_6  (
            .in0(N__9565),
            .in1(N__6006),
            .in2(N__5981),
            .in3(N__10643),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12099),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_12_7 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_12_7  (
            .in0(N__9839),
            .in1(N__9813),
            .in2(N__6648),
            .in3(N__8962),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12107),
            .ce(),
            .sr(N__11574));
    defparam \U712_REG_SM.C3_SYNC_1_LC_10_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_10_13_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_10_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6521),
            .lcout(U712_REG_SM_C3_SYNC_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12112),
            .ce(),
            .sr(N__11571));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_13_1 .LUT_INIT=16'b1010101001110111;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_10_13_1  (
            .in0(N__8963),
            .in1(N__8483),
            .in2(_gnd_net_),
            .in3(N__8846),
            .lcout(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12112),
            .ce(),
            .sr(N__11571));
    defparam \U712_REG_SM.C3_SYNC_0_LC_10_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_10_13_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_10_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6550),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12112),
            .ce(),
            .sr(N__11571));
    defparam \U712_CHIP_RAM.m11_e_LC_10_14_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m11_e_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m11_e_LC_10_14_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.m11_e_LC_10_14_1  (
            .in0(N__6971),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6995),
            .lcout(\U712_CHIP_RAM.N_329 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m174_LC_10_14_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m174_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m174_LC_10_14_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.m174_LC_10_14_2  (
            .in0(N__8096),
            .in1(N__9349),
            .in2(N__7003),
            .in3(N__6972),
            .lcout(N_175_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m27_LC_10_14_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m27_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m27_LC_10_14_3 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U712_CHIP_RAM.m27_LC_10_14_3  (
            .in0(N__9351),
            .in1(N__7502),
            .in2(N__8123),
            .in3(N__8841),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_28_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_14_4 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_10_14_4  (
            .in0(N__9678),
            .in1(N__6512),
            .in2(N__6515),
            .in3(N__7063),
            .lcout(U712_REG_SM_STATE_COUNT_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12120),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m15_LC_10_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m15_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m15_LC_10_14_5 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \U712_CHIP_RAM.m15_LC_10_14_5  (
            .in0(N__9350),
            .in1(N__8097),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_16_0 ),
            .ltout(\U712_CHIP_RAM.N_16_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_10_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_10_14_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_10_14_6 .LUT_INIT=16'b0000101010001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_10_14_6  (
            .in0(N__9677),
            .in1(N__7750),
            .in2(N__6506),
            .in3(N__7062),
            .lcout(U712_REG_SM_STATE_COUNT_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12120),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m65_LC_10_15_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m65_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m65_LC_10_15_1 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \U712_CHIP_RAM.m65_LC_10_15_1  (
            .in0(N__7454),
            .in1(N__7320),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_66_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m173_LC_10_15_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m173_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m173_LC_10_15_2 .LUT_INIT=16'b0000000011111011;
    LogicCell40 \U712_CHIP_RAM.m173_LC_10_15_2  (
            .in0(N__11411),
            .in1(N__6730),
            .in2(N__6734),
            .in3(N__9356),
            .lcout(N_174_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m143_LC_10_16_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m143_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m143_LC_10_16_0 .LUT_INIT=16'b0011000111000100;
    LogicCell40 \U712_CHIP_RAM.m143_LC_10_16_0  (
            .in0(N__7365),
            .in1(N__7319),
            .in2(N__6717),
            .in3(N__7442),
            .lcout(N_144_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m67_LC_10_17_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m67_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m67_LC_10_17_5 .LUT_INIT=16'b0101101001001000;
    LogicCell40 \U712_CHIP_RAM.m67_LC_10_17_5  (
            .in0(N__7303),
            .in1(N__7364),
            .in2(N__7440),
            .in3(N__6731),
            .lcout(N_68_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_7_5 .LUT_INIT=16'b1111101100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_11_7_5  (
            .in0(N__12347),
            .in1(N__10517),
            .in2(N__11125),
            .in3(N__7547),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12081),
            .ce(N__10326),
            .sr(N__11593));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_8_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_8_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__6674),
            .in2(_gnd_net_),
            .in3(N__6668),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__6936),
            .ce(),
            .sr(N__6905));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_8_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_8_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__6854),
            .in2(_gnd_net_),
            .in3(N__6665),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__6936),
            .ce(),
            .sr(N__6905));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_8_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_8_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__6881),
            .in2(_gnd_net_),
            .in3(N__6662),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__6936),
            .ce(),
            .sr(N__6905));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_8_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_8_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__6893),
            .in2(_gnd_net_),
            .in3(N__6659),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__6936),
            .ce(),
            .sr(N__6905));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_8_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_8_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__6868),
            .in2(_gnd_net_),
            .in3(N__6953),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__6936),
            .ce(),
            .sr(N__6905));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_8_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_8_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__6815),
            .in2(_gnd_net_),
            .in3(N__6950),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__6936),
            .ce(),
            .sr(N__6905));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_8_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_8_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__6830),
            .in2(_gnd_net_),
            .in3(N__6947),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__6936),
            .ce(),
            .sr(N__6905));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_8_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_8_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__6842),
            .in2(_gnd_net_),
            .in3(N__6944),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6936),
            .ce(),
            .sr(N__6905));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_9_1 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_9_1  (
            .in0(N__6892),
            .in1(N__6880),
            .in2(N__6869),
            .in3(N__6853),
            .lcout(),
            .ltout(\U712_CHIP_RAM.REFRESH5lt7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_11_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_11_9_2  (
            .in0(N__6841),
            .in1(N__6829),
            .in2(N__6818),
            .in3(N__6814),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12086),
            .ce(),
            .sr(N__11579));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_0_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_0_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_0_LC_11_9_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_0_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__11643),
            .in2(_gnd_net_),
            .in3(N__6755),
            .lcout(\U712_CHIP_RAM.N_168_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_START_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_START_LC_11_10_0 .SEQ_MODE=4'b1010;
    defparam \U712_CYCLE_TERM.TACK_START_LC_11_10_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CYCLE_TERM.TACK_START_LC_11_10_0  (
            .in0(N__7829),
            .in1(N__6749),
            .in2(_gnd_net_),
            .in3(N__9462),
            .lcout(\U712_CYCLE_TERM.TACK_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12092),
            .ce(),
            .sr(N__7034));
    defparam \U712_CYCLE_TERM.TACK_START_RNO_0_LC_11_11_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_START_RNO_0_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_START_RNO_0_LC_11_11_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_START_RNO_0_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__9563),
            .in2(_gnd_net_),
            .in3(N__9416),
            .lcout(\U712_CYCLE_TERM.TACK_RST_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__9669),
            .in2(_gnd_net_),
            .in3(N__7103),
            .lcout(U712_REG_SM_STATE_COUNT_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12100),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_7_LC_11_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_7_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_7_LC_11_12_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_7_LC_11_12_3  (
            .in0(N__9671),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7016),
            .lcout(U712_REG_SM_STATE_COUNT_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12100),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m45_0_LC_11_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m45_0_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m45_0_LC_11_12_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.m45_0_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__7024),
            .in2(_gnd_net_),
            .in3(N__6973),
            .lcout(U712_CHIP_RAM_m45_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_11_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_11_12_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_11_12_7  (
            .in0(N__9670),
            .in1(_gnd_net_),
            .in2(N__7028),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12100),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m9_LC_11_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m9_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m9_LC_11_13_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.m9_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__8107),
            .in2(_gnd_net_),
            .in3(N__9362),
            .lcout(N_10_0),
            .ltout(N_10_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_11_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_11_13_1 .LUT_INIT=16'b0000110010001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_11_13_1  (
            .in0(N__7490),
            .in1(N__9675),
            .in2(N__7010),
            .in3(N__7778),
            .lcout(U712_REG_SM_STATE_COUNT_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12108),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m83_LC_11_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m83_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m83_LC_11_13_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.m83_LC_11_13_2  (
            .in0(N__7007),
            .in1(N__9363),
            .in2(_gnd_net_),
            .in3(N__8108),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_84_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_13_3 .LUT_INIT=16'b0011111110111011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_11_13_3  (
            .in0(N__7076),
            .in1(N__9674),
            .in2(N__6977),
            .in3(N__6974),
            .lcout(U712_REG_SM_STATE_COUNT_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12108),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m40_ns_LC_11_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m40_ns_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m40_ns_LC_11_13_4 .LUT_INIT=16'b1100000011000101;
    LogicCell40 \U712_CHIP_RAM.m40_ns_LC_11_13_4  (
            .in0(N__11150),
            .in1(N__7115),
            .in2(N__7808),
            .in3(N__7489),
            .lcout(),
            .ltout(i66_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_11_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_11_13_5 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_11_13_5  (
            .in0(N__9672),
            .in1(_gnd_net_),
            .in2(N__7118),
            .in3(N__11151),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12108),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m40_ns_1_LC_11_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m40_ns_1_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m40_ns_1_LC_11_13_6 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \U712_CHIP_RAM.m40_ns_1_LC_11_13_6  (
            .in0(N__8177),
            .in1(N__8106),
            .in2(_gnd_net_),
            .in3(N__9361),
            .lcout(\U712_CHIP_RAM.m40_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_13_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_11_13_7  (
            .in0(N__9673),
            .in1(N__7777),
            .in2(_gnd_net_),
            .in3(N__7109),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12108),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m32_LC_11_14_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m32_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m32_LC_11_14_0 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \U712_CHIP_RAM.m32_LC_11_14_0  (
            .in0(N__7057),
            .in1(N__9338),
            .in2(N__8113),
            .in3(N__7800),
            .lcout(N_33_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_8_LC_11_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_8_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_8_LC_11_14_1 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_8_LC_11_14_1  (
            .in0(N__7802),
            .in1(N__9676),
            .in2(N__7097),
            .in3(N__7085),
            .lcout(U712_REG_SM_STATE_COUNT_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12113),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m20_LC_11_14_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m20_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m20_LC_11_14_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.m20_LC_11_14_2  (
            .in0(N__8095),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9340),
            .lcout(\U712_CHIP_RAM.N_21_0 ),
            .ltout(\U712_CHIP_RAM.N_21_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m30_LC_11_14_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m30_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m30_LC_11_14_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U712_CHIP_RAM.m30_LC_11_14_3  (
            .in0(N__7801),
            .in1(_gnd_net_),
            .in2(N__7079),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_31_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m19_LC_11_14_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m19_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m19_LC_11_14_4 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \U712_CHIP_RAM.m19_LC_11_14_4  (
            .in0(N__8094),
            .in1(N__7070),
            .in2(N__7064),
            .in3(N__9339),
            .lcout(N_20_0),
            .ltout(N_20_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_ess_RNO_LC_11_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_ess_RNO_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REGENn_ess_RNO_LC_11_14_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_REG_SM.REGENn_ess_RNO_LC_11_14_5  (
            .in0(N__11642),
            .in1(_gnd_net_),
            .in2(N__7037),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.N_20_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m36_LC_11_14_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m36_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m36_LC_11_14_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.m36_LC_11_14_6  (
            .in0(N__7501),
            .in1(N__9341),
            .in2(N__8840),
            .in3(N__8109),
            .lcout(\U712_CHIP_RAM.N_37_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_15_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_11_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7241),
            .lcout(U712_REG_SM_C1_SYNC_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12121),
            .ce(),
            .sr(N__11563));
    defparam \U712_REG_SM.UDSn_LC_11_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_LC_11_15_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.UDSn_LC_11_15_6 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \U712_REG_SM.UDSn_LC_11_15_6  (
            .in0(N__7465),
            .in1(N__7481),
            .in2(_gnd_net_),
            .in3(N__8766),
            .lcout(UDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12121),
            .ce(),
            .sr(N__11563));
    defparam \U712_CHIP_RAM.m144_LC_11_16_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m144_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m144_LC_11_16_3 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \U712_CHIP_RAM.m144_LC_11_16_3  (
            .in0(N__7452),
            .in1(N__7366),
            .in2(N__7390),
            .in3(N__7333),
            .lcout(N_145_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m171_LC_11_16_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m171_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m171_LC_11_16_5 .LUT_INIT=16'b0000000010101111;
    LogicCell40 \U712_CHIP_RAM.m171_LC_11_16_5  (
            .in0(N__11398),
            .in1(_gnd_net_),
            .in2(N__7391),
            .in3(N__9355),
            .lcout(N_172_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m70_LC_11_16_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m70_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m70_LC_11_16_6 .LUT_INIT=16'b0101110010101100;
    LogicCell40 \U712_CHIP_RAM.m70_LC_11_16_6  (
            .in0(N__7453),
            .in1(N__7389),
            .in2(N__7370),
            .in3(N__7334),
            .lcout(N_71_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_17_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_17_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_11_17_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_11_17_4  (
            .in0(N__7267),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12129),
            .ce(),
            .sr(N__11557));
    defparam CLK40_PLL_derived_clock_RNIIOT_LC_12_1_5.C_ON=1'b0;
    defparam CLK40_PLL_derived_clock_RNIIOT_LC_12_1_5.SEQ_MODE=4'b0000;
    defparam CLK40_PLL_derived_clock_RNIIOT_LC_12_1_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLK40_PLL_derived_clock_RNIIOT_LC_12_1_5 (
            .in0(N__7209),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_iso_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_6_1 .LUT_INIT=16'b0000100011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_6_1  (
            .in0(N__8616),
            .in1(N__12203),
            .in2(N__11102),
            .in3(N__7682),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12078),
            .ce(N__10320),
            .sr(N__11590));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_7_1 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_7_1  (
            .in0(N__10038),
            .in1(N__7658),
            .in2(N__9707),
            .in3(N__7610),
            .lcout(\U712_CHIP_RAM.m154_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_8_2 .LUT_INIT=16'b1010101010111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_8_2  (
            .in0(N__10548),
            .in1(N__7676),
            .in2(N__11119),
            .in3(N__10232),
            .lcout(\U712_CHIP_RAM.m154_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_8_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_8_5  (
            .in0(N__11095),
            .in1(N__10549),
            .in2(N__10242),
            .in3(N__7642),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_2_LC_12_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_2_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_2_LC_12_8_6 .LUT_INIT=16'b0000000010111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_2_LC_12_8_6  (
            .in0(N__7591),
            .in1(N__11096),
            .in2(N__10570),
            .in3(N__10233),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m157_xx_mm_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_7 .LUT_INIT=16'b0101000000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_7  (
            .in0(N__7562),
            .in1(N__10034),
            .in2(N__7550),
            .in3(N__10766),
            .lcout(\U712_CHIP_RAM.m157_xx_mm_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_9_0 .LUT_INIT=16'b0101000000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_9_0  (
            .in0(N__7541),
            .in1(N__10020),
            .in2(N__8282),
            .in3(N__10694),
            .lcout(\U712_CHIP_RAM.m156_xx_mm_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_9_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_9_1  (
            .in0(N__7532),
            .in1(N__11093),
            .in2(_gnd_net_),
            .in3(N__10542),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_9_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_9_7  (
            .in0(N__7517),
            .in1(N__11094),
            .in2(_gnd_net_),
            .in3(N__10541),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_8_LC_12_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_8_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_8_LC_12_10_2 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_8_LC_12_10_2  (
            .in0(N__10996),
            .in1(N__10234),
            .in2(N__10540),
            .in3(N__7892),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m162_xx_mm_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_12_10_3 .LUT_INIT=16'b0011000000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_12_10_3  (
            .in0(N__10028),
            .in1(N__7877),
            .in2(N__7865),
            .in3(N__8191),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m162_xx_mm_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_10_4 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_12_10_4  (
            .in0(N__10997),
            .in1(N__10106),
            .in2(N__7862),
            .in3(N__10490),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12085),
            .ce(N__10293),
            .sr(N__11572));
    defparam \U712_REG_SM.REG_TACK_LC_12_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_12_12_4 .LUT_INIT=16'b0101110101010001;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_12_12_4  (
            .in0(N__7814),
            .in1(N__7835),
            .in2(N__7760),
            .in3(N__7825),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12094),
            .ce(),
            .sr(N__11568));
    defparam \U712_CHIP_RAM.m35_LC_12_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m35_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m35_LC_12_13_1 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \U712_CHIP_RAM.m35_LC_12_13_1  (
            .in0(N__7803),
            .in1(N__7776),
            .in2(_gnd_net_),
            .in3(N__8178),
            .lcout(U712_REG_SM_REG_TACK_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m43_LC_12_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m43_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m43_LC_12_13_3 .LUT_INIT=16'b0011100000001000;
    LogicCell40 \U712_CHIP_RAM.m43_LC_12_13_3  (
            .in0(N__7804),
            .in1(N__9364),
            .in2(N__8124),
            .in3(N__7775),
            .lcout(N_44_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.WRITE_CYCLE_LC_12_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_12_14_2 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \U712_REG_SM.WRITE_CYCLE_LC_12_14_2  (
            .in0(N__11425),
            .in1(N__7751),
            .in2(_gnd_net_),
            .in3(N__8179),
            .lcout(U712_REG_SM_WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12103),
            .ce(),
            .sr(N__11562));
    defparam DBR_SYNC_0_LC_12_14_4.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_12_14_4.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_12_14_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 DBR_SYNC_0_LC_12_14_4 (
            .in0(N__7730),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12103),
            .ce(),
            .sr(N__11562));
    defparam DBR_SYNC_1_LC_12_14_5.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_12_14_5.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_12_14_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_12_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7700),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12103),
            .ce(),
            .sr(N__11562));
    defparam \U712_REG_SM.PRnW_LC_12_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.PRnW_LC_12_14_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.PRnW_LC_12_14_7 .LUT_INIT=16'b1111110001011100;
    LogicCell40 \U712_REG_SM.PRnW_LC_12_14_7  (
            .in0(N__8180),
            .in1(N__8137),
            .in2(N__8159),
            .in3(N__8126),
            .lcout(PRnW_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12103),
            .ce(),
            .sr(N__11562));
    defparam \U712_REG_SM.REGENn_ess_LC_12_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_ess_LC_12_15_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_ess_LC_12_15_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_REG_SM.REGENn_ess_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__8125),
            .in2(_gnd_net_),
            .in3(N__9360),
            .lcout(BLSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12111),
            .ce(N__8012),
            .sr(N__11558));
    defparam \U712_REG_SM.LDSn_LC_12_16_1 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_LC_12_16_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.LDSn_LC_12_16_1 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_REG_SM.LDSn_LC_12_16_1  (
            .in0(N__8000),
            .in1(N__7984),
            .in2(_gnd_net_),
            .in3(N__8774),
            .lcout(LDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12116),
            .ce(),
            .sr(N__11556));
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_5.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_5.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9666),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WEn_LC_13_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_13_6_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_13_6_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_13_6_6  (
            .in0(N__8366),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12080),
            .ce(),
            .sr(N__11600));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_1_LC_13_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_1_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_1_LC_13_7_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_1_LC_13_7_0  (
            .in0(N__10539),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10241),
            .lcout(\U712_CHIP_RAM.m164_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_7_LC_13_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_7_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_7_LC_13_8_0 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_7_LC_13_8_0  (
            .in0(N__11065),
            .in1(N__10227),
            .in2(N__10568),
            .in3(N__7937),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m161_xx_mm_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_8_1 .LUT_INIT=16'b0011000000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_8_1  (
            .in0(N__10032),
            .in1(N__7919),
            .in2(N__7913),
            .in3(N__9695),
            .lcout(\U712_CHIP_RAM.m161_xx_mm_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_4_LC_13_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_4_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_4_LC_13_8_3 .LUT_INIT=16'b0100010101010101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_4_LC_13_8_3  (
            .in0(N__10228),
            .in1(N__7910),
            .in2(N__10571),
            .in3(N__11066),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m159_xx_mm_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_8_4 .LUT_INIT=16'b0101000000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_8_4  (
            .in0(N__8423),
            .in1(N__10033),
            .in2(N__8417),
            .in3(N__9851),
            .lcout(\U712_CHIP_RAM.m159_xx_mm_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_6_LC_13_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_6_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_6_LC_13_8_6 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_6_LC_13_8_6  (
            .in0(N__8414),
            .in1(N__10226),
            .in2(N__11108),
            .in3(N__10553),
            .lcout(\U712_CHIP_RAM.m160_xx_mm_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_9_0 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_13_9_0  (
            .in0(N__11735),
            .in1(N__11114),
            .in2(N__8393),
            .in3(N__10544),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12087),
            .ce(N__10315),
            .sr(N__11580));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_9_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__8748),
            .in2(_gnd_net_),
            .in3(N__8362),
            .lcout(\U712_CHIP_RAM.N_3_0 ),
            .ltout(\U712_CHIP_RAM.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_0_LC_13_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_0_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_0_LC_13_9_2 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_0_LC_13_9_2  (
            .in0(N__8320),
            .in1(N__11113),
            .in2(N__8285),
            .in3(N__10543),
            .lcout(\U712_CHIP_RAM.m156_xx_mm_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNI8DDB1_LC_13_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNI8DDB1_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNI8DDB1_LC_13_10_1 .LUT_INIT=16'b1010111100100011;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNI8DDB1_LC_13_10_1  (
            .in0(N__8266),
            .in1(N__9746),
            .in2(N__11058),
            .in3(N__9072),
            .lcout(CLMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_13_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_13_10_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIHMEA_1_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(N__10993),
            .in2(_gnd_net_),
            .in3(N__10461),
            .lcout(\U712_CHIP_RAM.m154_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_11_0 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_11_0  (
            .in0(N__10837),
            .in1(N__11924),
            .in2(N__8219),
            .in3(N__8192),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .ce(),
            .sr(N__11575));
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_13_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_13_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_13_12_0 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_2_LC_13_12_0  (
            .in0(N__9619),
            .in1(N__8504),
            .in2(N__8956),
            .in3(N__8845),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12101),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_13_13_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_13_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__8431),
            .in2(N__8791),
            .in3(N__8792),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_13_13_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_13_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__8464),
            .in2(_gnd_net_),
            .in3(N__8507),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_13_13_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_13_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__8491),
            .in2(_gnd_net_),
            .in3(N__8498),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_13_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_13_13_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__8446),
            .in2(_gnd_net_),
            .in3(N__8495),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_13_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_13_13_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_13_13_4  (
            .in0(N__8447),
            .in1(N__8492),
            .in2(N__8468),
            .in3(N__8432),
            .lcout(\U712_CHIP_RAM.N_325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_13_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_13_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_13_13_5 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_1_LC_13_13_5  (
            .in0(N__9621),
            .in1(N__8474),
            .in2(N__8958),
            .in3(N__8839),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12109),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_13_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_13_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_13_13_6 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_3_LC_13_13_6  (
            .in0(N__8837),
            .in1(N__9622),
            .in2(N__8456),
            .in3(N__8949),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12109),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_13_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_13_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_13_13_7 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_0_LC_13_13_7  (
            .in0(N__9620),
            .in1(N__8438),
            .in2(N__8957),
            .in3(N__8838),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12109),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_RNITKK4_1_LC_13_14_1.C_ON=1'b0;
    defparam DBR_SYNC_RNITKK4_1_LC_13_14_1.SEQ_MODE=4'b0000;
    defparam DBR_SYNC_RNITKK4_1_LC_13_14_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBR_SYNC_RNITKK4_1_LC_13_14_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8824),
            .lcout(DBR_SYNC_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_RNO_LC_13_16_3 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_13_16_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.ASn_ess_RNO_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(N__11641),
            .in2(_gnd_net_),
            .in3(N__8773),
            .lcout(\U712_REG_SM.N_33_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RASn_LC_14_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_14_4_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_14_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_14_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8750),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12079),
            .ce(),
            .sr(N__11619));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1  (
            .in0(N__8618),
            .in1(N__8681),
            .in2(N__11103),
            .in3(N__10787),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12082),
            .ce(N__10319),
            .sr(N__11607));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_7_5 .LUT_INIT=16'b0100010000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_7_5  (
            .in0(N__8639),
            .in1(N__8624),
            .in2(N__10045),
            .in3(N__9218),
            .lcout(\U712_CHIP_RAM.m160_xx_mm_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_14_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_14_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_14_8_1 .LUT_INIT=16'b0000100011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_14_8_1  (
            .in0(N__8617),
            .in1(N__9212),
            .in2(N__11131),
            .in3(N__9182),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12088),
            .ce(N__10321),
            .sr(N__11594));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_8_5 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_14_8_5  (
            .in0(N__10775),
            .in1(N__11124),
            .in2(N__8579),
            .in3(N__10535),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12088),
            .ce(N__10321),
            .sr(N__11594));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_8_6 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_14_8_6  (
            .in0(N__10534),
            .in1(N__11123),
            .in2(N__8552),
            .in3(N__9863),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12088),
            .ce(N__10321),
            .sr(N__11594));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_14_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_14_9_1 .LUT_INIT=16'b1111111100010101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_14_9_1  (
            .in0(N__10224),
            .in1(N__8521),
            .in2(N__11129),
            .in3(N__10530),
            .lcout(\U712_CHIP_RAM.m155_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_9_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_9_4  (
            .in0(N__9206),
            .in1(N__10225),
            .in2(N__10567),
            .in3(N__11112),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_9_5 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_9_5  (
            .in0(N__10021),
            .in1(N__9191),
            .in2(N__9185),
            .in3(N__9857),
            .lcout(\U712_CHIP_RAM.m155_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNI8DDB1_0_LC_14_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNI8DDB1_0_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNI8DDB1_0_LC_14_10_3 .LUT_INIT=16'b0111000001110111;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNI8DDB1_0_LC_14_10_3  (
            .in0(N__9073),
            .in1(N__9742),
            .in2(N__9172),
            .in3(N__11001),
            .lcout(CUUBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNI6U6F1_LC_14_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNI6U6F1_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNI6U6F1_LC_14_11_0 .LUT_INIT=16'b1100111101000101;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNI6U6F1_LC_14_11_0  (
            .in0(N__9824),
            .in1(N__9122),
            .in2(N__11130),
            .in3(N__9053),
            .lcout(CLLBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNI6U6F1_0_LC_14_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNI6U6F1_0_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNI6U6F1_0_LC_14_11_1 .LUT_INIT=16'b0111000001110111;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNI6U6F1_0_LC_14_11_1  (
            .in0(N__9052),
            .in1(N__9823),
            .in2(N__9020),
            .in3(N__11115),
            .lcout(CUMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_14_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_14_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_14_12_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_14_12_0  (
            .in0(N__11286),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11224),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12110),
            .ce(),
            .sr(N__11576));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_14_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_14_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_14_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_14_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8969),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12110),
            .ce(),
            .sr(N__11576));
    defparam \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_14_13_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_14_13_3 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_14_13_3  (
            .in0(N__9486),
            .in1(N__9508),
            .in2(_gnd_net_),
            .in3(N__9471),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_36_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUT_LC_14_13_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUT_LC_14_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_OUT_LC_14_13_4 .LUT_INIT=16'b1011111110110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUT_LC_14_13_4  (
            .in0(N__9511),
            .in1(N__9632),
            .in2(N__8915),
            .in3(N__8864),
            .lcout(TACK_OUT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_14_13_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_14_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_14_13_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_14_13_5  (
            .in0(N__9633),
            .in1(N__9510),
            .in2(N__9491),
            .in3(N__9472),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_14_13_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_14_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_14_13_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_14_13_6  (
            .in0(N__9509),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9634),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_OUTC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_LC_14_14_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_14_14_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_14_14_0 .LUT_INIT=16'b0011000100110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_LC_14_14_0  (
            .in0(N__9512),
            .in1(N__9490),
            .in2(N__9406),
            .in3(N__9473),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CYCLE_TERM.TACK_ENC_net ),
            .ce(),
            .sr(N__11569));
    defparam \U712_REG_SM.ASn_ess_LC_14_16_6 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_LC_14_16_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_ess_LC_14_16_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.ASn_ess_LC_14_16_6  (
            .in0(N__9368),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12130),
            .ce(N__9266),
            .sr(N__11564));
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIVHJN_LC_14_19_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIVHJN_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIVHJN_LC_14_19_3 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIVHJN_LC_14_19_3  (
            .in0(N__11223),
            .in1(N__11293),
            .in2(_gnd_net_),
            .in3(N__11354),
            .lcout(DMA_LATCH_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_15_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_15_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_15_6_4 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_15_6_4  (
            .in0(N__9875),
            .in1(N__11048),
            .in2(N__10574),
            .in3(N__9239),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12083),
            .ce(N__10328),
            .sr(N__11615));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_7_5  (
            .in0(N__9970),
            .in1(N__11919),
            .in2(_gnd_net_),
            .in3(N__10154),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__11689),
            .sr(N__11608));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_8_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_8_5  (
            .in0(N__9926),
            .in1(N__11928),
            .in2(_gnd_net_),
            .in3(N__10750),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11723),
            .ce(N__11687),
            .sr(N__11601));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_8_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_8_7  (
            .in0(N__9969),
            .in1(N__11929),
            .in2(_gnd_net_),
            .in3(N__10153),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11723),
            .ce(N__11687),
            .sr(N__11601));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_9_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_9_0  (
            .in0(N__9968),
            .in1(N__11927),
            .in2(_gnd_net_),
            .in3(N__9922),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__11684),
            .sr(N__11595));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_10_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_10_6  (
            .in0(N__10751),
            .in1(N__11926),
            .in2(_gnd_net_),
            .in3(N__9915),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__11682),
            .sr(N__11585));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_15_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_15_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__10091),
            .in2(_gnd_net_),
            .in3(N__10078),
            .lcout(\U712_CHIP_RAM.m228_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIMKV8_LC_15_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIMKV8_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIMKV8_LC_15_11_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_RNIMKV8_LC_15_11_6  (
            .in0(N__9815),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11300),
            .lcout(\U712_CHIP_RAM.N_343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIVA8H_LC_15_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIVA8H_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_RNIVA8H_LC_15_12_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_RNIVA8H_LC_15_12_7  (
            .in0(_gnd_net_),
            .in1(N__11234),
            .in2(_gnd_net_),
            .in3(N__9814),
            .lcout(\U712_CHIP_RAM.N_342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_3_LC_16_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_3_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_3_LC_16_6_7 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_3_LC_16_6_7  (
            .in0(N__9725),
            .in1(N__10244),
            .in2(N__11101),
            .in3(N__10557),
            .lcout(\U712_CHIP_RAM.m158_xx_mm_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_16_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_16_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_16_7_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_16_7_0  (
            .in0(N__12338),
            .in1(N__11918),
            .in2(_gnd_net_),
            .in3(N__12242),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__11692),
            .sr(N__11616));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_8_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_8_2  (
            .in0(N__10145),
            .in1(N__11902),
            .in2(_gnd_net_),
            .in3(N__10838),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__11690),
            .sr(N__11609));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_16_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_16_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_16_9_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_16_9_5  (
            .in0(N__10243),
            .in1(N__10657),
            .in2(_gnd_net_),
            .in3(N__10569),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12102),
            .ce(N__10325),
            .sr(N__11602));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_10_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_10_4  (
            .in0(N__10829),
            .in1(N__11894),
            .in2(_gnd_net_),
            .in3(N__10146),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11718),
            .ce(N__11685),
            .sr(N__11596));
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_16_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_16_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_16_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_2_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12146),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12114),
            .ce(),
            .sr(N__11586));
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_16_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_16_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_16_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_3_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10097),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12114),
            .ce(),
            .sr(N__11586));
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_16_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_16_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_16_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_5_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10079),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12114),
            .ce(),
            .sr(N__11586));
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_16_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_16_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_16_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_4_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10085),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12114),
            .ce(),
            .sr(N__11586));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_17_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_17_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_17_6_3 .LUT_INIT=16'b0100010000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_17_6_3  (
            .in0(N__10067),
            .in1(N__10052),
            .in2(N__10046),
            .in3(N__10706),
            .lcout(\U712_CHIP_RAM.m158_xx_mm_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_7_4  (
            .in0(N__11870),
            .in1(N__9971),
            .in2(_gnd_net_),
            .in3(N__9914),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11722),
            .ce(N__11694),
            .sr(N__11620));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_8_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_8_0  (
            .in0(N__10833),
            .in1(_gnd_net_),
            .in2(N__11923),
            .in3(N__12175),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11720),
            .ce(N__11693),
            .sr(N__11617));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_17_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_17_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_17_8_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_17_8_5  (
            .in0(N__10749),
            .in1(N__11895),
            .in2(_gnd_net_),
            .in3(N__12302),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11720),
            .ce(N__11693),
            .sr(N__11617));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_17_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_17_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_17_9_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_17_9_1  (
            .in0(N__11893),
            .in1(N__12301),
            .in2(_gnd_net_),
            .in3(N__12333),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__11691),
            .sr(N__11610));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_17_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_17_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_17_10_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_17_10_4  (
            .in0(N__12300),
            .in1(N__11892),
            .in2(_gnd_net_),
            .in3(N__10739),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__11688),
            .sr(N__11603));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_17_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_17_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_17_11_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_17_11_1  (
            .in0(N__12238),
            .in1(N__11817),
            .in2(_gnd_net_),
            .in3(N__11764),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__11683),
            .sr(N__11597));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_17_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_17_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_17_11_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_17_11_5  (
            .in0(N__11972),
            .in1(N__11816),
            .in2(_gnd_net_),
            .in3(N__11763),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__11683),
            .sr(N__11597));
    defparam \U712_CHIP_RAM.CRCSn_LC_18_3_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_18_3_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_18_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_18_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10664),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12084),
            .ce(),
            .sr(N__11625));
    defparam \U712_CHIP_RAM.CASn_LC_18_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_18_5_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_18_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_18_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10573),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12093),
            .ce(),
            .sr(N__11624));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_18_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_18_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_18_6_0 .LUT_INIT=16'b1111101100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_18_6_0  (
            .in0(N__12251),
            .in1(N__10572),
            .in2(N__11104),
            .in3(N__10352),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12096),
            .ce(N__10327),
            .sr(N__11623));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_18_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_18_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_18_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_18_7_5  (
            .in0(N__12234),
            .in1(N__11869),
            .in2(_gnd_net_),
            .in3(N__12332),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11721),
            .ce(N__11696),
            .sr(N__11622));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_18_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_18_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_18_8_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_18_8_3  (
            .in0(N__12334),
            .in1(_gnd_net_),
            .in2(N__11925),
            .in3(N__12299),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11719),
            .ce(N__11695),
            .sr(N__11621));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_18_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_18_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_18_8_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_18_8_6  (
            .in0(N__11768),
            .in1(N__11903),
            .in2(_gnd_net_),
            .in3(N__12233),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11719),
            .ce(N__11695),
            .sr(N__11621));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_18_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_18_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_18_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_18_9_6  (
            .in0(N__12188),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12176),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12115),
            .ce(),
            .sr(N__11618));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_18_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_18_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_18_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_18_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12152),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12122),
            .ce(),
            .sr(N__11611));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_18_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_18_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_18_11_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_18_11_1  (
            .in0(N__11971),
            .in1(N__11815),
            .in2(_gnd_net_),
            .in3(N__11754),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11717),
            .ce(N__11686),
            .sr(N__11604));
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIRVG61_LC_24_19_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIRVG61_LC_24_19_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIRVG61_LC_24_19_5 .LUT_INIT=16'b0000100001111111;
    LogicCell40 \U712_CHIP_RAM.DMA_WRITE_CYCLE_RNIRVG61_LC_24_19_5  (
            .in0(N__11219),
            .in1(N__11280),
            .in2(N__11429),
            .in3(N__11353),
            .lcout(N_323_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIQ44J_LC_24_19_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIQ44J_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIQ44J_LC_24_19_6 .LUT_INIT=16'b0000111100001000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNIQ44J_LC_24_19_6  (
            .in0(N__11279),
            .in1(N__11218),
            .in2(N__11177),
            .in3(N__11132),
            .lcout(N_333_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Nov 28 2024 19:11:39

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    A,
    RnW,
    TT1,
    TICK50,
    nROMEN,
    nCIACS1,
    TT0,
    TICK60,
    LBENn,
    CLKCIA,
    CLK6,
    CLK40_IN,
    CLK28_IN,
    TSn,
    nBUFEN,
    nREGSPACE,
    nRAMSPACE,
    RESETn,
    OVL,
    TACKn,
    nCIACS0,
    PORTSIZE);

    input [31:1] A;
    input RnW;
    input TT1;
    output TICK50;
    output nROMEN;
    output nCIACS1;
    input TT0;
    output TICK60;
    input LBENn;
    output CLKCIA;
    input CLK6;
    input CLK40_IN;
    input CLK28_IN;
    input TSn;
    output nBUFEN;
    output nREGSPACE;
    output nRAMSPACE;
    input RESETn;
    input OVL;
    inout TACKn;
    output nCIACS0;
    output PORTSIZE;

    wire N__6367;
    wire N__6366;
    wire N__6365;
    wire N__6357;
    wire N__6356;
    wire N__6355;
    wire N__6346;
    wire N__6345;
    wire N__6344;
    wire N__6337;
    wire N__6336;
    wire N__6335;
    wire N__6328;
    wire N__6327;
    wire N__6326;
    wire N__6319;
    wire N__6318;
    wire N__6317;
    wire N__6310;
    wire N__6309;
    wire N__6308;
    wire N__6301;
    wire N__6300;
    wire N__6299;
    wire N__6292;
    wire N__6291;
    wire N__6290;
    wire N__6283;
    wire N__6282;
    wire N__6281;
    wire N__6274;
    wire N__6273;
    wire N__6272;
    wire N__6265;
    wire N__6264;
    wire N__6263;
    wire N__6256;
    wire N__6255;
    wire N__6254;
    wire N__6247;
    wire N__6246;
    wire N__6245;
    wire N__6238;
    wire N__6237;
    wire N__6236;
    wire N__6229;
    wire N__6228;
    wire N__6227;
    wire N__6220;
    wire N__6219;
    wire N__6218;
    wire N__6211;
    wire N__6210;
    wire N__6209;
    wire N__6202;
    wire N__6201;
    wire N__6200;
    wire N__6193;
    wire N__6192;
    wire N__6191;
    wire N__6184;
    wire N__6183;
    wire N__6182;
    wire N__6175;
    wire N__6174;
    wire N__6173;
    wire N__6166;
    wire N__6165;
    wire N__6164;
    wire N__6157;
    wire N__6156;
    wire N__6155;
    wire N__6148;
    wire N__6147;
    wire N__6146;
    wire N__6139;
    wire N__6138;
    wire N__6137;
    wire N__6130;
    wire N__6129;
    wire N__6128;
    wire N__6121;
    wire N__6120;
    wire N__6119;
    wire N__6112;
    wire N__6111;
    wire N__6110;
    wire N__6103;
    wire N__6102;
    wire N__6101;
    wire N__6094;
    wire N__6093;
    wire N__6092;
    wire N__6085;
    wire N__6084;
    wire N__6083;
    wire N__6076;
    wire N__6075;
    wire N__6074;
    wire N__6067;
    wire N__6066;
    wire N__6065;
    wire N__6058;
    wire N__6057;
    wire N__6056;
    wire N__6039;
    wire N__6036;
    wire N__6035;
    wire N__6034;
    wire N__6033;
    wire N__6030;
    wire N__6027;
    wire N__6024;
    wire N__6021;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6002;
    wire N__6001;
    wire N__6000;
    wire N__5999;
    wire N__5998;
    wire N__5997;
    wire N__5994;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5982;
    wire N__5975;
    wire N__5972;
    wire N__5961;
    wire N__5960;
    wire N__5957;
    wire N__5956;
    wire N__5955;
    wire N__5952;
    wire N__5951;
    wire N__5950;
    wire N__5945;
    wire N__5938;
    wire N__5935;
    wire N__5928;
    wire N__5925;
    wire N__5924;
    wire N__5923;
    wire N__5920;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5900;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5886;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5874;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5866;
    wire N__5865;
    wire N__5862;
    wire N__5859;
    wire N__5856;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5843;
    wire N__5842;
    wire N__5841;
    wire N__5840;
    wire N__5839;
    wire N__5838;
    wire N__5835;
    wire N__5834;
    wire N__5833;
    wire N__5832;
    wire N__5829;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5809;
    wire N__5806;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5792;
    wire N__5785;
    wire N__5778;
    wire N__5775;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5757;
    wire N__5754;
    wire N__5751;
    wire N__5750;
    wire N__5749;
    wire N__5746;
    wire N__5745;
    wire N__5742;
    wire N__5739;
    wire N__5736;
    wire N__5733;
    wire N__5730;
    wire N__5727;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5709;
    wire N__5706;
    wire N__5703;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5682;
    wire N__5681;
    wire N__5680;
    wire N__5677;
    wire N__5672;
    wire N__5667;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5652;
    wire N__5651;
    wire N__5650;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5638;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5622;
    wire N__5619;
    wire N__5618;
    wire N__5617;
    wire N__5614;
    wire N__5613;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5586;
    wire N__5583;
    wire N__5582;
    wire N__5581;
    wire N__5580;
    wire N__5577;
    wire N__5574;
    wire N__5569;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5552;
    wire N__5551;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5529;
    wire N__5526;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5516;
    wire N__5515;
    wire N__5514;
    wire N__5513;
    wire N__5512;
    wire N__5509;
    wire N__5504;
    wire N__5499;
    wire N__5496;
    wire N__5487;
    wire N__5484;
    wire N__5481;
    wire N__5478;
    wire N__5475;
    wire N__5472;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5460;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5442;
    wire N__5441;
    wire N__5438;
    wire N__5437;
    wire N__5434;
    wire N__5433;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5406;
    wire N__5403;
    wire N__5400;
    wire N__5397;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5367;
    wire N__5364;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5349;
    wire N__5346;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5334;
    wire N__5331;
    wire N__5330;
    wire N__5329;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5315;
    wire N__5314;
    wire N__5311;
    wire N__5306;
    wire N__5301;
    wire N__5298;
    wire N__5295;
    wire N__5292;
    wire N__5289;
    wire N__5286;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5274;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5262;
    wire N__5259;
    wire N__5256;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5213;
    wire N__5212;
    wire N__5211;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5196;
    wire N__5187;
    wire N__5186;
    wire N__5185;
    wire N__5184;
    wire N__5183;
    wire N__5180;
    wire N__5179;
    wire N__5172;
    wire N__5165;
    wire N__5160;
    wire N__5159;
    wire N__5158;
    wire N__5157;
    wire N__5154;
    wire N__5151;
    wire N__5148;
    wire N__5145;
    wire N__5142;
    wire N__5139;
    wire N__5134;
    wire N__5127;
    wire N__5124;
    wire N__5121;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5102;
    wire N__5101;
    wire N__5100;
    wire N__5099;
    wire N__5094;
    wire N__5087;
    wire N__5082;
    wire N__5079;
    wire N__5078;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire N__5044;
    wire N__5043;
    wire N__5038;
    wire N__5035;
    wire N__5032;
    wire N__5027;
    wire N__5024;
    wire N__5023;
    wire N__5020;
    wire N__5017;
    wire N__5014;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4968;
    wire N__4967;
    wire N__4966;
    wire N__4965;
    wire N__4964;
    wire N__4963;
    wire N__4962;
    wire N__4961;
    wire N__4952;
    wire N__4949;
    wire N__4942;
    wire N__4935;
    wire N__4934;
    wire N__4933;
    wire N__4932;
    wire N__4931;
    wire N__4930;
    wire N__4925;
    wire N__4924;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4912;
    wire N__4909;
    wire N__4900;
    wire N__4893;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4881;
    wire N__4880;
    wire N__4879;
    wire N__4878;
    wire N__4877;
    wire N__4876;
    wire N__4875;
    wire N__4874;
    wire N__4863;
    wire N__4856;
    wire N__4851;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4839;
    wire N__4838;
    wire N__4837;
    wire N__4836;
    wire N__4835;
    wire N__4834;
    wire N__4833;
    wire N__4832;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4805;
    wire N__4804;
    wire N__4801;
    wire N__4798;
    wire N__4795;
    wire N__4788;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4755;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4743;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4731;
    wire N__4730;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4718;
    wire N__4715;
    wire N__4710;
    wire N__4707;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4689;
    wire N__4688;
    wire N__4685;
    wire N__4682;
    wire N__4677;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4665;
    wire N__4664;
    wire N__4661;
    wire N__4660;
    wire N__4659;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4623;
    wire N__4620;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4575;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4530;
    wire N__4529;
    wire N__4528;
    wire N__4527;
    wire N__4526;
    wire N__4523;
    wire N__4518;
    wire N__4513;
    wire N__4506;
    wire N__4505;
    wire N__4504;
    wire N__4503;
    wire N__4496;
    wire N__4493;
    wire N__4488;
    wire N__4485;
    wire N__4482;
    wire N__4481;
    wire N__4480;
    wire N__4479;
    wire N__4472;
    wire N__4469;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4443;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4431;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4373;
    wire N__4372;
    wire N__4369;
    wire N__4366;
    wire N__4363;
    wire N__4358;
    wire N__4355;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4333;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4302;
    wire N__4299;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4291;
    wire N__4286;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4276;
    wire N__4273;
    wire N__4266;
    wire N__4263;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4255;
    wire N__4250;
    wire N__4247;
    wire N__4242;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4219;
    wire N__4216;
    wire N__4213;
    wire N__4210;
    wire N__4203;
    wire N__4200;
    wire N__4197;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4164;
    wire N__4161;
    wire N__4158;
    wire N__4155;
    wire N__4152;
    wire N__4151;
    wire N__4148;
    wire N__4145;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4122;
    wire N__4119;
    wire N__4116;
    wire N__4113;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4101;
    wire N__4098;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4065;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4041;
    wire N__4038;
    wire N__4037;
    wire N__4034;
    wire N__4031;
    wire N__4026;
    wire N__4023;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4011;
    wire N__4008;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__3996;
    wire N__3993;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire N__3981;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3963;
    wire N__3960;
    wire N__3957;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3900;
    wire N__3897;
    wire N__3894;
    wire N__3891;
    wire N__3890;
    wire N__3889;
    wire N__3886;
    wire N__3883;
    wire N__3880;
    wire N__3873;
    wire N__3872;
    wire N__3871;
    wire N__3870;
    wire N__3867;
    wire N__3862;
    wire N__3859;
    wire N__3856;
    wire N__3849;
    wire N__3846;
    wire N__3845;
    wire N__3842;
    wire N__3839;
    wire N__3834;
    wire N__3831;
    wire N__3830;
    wire N__3827;
    wire N__3824;
    wire N__3819;
    wire N__3816;
    wire N__3815;
    wire N__3812;
    wire N__3809;
    wire N__3804;
    wire N__3801;
    wire N__3798;
    wire N__3795;
    wire N__3794;
    wire N__3791;
    wire N__3788;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3776;
    wire N__3773;
    wire N__3770;
    wire N__3765;
    wire N__3762;
    wire N__3759;
    wire N__3756;
    wire N__3753;
    wire N__3750;
    wire N__3747;
    wire N__3744;
    wire N__3743;
    wire N__3742;
    wire N__3741;
    wire N__3740;
    wire N__3739;
    wire N__3738;
    wire N__3727;
    wire N__3722;
    wire N__3717;
    wire N__3714;
    wire N__3713;
    wire N__3712;
    wire N__3709;
    wire N__3706;
    wire N__3705;
    wire N__3704;
    wire N__3703;
    wire N__3700;
    wire N__3699;
    wire N__3696;
    wire N__3691;
    wire N__3688;
    wire N__3681;
    wire N__3672;
    wire N__3671;
    wire N__3670;
    wire N__3667;
    wire N__3666;
    wire N__3665;
    wire N__3664;
    wire N__3663;
    wire N__3658;
    wire N__3647;
    wire N__3642;
    wire N__3639;
    wire N__3636;
    wire N__3635;
    wire N__3634;
    wire N__3633;
    wire N__3632;
    wire N__3631;
    wire N__3630;
    wire N__3621;
    wire N__3614;
    wire N__3609;
    wire N__3606;
    wire N__3605;
    wire N__3600;
    wire N__3597;
    wire N__3594;
    wire N__3591;
    wire N__3590;
    wire N__3589;
    wire N__3588;
    wire N__3587;
    wire N__3586;
    wire N__3585;
    wire N__3584;
    wire N__3581;
    wire N__3578;
    wire N__3569;
    wire N__3562;
    wire N__3555;
    wire N__3552;
    wire N__3551;
    wire N__3550;
    wire N__3549;
    wire N__3548;
    wire N__3547;
    wire N__3544;
    wire N__3537;
    wire N__3532;
    wire N__3525;
    wire N__3524;
    wire N__3523;
    wire N__3522;
    wire N__3513;
    wire N__3510;
    wire N__3507;
    wire N__3504;
    wire N__3501;
    wire N__3498;
    wire N__3495;
    wire N__3494;
    wire N__3491;
    wire N__3488;
    wire N__3483;
    wire N__3480;
    wire N__3477;
    wire N__3474;
    wire N__3471;
    wire N__3468;
    wire N__3467;
    wire N__3462;
    wire N__3459;
    wire N__3458;
    wire N__3457;
    wire N__3456;
    wire N__3453;
    wire N__3448;
    wire N__3445;
    wire N__3438;
    wire N__3437;
    wire N__3436;
    wire N__3435;
    wire N__3430;
    wire N__3425;
    wire N__3420;
    wire N__3419;
    wire N__3416;
    wire N__3415;
    wire N__3412;
    wire N__3411;
    wire N__3406;
    wire N__3401;
    wire N__3396;
    wire N__3393;
    wire N__3390;
    wire N__3387;
    wire N__3384;
    wire N__3381;
    wire N__3378;
    wire N__3375;
    wire N__3374;
    wire N__3373;
    wire N__3370;
    wire N__3369;
    wire N__3368;
    wire N__3361;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3351;
    wire N__3350;
    wire N__3347;
    wire N__3344;
    wire N__3341;
    wire N__3338;
    wire N__3335;
    wire N__3330;
    wire N__3323;
    wire N__3318;
    wire N__3315;
    wire N__3312;
    wire N__3311;
    wire N__3308;
    wire N__3305;
    wire N__3300;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3279;
    wire N__3276;
    wire N__3273;
    wire N__3270;
    wire N__3269;
    wire N__3268;
    wire N__3267;
    wire N__3264;
    wire N__3263;
    wire N__3262;
    wire N__3261;
    wire N__3258;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3244;
    wire N__3241;
    wire N__3238;
    wire N__3233;
    wire N__3228;
    wire N__3225;
    wire N__3224;
    wire N__3219;
    wire N__3214;
    wire N__3211;
    wire N__3204;
    wire N__3201;
    wire N__3198;
    wire N__3195;
    wire N__3192;
    wire N__3191;
    wire N__3188;
    wire N__3185;
    wire N__3180;
    wire N__3177;
    wire N__3174;
    wire N__3171;
    wire N__3168;
    wire N__3165;
    wire N__3162;
    wire N__3159;
    wire N__3156;
    wire N__3155;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3145;
    wire N__3144;
    wire N__3141;
    wire N__3138;
    wire N__3135;
    wire N__3132;
    wire N__3131;
    wire N__3130;
    wire N__3127;
    wire N__3122;
    wire N__3119;
    wire N__3114;
    wire N__3105;
    wire N__3102;
    wire N__3101;
    wire N__3100;
    wire N__3099;
    wire N__3096;
    wire N__3093;
    wire N__3090;
    wire N__3089;
    wire N__3086;
    wire N__3081;
    wire N__3078;
    wire N__3075;
    wire N__3074;
    wire N__3071;
    wire N__3068;
    wire N__3065;
    wire N__3060;
    wire N__3051;
    wire N__3050;
    wire N__3047;
    wire N__3044;
    wire N__3041;
    wire N__3036;
    wire N__3033;
    wire N__3030;
    wire N__3027;
    wire N__3024;
    wire N__3021;
    wire N__3018;
    wire N__3015;
    wire N__3012;
    wire N__3009;
    wire N__3006;
    wire N__3003;
    wire N__3000;
    wire N__2997;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2982;
    wire N__2979;
    wire N__2976;
    wire N__2973;
    wire N__2972;
    wire N__2971;
    wire N__2970;
    wire N__2963;
    wire N__2960;
    wire N__2959;
    wire N__2954;
    wire N__2951;
    wire N__2950;
    wire N__2945;
    wire N__2942;
    wire N__2937;
    wire N__2934;
    wire N__2931;
    wire N__2928;
    wire N__2925;
    wire N__2922;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2912;
    wire N__2907;
    wire N__2904;
    wire N__2901;
    wire N__2900;
    wire N__2895;
    wire N__2892;
    wire N__2889;
    wire N__2888;
    wire N__2885;
    wire N__2880;
    wire N__2877;
    wire N__2874;
    wire N__2871;
    wire N__2868;
    wire N__2865;
    wire N__2862;
    wire N__2861;
    wire N__2856;
    wire N__2853;
    wire N__2850;
    wire N__2847;
    wire N__2844;
    wire N__2841;
    wire N__2840;
    wire N__2835;
    wire N__2832;
    wire N__2829;
    wire N__2826;
    wire N__2823;
    wire N__2822;
    wire N__2817;
    wire N__2814;
    wire N__2811;
    wire N__2808;
    wire N__2805;
    wire N__2802;
    wire N__2801;
    wire N__2798;
    wire N__2795;
    wire N__2792;
    wire N__2789;
    wire N__2784;
    wire N__2781;
    wire N__2778;
    wire N__2775;
    wire N__2774;
    wire N__2771;
    wire N__2768;
    wire N__2763;
    wire N__2760;
    wire N__2757;
    wire N__2754;
    wire N__2751;
    wire N__2750;
    wire N__2745;
    wire N__2742;
    wire N__2739;
    wire N__2736;
    wire N__2733;
    wire N__2730;
    wire N__2727;
    wire N__2726;
    wire N__2723;
    wire N__2720;
    wire N__2717;
    wire N__2714;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2700;
    wire N__2697;
    wire N__2696;
    wire N__2691;
    wire N__2688;
    wire N__2685;
    wire N__2682;
    wire N__2679;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2667;
    wire N__2664;
    wire N__2663;
    wire N__2662;
    wire N__2659;
    wire N__2654;
    wire N__2651;
    wire N__2648;
    wire N__2645;
    wire N__2642;
    wire N__2637;
    wire N__2634;
    wire N__2631;
    wire N__2628;
    wire N__2625;
    wire N__2622;
    wire N__2621;
    wire N__2618;
    wire N__2615;
    wire N__2610;
    wire N__2607;
    wire N__2604;
    wire N__2601;
    wire N__2598;
    wire N__2595;
    wire N__2592;
    wire N__2589;
    wire N__2588;
    wire N__2583;
    wire N__2580;
    wire N__2577;
    wire N__2576;
    wire N__2575;
    wire N__2572;
    wire N__2569;
    wire N__2564;
    wire N__2561;
    wire N__2558;
    wire N__2557;
    wire N__2552;
    wire N__2549;
    wire N__2544;
    wire N__2541;
    wire N__2540;
    wire N__2539;
    wire N__2538;
    wire N__2537;
    wire N__2536;
    wire N__2535;
    wire N__2534;
    wire N__2533;
    wire N__2532;
    wire N__2531;
    wire N__2530;
    wire N__2505;
    wire CLK80_OUT;
    wire GNDG0;
    wire VCCG0;
    wire A_c_18;
    wire A_c_16;
    wire A_c_17;
    wire \U409_CIA.g0Z0Z_11_cascade_ ;
    wire \U409_CIA.g0Z0Z_8 ;
    wire A_c_19;
    wire \U409_ADDRESS_DECODE.ROMEN_0_a2_0Z0Z_2_cascade_ ;
    wire \U409_ADDRESS_DECODE.N_58 ;
    wire OVL_c;
    wire \U409_ADDRESS_DECODE.CIA_SPACEm_6 ;
    wire A_c_20;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ;
    wire \U409_ADDRESS_DECODE.un1_nREGSPACEZ0_cascade_ ;
    wire PORTSIZE_0_i;
    wire A_c_22;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ;
    wire \U409_CIA.g0Z0Z_2_cascade_ ;
    wire \U409_CIA.g0Z0Z_10 ;
    wire A_c_27;
    wire A_c_25;
    wire A_c_26;
    wire A_c_24;
    wire A_c_31;
    wire A_c_29;
    wire A_c_30;
    wire A_c_28;
    wire U409_ADDRESS_DECODE_un1_nRAMSPACE_i;
    wire A_c_21;
    wire \U409_ADDRESS_DECODE.un1_nRAMSPACEZ0Z_2 ;
    wire \U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ;
    wire nBUFEN_c;
    wire A_c_23;
    wire \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ;
    wire U409_ADDRESS_DECODE_un1_nREGSPACE_i;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ;
    wire \U409_ADDRESS_DECODE.N_23 ;
    wire ROMENm_i;
    wire bfn_7_6_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ;
    wire \U409_CIA.CIA_CLK_COUNT11_0_a2_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.N_9_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.N_20_cascade_ ;
    wire \U409_CIA.CLKCIA8_0_a2_0 ;
    wire \U409_CIA.CLKCIA6_0_a2_1 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CLKCIAZ0_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire CLK28_IN_c_g;
    wire TICK60_c;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire \U409_TICK.TICK603_10_cascade_ ;
    wire \U409_TICK.TICK603_8_cascade_ ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.TICK603_11 ;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_nCIACS1_i;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_nCIACS0_i;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire bfn_9_7_0_;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire bfn_9_8_0_;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire ROMENm;
    wire \U409_TRANSFER_ACK.N_24_cascade_ ;
    wire \U409_TRANSFER_ACK.N_22 ;
    wire bfn_10_5_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire bfn_10_6_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire CIA_ENABLEm;
    wire \U409_CIA.g0Z0Z_14 ;
    wire \U409_CIA.g0Z0Z_13 ;
    wire \U409_CIA.VMAZ0 ;
    wire \U409_CIA.CIA_HOLDZ0 ;
    wire CLKCIA_c;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_EN_nesrC_net ;
    wire \U409_TRANSFER_ACK.N_22_0_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_24 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire TICK50_c;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire \U409_TICK.TICK503_11 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire CLK6_c_g;
    wire \U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_49 ;
    wire \U409_TRANSFER_ACK.N_29_cascade_ ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_1C_net ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_53 ;
    wire \U409_TRANSFER_ACK.N_52_cascade_ ;
    wire \U409_TRANSFER_ACK.N_29 ;
    wire \U409_TRANSFER_ACK.m9_i_1_cascade_ ;
    wire \U409_TRANSFER_ACK.N_54 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire \U409_TRANSFER_ACK.N_60 ;
    wire \U409_TRANSFER_ACK.N_55 ;
    wire \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ;
    wire RESETn_c_i;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_ ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire TACK_OUTn;
    wire \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ;
    wire \INVU409_TRANSFER_ACK.TACK_EN_iC_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ;
    wire CONSTANT_ONE_NET;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.N_41 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_4_cascade_ ;
    wire TSn_c;
    wire \U409_TRANSFER_ACK.N_41_4_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a4_0_2_0_cascade_ ;
    wire CLK40_IN_c;
    wire \U409_TRANSFER_ACK.N_44_cascade_ ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0_cascade_ ;
    wire \U409_TRANSFER_ACK.N_41_4 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_41_i ;
    wire bfn_14_14_0_;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_THRU_CO ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2_THRU_CO ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3_THRU_CO ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4_THRU_CO ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5_THRU_CO ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5 ;
    wire \U409_TRANSFER_ACK.N_35 ;
    wire \U409_TRANSFER_ACK.N_44 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ;
    wire TACKn_in;
    wire RESETn_c;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire TACK_EN_i;
    wire N_391_i;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__5445),
            .RESETB(N__5250),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6365),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__6367),
            .DIN(N__6366),
            .DOUT(N__6365),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__6367),
            .PADOUT(N__6366),
            .PADIN(N__6365),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6355),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__6357),
            .DIN(N__6356),
            .DOUT(N__6355),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__6357),
            .PADOUT(N__6356),
            .PADIN(N__6355),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKCIA_obuf_iopad (
            .OE(N__6346),
            .DIN(N__6345),
            .DOUT(N__6344),
            .PACKAGEPIN(CLKCIA));
    defparam CLKCIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKCIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKCIA_obuf_preio (
            .PADOEN(N__6346),
            .PADOUT(N__6345),
            .PADIN(N__6344),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4242),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_24_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_24_iopad (
            .OE(N__6337),
            .DIN(N__6336),
            .DOUT(N__6335),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__6337),
            .PADOUT(N__6336),
            .PADIN(N__6335),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nCIACS0_obuf_iopad (
            .OE(N__6328),
            .DIN(N__6327),
            .DOUT(N__6326),
            .PACKAGEPIN(nCIACS0));
    defparam nCIACS0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCIACS0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCIACS0_obuf_preio (
            .PADOEN(N__6328),
            .PADOUT(N__6327),
            .PADIN(N__6326),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3912),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nCIACS1_obuf_iopad (
            .OE(N__6319),
            .DIN(N__6318),
            .DOUT(N__6317),
            .PACKAGEPIN(nCIACS1));
    defparam nCIACS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCIACS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCIACS1_obuf_preio (
            .PADOEN(N__6319),
            .PADOUT(N__6318),
            .PADIN(N__6317),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3948),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_31_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_31_iopad (
            .OE(N__6310),
            .DIN(N__6309),
            .DOUT(N__6308),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__6310),
            .PADOUT(N__6309),
            .PADIN(N__6308),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_17_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_17_iopad (
            .OE(N__6301),
            .DIN(N__6300),
            .DOUT(N__6299),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__6301),
            .PADOUT(N__6300),
            .PADIN(N__6299),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_21_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_21_iopad (
            .OE(N__6292),
            .DIN(N__6291),
            .DOUT(N__6290),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__6292),
            .PADOUT(N__6291),
            .PADIN(N__6290),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TACKn_iobuf_iopad.PULLUP=1'b1;
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__6283),
            .DIN(N__6282),
            .DOUT(N__6281),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__6283),
            .PADOUT(N__6282),
            .PADIN(N__6281),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5700),
            .DIN0(TACKn_in),
            .DOUT0(N__5301),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_12_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_12_iopad (
            .OE(N__6274),
            .DIN(N__6273),
            .DOUT(N__6272),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__6274),
            .PADOUT(N__6273),
            .PADIN(N__6272),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__6265),
            .DIN(N__6264),
            .DOUT(N__6263),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__6265),
            .PADOUT(N__6264),
            .PADIN(N__6263),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PORTSIZE_obuf_iopad.PULLUP=1'b1;
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__6256),
            .DIN(N__6255),
            .DOUT(N__6254),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__6256),
            .PADOUT(N__6255),
            .PADIN(N__6254),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2991),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nRAMSPACE_obuf_iopad (
            .OE(N__6247),
            .DIN(N__6246),
            .DOUT(N__6245),
            .PACKAGEPIN(nRAMSPACE));
    defparam nRAMSPACE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nRAMSPACE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nRAMSPACE_obuf_preio (
            .PADOEN(N__6247),
            .PADOUT(N__6246),
            .PADIN(N__6245),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3396),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nROMEN_obuf_iopad (
            .OE(N__6238),
            .DIN(N__6237),
            .DOUT(N__6236),
            .PACKAGEPIN(nROMEN));
    defparam nROMEN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nROMEN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nROMEN_obuf_preio (
            .PADOEN(N__6238),
            .PADOUT(N__6237),
            .PADIN(N__6236),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3030),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_18_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_18_iopad (
            .OE(N__6229),
            .DIN(N__6228),
            .DOUT(N__6227),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__6229),
            .PADOUT(N__6228),
            .PADIN(N__6227),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_29_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_29_iopad (
            .OE(N__6220),
            .DIN(N__6219),
            .DOUT(N__6218),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__6220),
            .PADOUT(N__6219),
            .PADIN(N__6218),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nBUFEN_obuf_iopad (
            .OE(N__6211),
            .DIN(N__6210),
            .DOUT(N__6209),
            .PACKAGEPIN(nBUFEN));
    defparam nBUFEN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nBUFEN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nBUFEN_obuf_preio (
            .PADOEN(N__6211),
            .PADOUT(N__6210),
            .PADIN(N__6209),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3294),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_22_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_22_iopad (
            .OE(N__6202),
            .DIN(N__6201),
            .DOUT(N__6200),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__6202),
            .PADOUT(N__6201),
            .PADIN(N__6200),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_27_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_27_iopad (
            .OE(N__6193),
            .DIN(N__6192),
            .DOUT(N__6191),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__6193),
            .PADOUT(N__6192),
            .PADIN(N__6191),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__6184),
            .DIN(N__6183),
            .DOUT(N__6182),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__6184),
            .PADOUT(N__6183),
            .PADIN(N__6182),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__6175),
            .DIN(N__6174),
            .DOUT(N__6173),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__6175),
            .PADOUT(N__6174),
            .PADIN(N__6173),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_20_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_20_iopad (
            .OE(N__6166),
            .DIN(N__6165),
            .DOUT(N__6164),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__6166),
            .PADOUT(N__6165),
            .PADIN(N__6164),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_13_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_13_iopad (
            .OE(N__6157),
            .DIN(N__6156),
            .DOUT(N__6155),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__6157),
            .PADOUT(N__6156),
            .PADIN(N__6155),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_25_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_25_iopad (
            .OE(N__6148),
            .DIN(N__6147),
            .DOUT(N__6146),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__6148),
            .PADOUT(N__6147),
            .PADIN(N__6146),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD nREGSPACE_obuf_iopad (
            .OE(N__6139),
            .DIN(N__6138),
            .DOUT(N__6137),
            .PACKAGEPIN(nREGSPACE));
    defparam nREGSPACE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nREGSPACE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nREGSPACE_obuf_preio (
            .PADOEN(N__6139),
            .PADOUT(N__6138),
            .PADIN(N__6137),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3180),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__6130),
            .DIN(N__6129),
            .DOUT(N__6128),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__6130),
            .PADOUT(N__6129),
            .PADIN(N__6128),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4710),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_19_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_19_iopad (
            .OE(N__6121),
            .DIN(N__6120),
            .DOUT(N__6119),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__6121),
            .PADOUT(N__6120),
            .PADIN(N__6119),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_28_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_28_iopad (
            .OE(N__6112),
            .DIN(N__6111),
            .DOUT(N__6110),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__6112),
            .PADOUT(N__6111),
            .PADIN(N__6110),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_30_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_30_iopad (
            .OE(N__6103),
            .DIN(N__6102),
            .DOUT(N__6101),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__6103),
            .PADOUT(N__6102),
            .PADIN(N__6101),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__6094),
            .DIN(N__6093),
            .DOUT(N__6092),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__6094),
            .PADOUT(N__6093),
            .PADIN(N__6092),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_16_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_16_iopad (
            .OE(N__6085),
            .DIN(N__6084),
            .DOUT(N__6083),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__6085),
            .PADOUT(N__6084),
            .PADIN(N__6083),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__6076),
            .DIN(N__6075),
            .DOUT(N__6074),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__6076),
            .PADOUT(N__6075),
            .PADIN(N__6074),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3507),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_26_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_26_iopad (
            .OE(N__6067),
            .DIN(N__6066),
            .DOUT(N__6065),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__6067),
            .PADOUT(N__6066),
            .PADIN(N__6065),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_23_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_23_iopad (
            .OE(N__6058),
            .DIN(N__6057),
            .DOUT(N__6056),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__6058),
            .PADOUT(N__6057),
            .PADIN(N__6056),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__1397 (
            .O(N__6039),
            .I(N__6036));
    InMux I__1396 (
            .O(N__6036),
            .I(N__6030));
    InMux I__1395 (
            .O(N__6035),
            .I(N__6027));
    InMux I__1394 (
            .O(N__6034),
            .I(N__6024));
    InMux I__1393 (
            .O(N__6033),
            .I(N__6021));
    LocalMux I__1392 (
            .O(N__6030),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__1391 (
            .O(N__6027),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__1390 (
            .O(N__6024),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__1389 (
            .O(N__6021),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    InMux I__1388 (
            .O(N__6012),
            .I(N__6009));
    LocalMux I__1387 (
            .O(N__6009),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5_THRU_CO ));
    InMux I__1386 (
            .O(N__6006),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5 ));
    CascadeMux I__1385 (
            .O(N__6003),
            .I(N__5994));
    InMux I__1384 (
            .O(N__6002),
            .I(N__5990));
    InMux I__1383 (
            .O(N__6001),
            .I(N__5987));
    InMux I__1382 (
            .O(N__6000),
            .I(N__5982));
    InMux I__1381 (
            .O(N__5999),
            .I(N__5982));
    InMux I__1380 (
            .O(N__5998),
            .I(N__5975));
    InMux I__1379 (
            .O(N__5997),
            .I(N__5975));
    InMux I__1378 (
            .O(N__5994),
            .I(N__5975));
    InMux I__1377 (
            .O(N__5993),
            .I(N__5972));
    LocalMux I__1376 (
            .O(N__5990),
            .I(\U409_TRANSFER_ACK.N_35 ));
    LocalMux I__1375 (
            .O(N__5987),
            .I(\U409_TRANSFER_ACK.N_35 ));
    LocalMux I__1374 (
            .O(N__5982),
            .I(\U409_TRANSFER_ACK.N_35 ));
    LocalMux I__1373 (
            .O(N__5975),
            .I(\U409_TRANSFER_ACK.N_35 ));
    LocalMux I__1372 (
            .O(N__5972),
            .I(\U409_TRANSFER_ACK.N_35 ));
    CascadeMux I__1371 (
            .O(N__5961),
            .I(N__5957));
    CascadeMux I__1370 (
            .O(N__5960),
            .I(N__5952));
    InMux I__1369 (
            .O(N__5957),
            .I(N__5945));
    InMux I__1368 (
            .O(N__5956),
            .I(N__5945));
    InMux I__1367 (
            .O(N__5955),
            .I(N__5938));
    InMux I__1366 (
            .O(N__5952),
            .I(N__5938));
    InMux I__1365 (
            .O(N__5951),
            .I(N__5938));
    InMux I__1364 (
            .O(N__5950),
            .I(N__5935));
    LocalMux I__1363 (
            .O(N__5945),
            .I(\U409_TRANSFER_ACK.N_44 ));
    LocalMux I__1362 (
            .O(N__5938),
            .I(\U409_TRANSFER_ACK.N_44 ));
    LocalMux I__1361 (
            .O(N__5935),
            .I(\U409_TRANSFER_ACK.N_44 ));
    InMux I__1360 (
            .O(N__5928),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_6 ));
    CascadeMux I__1359 (
            .O(N__5925),
            .I(N__5920));
    CascadeMux I__1358 (
            .O(N__5924),
            .I(N__5917));
    InMux I__1357 (
            .O(N__5923),
            .I(N__5914));
    InMux I__1356 (
            .O(N__5920),
            .I(N__5911));
    InMux I__1355 (
            .O(N__5917),
            .I(N__5908));
    LocalMux I__1354 (
            .O(N__5914),
            .I(N__5905));
    LocalMux I__1353 (
            .O(N__5911),
            .I(N__5900));
    LocalMux I__1352 (
            .O(N__5908),
            .I(N__5900));
    Odrv4 I__1351 (
            .O(N__5905),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    Odrv4 I__1350 (
            .O(N__5900),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    InMux I__1349 (
            .O(N__5895),
            .I(N__5892));
    LocalMux I__1348 (
            .O(N__5892),
            .I(N__5889));
    Span4Mux_v I__1347 (
            .O(N__5889),
            .I(N__5886));
    Sp12to4 I__1346 (
            .O(N__5886),
            .I(N__5883));
    Span12Mux_h I__1345 (
            .O(N__5883),
            .I(N__5880));
    Span12Mux_v I__1344 (
            .O(N__5880),
            .I(N__5877));
    Odrv12 I__1343 (
            .O(N__5877),
            .I(TACKn_in));
    InMux I__1342 (
            .O(N__5874),
            .I(N__5870));
    CascadeMux I__1341 (
            .O(N__5873),
            .I(N__5867));
    LocalMux I__1340 (
            .O(N__5870),
            .I(N__5862));
    InMux I__1339 (
            .O(N__5867),
            .I(N__5859));
    InMux I__1338 (
            .O(N__5866),
            .I(N__5856));
    CascadeMux I__1337 (
            .O(N__5865),
            .I(N__5852));
    Span4Mux_v I__1336 (
            .O(N__5862),
            .I(N__5849));
    LocalMux I__1335 (
            .O(N__5859),
            .I(N__5846));
    LocalMux I__1334 (
            .O(N__5856),
            .I(N__5843));
    InMux I__1333 (
            .O(N__5855),
            .I(N__5835));
    InMux I__1332 (
            .O(N__5852),
            .I(N__5829));
    Span4Mux_h I__1331 (
            .O(N__5849),
            .I(N__5824));
    Span4Mux_v I__1330 (
            .O(N__5846),
            .I(N__5824));
    Span4Mux_h I__1329 (
            .O(N__5843),
            .I(N__5821));
    InMux I__1328 (
            .O(N__5842),
            .I(N__5818));
    InMux I__1327 (
            .O(N__5841),
            .I(N__5809));
    InMux I__1326 (
            .O(N__5840),
            .I(N__5809));
    InMux I__1325 (
            .O(N__5839),
            .I(N__5809));
    InMux I__1324 (
            .O(N__5838),
            .I(N__5809));
    LocalMux I__1323 (
            .O(N__5835),
            .I(N__5806));
    InMux I__1322 (
            .O(N__5834),
            .I(N__5803));
    InMux I__1321 (
            .O(N__5833),
            .I(N__5800));
    InMux I__1320 (
            .O(N__5832),
            .I(N__5797));
    LocalMux I__1319 (
            .O(N__5829),
            .I(N__5792));
    Sp12to4 I__1318 (
            .O(N__5824),
            .I(N__5792));
    Span4Mux_h I__1317 (
            .O(N__5821),
            .I(N__5785));
    LocalMux I__1316 (
            .O(N__5818),
            .I(N__5785));
    LocalMux I__1315 (
            .O(N__5809),
            .I(N__5785));
    Span4Mux_h I__1314 (
            .O(N__5806),
            .I(N__5778));
    LocalMux I__1313 (
            .O(N__5803),
            .I(N__5778));
    LocalMux I__1312 (
            .O(N__5800),
            .I(N__5778));
    LocalMux I__1311 (
            .O(N__5797),
            .I(N__5775));
    Span12Mux_h I__1310 (
            .O(N__5792),
            .I(N__5768));
    Sp12to4 I__1309 (
            .O(N__5785),
            .I(N__5768));
    Sp12to4 I__1308 (
            .O(N__5778),
            .I(N__5768));
    Span12Mux_h I__1307 (
            .O(N__5775),
            .I(N__5765));
    Span12Mux_v I__1306 (
            .O(N__5768),
            .I(N__5762));
    Span12Mux_v I__1305 (
            .O(N__5765),
            .I(N__5757));
    Span12Mux_h I__1304 (
            .O(N__5762),
            .I(N__5757));
    Odrv12 I__1303 (
            .O(N__5757),
            .I(RESETn_c));
    SRMux I__1302 (
            .O(N__5754),
            .I(N__5751));
    LocalMux I__1301 (
            .O(N__5751),
            .I(N__5746));
    SRMux I__1300 (
            .O(N__5750),
            .I(N__5742));
    SRMux I__1299 (
            .O(N__5749),
            .I(N__5739));
    Span4Mux_v I__1298 (
            .O(N__5746),
            .I(N__5736));
    SRMux I__1297 (
            .O(N__5745),
            .I(N__5733));
    LocalMux I__1296 (
            .O(N__5742),
            .I(N__5730));
    LocalMux I__1295 (
            .O(N__5739),
            .I(N__5727));
    Odrv4 I__1294 (
            .O(N__5736),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    LocalMux I__1293 (
            .O(N__5733),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv12 I__1292 (
            .O(N__5730),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv4 I__1291 (
            .O(N__5727),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__1290 (
            .O(N__5718),
            .I(N__5715));
    LocalMux I__1289 (
            .O(N__5715),
            .I(N__5712));
    Span4Mux_v I__1288 (
            .O(N__5712),
            .I(N__5709));
    Span4Mux_h I__1287 (
            .O(N__5709),
            .I(N__5706));
    Span4Mux_v I__1286 (
            .O(N__5706),
            .I(N__5703));
    Odrv4 I__1285 (
            .O(N__5703),
            .I(TACK_EN_i));
    IoInMux I__1284 (
            .O(N__5700),
            .I(N__5697));
    LocalMux I__1283 (
            .O(N__5697),
            .I(N__5694));
    Span4Mux_s3_v I__1282 (
            .O(N__5694),
            .I(N__5691));
    Span4Mux_v I__1281 (
            .O(N__5691),
            .I(N__5688));
    Sp12to4 I__1280 (
            .O(N__5688),
            .I(N__5685));
    Odrv12 I__1279 (
            .O(N__5685),
            .I(N_391_i));
    InMux I__1278 (
            .O(N__5682),
            .I(N__5677));
    InMux I__1277 (
            .O(N__5681),
            .I(N__5672));
    InMux I__1276 (
            .O(N__5680),
            .I(N__5672));
    LocalMux I__1275 (
            .O(N__5677),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1274 (
            .O(N__5672),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    CascadeMux I__1273 (
            .O(N__5667),
            .I(N__5663));
    InMux I__1272 (
            .O(N__5666),
            .I(N__5660));
    InMux I__1271 (
            .O(N__5663),
            .I(N__5657));
    LocalMux I__1270 (
            .O(N__5660),
            .I(\U409_TRANSFER_ACK.N_41_i ));
    LocalMux I__1269 (
            .O(N__5657),
            .I(\U409_TRANSFER_ACK.N_41_i ));
    InMux I__1268 (
            .O(N__5652),
            .I(N__5646));
    InMux I__1267 (
            .O(N__5651),
            .I(N__5643));
    InMux I__1266 (
            .O(N__5650),
            .I(N__5638));
    InMux I__1265 (
            .O(N__5649),
            .I(N__5638));
    LocalMux I__1264 (
            .O(N__5646),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1263 (
            .O(N__5643),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1262 (
            .O(N__5638),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    CascadeMux I__1261 (
            .O(N__5631),
            .I(N__5628));
    InMux I__1260 (
            .O(N__5628),
            .I(N__5625));
    LocalMux I__1259 (
            .O(N__5625),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_THRU_CO ));
    InMux I__1258 (
            .O(N__5622),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0 ));
    CascadeMux I__1257 (
            .O(N__5619),
            .I(N__5614));
    InMux I__1256 (
            .O(N__5618),
            .I(N__5609));
    InMux I__1255 (
            .O(N__5617),
            .I(N__5606));
    InMux I__1254 (
            .O(N__5614),
            .I(N__5603));
    InMux I__1253 (
            .O(N__5613),
            .I(N__5600));
    InMux I__1252 (
            .O(N__5612),
            .I(N__5597));
    LocalMux I__1251 (
            .O(N__5609),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1250 (
            .O(N__5606),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1249 (
            .O(N__5603),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1248 (
            .O(N__5600),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1247 (
            .O(N__5597),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    InMux I__1246 (
            .O(N__5586),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_1 ));
    InMux I__1245 (
            .O(N__5583),
            .I(N__5577));
    InMux I__1244 (
            .O(N__5582),
            .I(N__5574));
    InMux I__1243 (
            .O(N__5581),
            .I(N__5569));
    InMux I__1242 (
            .O(N__5580),
            .I(N__5569));
    LocalMux I__1241 (
            .O(N__5577),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1240 (
            .O(N__5574),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1239 (
            .O(N__5569),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    InMux I__1238 (
            .O(N__5562),
            .I(N__5559));
    LocalMux I__1237 (
            .O(N__5559),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2_THRU_CO ));
    InMux I__1236 (
            .O(N__5556),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2 ));
    InMux I__1235 (
            .O(N__5553),
            .I(N__5547));
    InMux I__1234 (
            .O(N__5552),
            .I(N__5544));
    InMux I__1233 (
            .O(N__5551),
            .I(N__5541));
    InMux I__1232 (
            .O(N__5550),
            .I(N__5538));
    LocalMux I__1231 (
            .O(N__5547),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1230 (
            .O(N__5544),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1229 (
            .O(N__5541),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1228 (
            .O(N__5538),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    InMux I__1227 (
            .O(N__5529),
            .I(N__5526));
    LocalMux I__1226 (
            .O(N__5526),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3_THRU_CO ));
    InMux I__1225 (
            .O(N__5523),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3 ));
    CascadeMux I__1224 (
            .O(N__5520),
            .I(N__5517));
    InMux I__1223 (
            .O(N__5517),
            .I(N__5509));
    InMux I__1222 (
            .O(N__5516),
            .I(N__5504));
    InMux I__1221 (
            .O(N__5515),
            .I(N__5504));
    InMux I__1220 (
            .O(N__5514),
            .I(N__5499));
    InMux I__1219 (
            .O(N__5513),
            .I(N__5499));
    InMux I__1218 (
            .O(N__5512),
            .I(N__5496));
    LocalMux I__1217 (
            .O(N__5509),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__1216 (
            .O(N__5504),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__1215 (
            .O(N__5499),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__1214 (
            .O(N__5496),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    InMux I__1213 (
            .O(N__5487),
            .I(N__5484));
    LocalMux I__1212 (
            .O(N__5484),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4_THRU_CO ));
    InMux I__1211 (
            .O(N__5481),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4 ));
    InMux I__1210 (
            .O(N__5478),
            .I(N__5475));
    LocalMux I__1209 (
            .O(N__5475),
            .I(N__5472));
    Span4Mux_v I__1208 (
            .O(N__5472),
            .I(N__5468));
    InMux I__1207 (
            .O(N__5471),
            .I(N__5465));
    Sp12to4 I__1206 (
            .O(N__5468),
            .I(N__5460));
    LocalMux I__1205 (
            .O(N__5465),
            .I(N__5460));
    Span12Mux_h I__1204 (
            .O(N__5460),
            .I(N__5457));
    Span12Mux_v I__1203 (
            .O(N__5457),
            .I(N__5454));
    Odrv12 I__1202 (
            .O(N__5454),
            .I(TSn_c));
    CascadeMux I__1201 (
            .O(N__5451),
            .I(\U409_TRANSFER_ACK.N_41_4_cascade_ ));
    CascadeMux I__1200 (
            .O(N__5448),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a4_0_2_0_cascade_ ));
    IoInMux I__1199 (
            .O(N__5445),
            .I(N__5442));
    LocalMux I__1198 (
            .O(N__5442),
            .I(N__5438));
    InMux I__1197 (
            .O(N__5441),
            .I(N__5434));
    IoSpan4Mux I__1196 (
            .O(N__5438),
            .I(N__5429));
    InMux I__1195 (
            .O(N__5437),
            .I(N__5426));
    LocalMux I__1194 (
            .O(N__5434),
            .I(N__5423));
    InMux I__1193 (
            .O(N__5433),
            .I(N__5420));
    InMux I__1192 (
            .O(N__5432),
            .I(N__5417));
    Span4Mux_s0_v I__1191 (
            .O(N__5429),
            .I(N__5414));
    LocalMux I__1190 (
            .O(N__5426),
            .I(N__5411));
    Span4Mux_h I__1189 (
            .O(N__5423),
            .I(N__5406));
    LocalMux I__1188 (
            .O(N__5420),
            .I(N__5406));
    LocalMux I__1187 (
            .O(N__5417),
            .I(N__5403));
    Sp12to4 I__1186 (
            .O(N__5414),
            .I(N__5400));
    Span4Mux_v I__1185 (
            .O(N__5411),
            .I(N__5397));
    Span4Mux_v I__1184 (
            .O(N__5406),
            .I(N__5392));
    Span4Mux_h I__1183 (
            .O(N__5403),
            .I(N__5392));
    Span12Mux_v I__1182 (
            .O(N__5400),
            .I(N__5389));
    Sp12to4 I__1181 (
            .O(N__5397),
            .I(N__5386));
    Sp12to4 I__1180 (
            .O(N__5392),
            .I(N__5383));
    Span12Mux_v I__1179 (
            .O(N__5389),
            .I(N__5380));
    Span12Mux_h I__1178 (
            .O(N__5386),
            .I(N__5377));
    Span12Mux_v I__1177 (
            .O(N__5383),
            .I(N__5374));
    Odrv12 I__1176 (
            .O(N__5380),
            .I(CLK40_IN_c));
    Odrv12 I__1175 (
            .O(N__5377),
            .I(CLK40_IN_c));
    Odrv12 I__1174 (
            .O(N__5374),
            .I(CLK40_IN_c));
    CascadeMux I__1173 (
            .O(N__5367),
            .I(\U409_TRANSFER_ACK.N_44_cascade_ ));
    CascadeMux I__1172 (
            .O(N__5364),
            .I(N__5360));
    InMux I__1171 (
            .O(N__5363),
            .I(N__5357));
    InMux I__1170 (
            .O(N__5360),
            .I(N__5354));
    LocalMux I__1169 (
            .O(N__5357),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0 ));
    LocalMux I__1168 (
            .O(N__5354),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0 ));
    CascadeMux I__1167 (
            .O(N__5349),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0_cascade_ ));
    InMux I__1166 (
            .O(N__5346),
            .I(N__5342));
    InMux I__1165 (
            .O(N__5345),
            .I(N__5339));
    LocalMux I__1164 (
            .O(N__5342),
            .I(\U409_TRANSFER_ACK.N_41_4 ));
    LocalMux I__1163 (
            .O(N__5339),
            .I(\U409_TRANSFER_ACK.N_41_4 ));
    CascadeMux I__1162 (
            .O(N__5334),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ));
    InMux I__1161 (
            .O(N__5331),
            .I(N__5322));
    InMux I__1160 (
            .O(N__5330),
            .I(N__5322));
    InMux I__1159 (
            .O(N__5329),
            .I(N__5322));
    LocalMux I__1158 (
            .O(N__5322),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    CascadeMux I__1157 (
            .O(N__5319),
            .I(N__5316));
    InMux I__1156 (
            .O(N__5316),
            .I(N__5311));
    InMux I__1155 (
            .O(N__5315),
            .I(N__5306));
    InMux I__1154 (
            .O(N__5314),
            .I(N__5306));
    LocalMux I__1153 (
            .O(N__5311),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__1152 (
            .O(N__5306),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    IoInMux I__1151 (
            .O(N__5301),
            .I(N__5298));
    LocalMux I__1150 (
            .O(N__5298),
            .I(N__5295));
    IoSpan4Mux I__1149 (
            .O(N__5295),
            .I(N__5292));
    Span4Mux_s2_v I__1148 (
            .O(N__5292),
            .I(N__5289));
    Sp12to4 I__1147 (
            .O(N__5289),
            .I(N__5286));
    Span12Mux_v I__1146 (
            .O(N__5286),
            .I(N__5282));
    InMux I__1145 (
            .O(N__5285),
            .I(N__5279));
    Odrv12 I__1144 (
            .O(N__5282),
            .I(TACK_OUTn));
    LocalMux I__1143 (
            .O(N__5279),
            .I(TACK_OUTn));
    InMux I__1142 (
            .O(N__5274),
            .I(N__5270));
    InMux I__1141 (
            .O(N__5273),
            .I(N__5267));
    LocalMux I__1140 (
            .O(N__5270),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ));
    LocalMux I__1139 (
            .O(N__5267),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ));
    CEMux I__1138 (
            .O(N__5262),
            .I(N__5259));
    LocalMux I__1137 (
            .O(N__5259),
            .I(N__5256));
    Span4Mux_v I__1136 (
            .O(N__5256),
            .I(N__5253));
    Odrv4 I__1135 (
            .O(N__5253),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ));
    IoInMux I__1134 (
            .O(N__5250),
            .I(N__5247));
    LocalMux I__1133 (
            .O(N__5247),
            .I(N__5244));
    Span4Mux_s3_v I__1132 (
            .O(N__5244),
            .I(N__5241));
    Span4Mux_h I__1131 (
            .O(N__5241),
            .I(N__5238));
    Odrv4 I__1130 (
            .O(N__5238),
            .I(CONSTANT_ONE_NET));
    InMux I__1129 (
            .O(N__5235),
            .I(N__5231));
    InMux I__1128 (
            .O(N__5234),
            .I(N__5228));
    LocalMux I__1127 (
            .O(N__5231),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    LocalMux I__1126 (
            .O(N__5228),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    InMux I__1125 (
            .O(N__5223),
            .I(N__5220));
    LocalMux I__1124 (
            .O(N__5220),
            .I(\U409_TRANSFER_ACK.N_41 ));
    CascadeMux I__1123 (
            .O(N__5217),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_4_cascade_ ));
    InMux I__1122 (
            .O(N__5214),
            .I(N__5207));
    InMux I__1121 (
            .O(N__5213),
            .I(N__5204));
    InMux I__1120 (
            .O(N__5212),
            .I(N__5201));
    InMux I__1119 (
            .O(N__5211),
            .I(N__5196));
    InMux I__1118 (
            .O(N__5210),
            .I(N__5196));
    LocalMux I__1117 (
            .O(N__5207),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__1116 (
            .O(N__5204),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__1115 (
            .O(N__5201),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__1114 (
            .O(N__5196),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    CascadeMux I__1113 (
            .O(N__5187),
            .I(N__5180));
    InMux I__1112 (
            .O(N__5186),
            .I(N__5172));
    InMux I__1111 (
            .O(N__5185),
            .I(N__5172));
    InMux I__1110 (
            .O(N__5184),
            .I(N__5172));
    InMux I__1109 (
            .O(N__5183),
            .I(N__5165));
    InMux I__1108 (
            .O(N__5180),
            .I(N__5165));
    InMux I__1107 (
            .O(N__5179),
            .I(N__5165));
    LocalMux I__1106 (
            .O(N__5172),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__1105 (
            .O(N__5165),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    InMux I__1104 (
            .O(N__5160),
            .I(N__5154));
    CascadeMux I__1103 (
            .O(N__5159),
            .I(N__5151));
    CascadeMux I__1102 (
            .O(N__5158),
            .I(N__5148));
    CascadeMux I__1101 (
            .O(N__5157),
            .I(N__5145));
    LocalMux I__1100 (
            .O(N__5154),
            .I(N__5142));
    InMux I__1099 (
            .O(N__5151),
            .I(N__5139));
    InMux I__1098 (
            .O(N__5148),
            .I(N__5134));
    InMux I__1097 (
            .O(N__5145),
            .I(N__5134));
    Odrv4 I__1096 (
            .O(N__5142),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    LocalMux I__1095 (
            .O(N__5139),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    LocalMux I__1094 (
            .O(N__5134),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    InMux I__1093 (
            .O(N__5127),
            .I(N__5124));
    LocalMux I__1092 (
            .O(N__5124),
            .I(\U409_TRANSFER_ACK.N_53 ));
    CascadeMux I__1091 (
            .O(N__5121),
            .I(\U409_TRANSFER_ACK.N_52_cascade_ ));
    InMux I__1090 (
            .O(N__5118),
            .I(N__5115));
    LocalMux I__1089 (
            .O(N__5115),
            .I(\U409_TRANSFER_ACK.N_29 ));
    CascadeMux I__1088 (
            .O(N__5112),
            .I(\U409_TRANSFER_ACK.m9_i_1_cascade_ ));
    InMux I__1087 (
            .O(N__5109),
            .I(N__5106));
    LocalMux I__1086 (
            .O(N__5106),
            .I(\U409_TRANSFER_ACK.N_54 ));
    InMux I__1085 (
            .O(N__5103),
            .I(N__5094));
    InMux I__1084 (
            .O(N__5102),
            .I(N__5094));
    InMux I__1083 (
            .O(N__5101),
            .I(N__5087));
    InMux I__1082 (
            .O(N__5100),
            .I(N__5087));
    InMux I__1081 (
            .O(N__5099),
            .I(N__5087));
    LocalMux I__1080 (
            .O(N__5094),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1079 (
            .O(N__5087),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    InMux I__1078 (
            .O(N__5082),
            .I(N__5079));
    LocalMux I__1077 (
            .O(N__5079),
            .I(N__5074));
    InMux I__1076 (
            .O(N__5078),
            .I(N__5071));
    InMux I__1075 (
            .O(N__5077),
            .I(N__5068));
    Odrv4 I__1074 (
            .O(N__5074),
            .I(\U409_TRANSFER_ACK.N_60 ));
    LocalMux I__1073 (
            .O(N__5071),
            .I(\U409_TRANSFER_ACK.N_60 ));
    LocalMux I__1072 (
            .O(N__5068),
            .I(\U409_TRANSFER_ACK.N_60 ));
    InMux I__1071 (
            .O(N__5061),
            .I(N__5058));
    LocalMux I__1070 (
            .O(N__5058),
            .I(\U409_TRANSFER_ACK.N_55 ));
    SRMux I__1069 (
            .O(N__5055),
            .I(N__5052));
    LocalMux I__1068 (
            .O(N__5052),
            .I(N__5048));
    SRMux I__1067 (
            .O(N__5051),
            .I(N__5045));
    Span4Mux_v I__1066 (
            .O(N__5048),
            .I(N__5038));
    LocalMux I__1065 (
            .O(N__5045),
            .I(N__5038));
    SRMux I__1064 (
            .O(N__5044),
            .I(N__5035));
    SRMux I__1063 (
            .O(N__5043),
            .I(N__5032));
    Span4Mux_v I__1062 (
            .O(N__5038),
            .I(N__5027));
    LocalMux I__1061 (
            .O(N__5035),
            .I(N__5027));
    LocalMux I__1060 (
            .O(N__5032),
            .I(N__5024));
    Span4Mux_v I__1059 (
            .O(N__5027),
            .I(N__5020));
    Span4Mux_v I__1058 (
            .O(N__5024),
            .I(N__5017));
    InMux I__1057 (
            .O(N__5023),
            .I(N__5014));
    Odrv4 I__1056 (
            .O(N__5020),
            .I(RESETn_c_i));
    Odrv4 I__1055 (
            .O(N__5017),
            .I(RESETn_c_i));
    LocalMux I__1054 (
            .O(N__5014),
            .I(RESETn_c_i));
    InMux I__1053 (
            .O(N__5007),
            .I(N__5004));
    LocalMux I__1052 (
            .O(N__5004),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__1051 (
            .O(N__5001),
            .I(N__4997));
    InMux I__1050 (
            .O(N__5000),
            .I(N__4994));
    LocalMux I__1049 (
            .O(N__4997),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__1048 (
            .O(N__4994),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    CascadeMux I__1047 (
            .O(N__4989),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_ ));
    InMux I__1046 (
            .O(N__4986),
            .I(N__4983));
    LocalMux I__1045 (
            .O(N__4983),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__1044 (
            .O(N__4980),
            .I(N__4976));
    InMux I__1043 (
            .O(N__4979),
            .I(N__4973));
    LocalMux I__1042 (
            .O(N__4976),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__1041 (
            .O(N__4973),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    InMux I__1040 (
            .O(N__4968),
            .I(N__4952));
    InMux I__1039 (
            .O(N__4967),
            .I(N__4952));
    InMux I__1038 (
            .O(N__4966),
            .I(N__4952));
    InMux I__1037 (
            .O(N__4965),
            .I(N__4952));
    InMux I__1036 (
            .O(N__4964),
            .I(N__4949));
    InMux I__1035 (
            .O(N__4963),
            .I(N__4942));
    InMux I__1034 (
            .O(N__4962),
            .I(N__4942));
    InMux I__1033 (
            .O(N__4961),
            .I(N__4942));
    LocalMux I__1032 (
            .O(N__4952),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1031 (
            .O(N__4949),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1030 (
            .O(N__4942),
            .I(\U409_TICK.TICK503_9 ));
    InMux I__1029 (
            .O(N__4935),
            .I(N__4925));
    InMux I__1028 (
            .O(N__4934),
            .I(N__4925));
    CascadeMux I__1027 (
            .O(N__4933),
            .I(N__4920));
    CascadeMux I__1026 (
            .O(N__4932),
            .I(N__4917));
    InMux I__1025 (
            .O(N__4931),
            .I(N__4912));
    InMux I__1024 (
            .O(N__4930),
            .I(N__4912));
    LocalMux I__1023 (
            .O(N__4925),
            .I(N__4909));
    InMux I__1022 (
            .O(N__4924),
            .I(N__4900));
    InMux I__1021 (
            .O(N__4923),
            .I(N__4900));
    InMux I__1020 (
            .O(N__4920),
            .I(N__4900));
    InMux I__1019 (
            .O(N__4917),
            .I(N__4900));
    LocalMux I__1018 (
            .O(N__4912),
            .I(\U409_TICK.TICK503_14 ));
    Odrv4 I__1017 (
            .O(N__4909),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__1016 (
            .O(N__4900),
            .I(\U409_TICK.TICK503_14 ));
    CascadeMux I__1015 (
            .O(N__4893),
            .I(N__4890));
    InMux I__1014 (
            .O(N__4890),
            .I(N__4887));
    LocalMux I__1013 (
            .O(N__4887),
            .I(N__4884));
    Odrv4 I__1012 (
            .O(N__4884),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__1011 (
            .O(N__4881),
            .I(N__4863));
    InMux I__1010 (
            .O(N__4880),
            .I(N__4863));
    InMux I__1009 (
            .O(N__4879),
            .I(N__4863));
    InMux I__1008 (
            .O(N__4878),
            .I(N__4863));
    InMux I__1007 (
            .O(N__4877),
            .I(N__4863));
    InMux I__1006 (
            .O(N__4876),
            .I(N__4856));
    InMux I__1005 (
            .O(N__4875),
            .I(N__4856));
    InMux I__1004 (
            .O(N__4874),
            .I(N__4856));
    LocalMux I__1003 (
            .O(N__4863),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__1002 (
            .O(N__4856),
            .I(\U409_TICK.TICK503_10 ));
    InMux I__1001 (
            .O(N__4851),
            .I(N__4847));
    InMux I__1000 (
            .O(N__4850),
            .I(N__4844));
    LocalMux I__999 (
            .O(N__4847),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__998 (
            .O(N__4844),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    ClkMux I__997 (
            .O(N__4839),
            .I(N__4815));
    ClkMux I__996 (
            .O(N__4838),
            .I(N__4815));
    ClkMux I__995 (
            .O(N__4837),
            .I(N__4815));
    ClkMux I__994 (
            .O(N__4836),
            .I(N__4815));
    ClkMux I__993 (
            .O(N__4835),
            .I(N__4815));
    ClkMux I__992 (
            .O(N__4834),
            .I(N__4815));
    ClkMux I__991 (
            .O(N__4833),
            .I(N__4815));
    ClkMux I__990 (
            .O(N__4832),
            .I(N__4815));
    GlobalMux I__989 (
            .O(N__4815),
            .I(N__4812));
    gio2CtrlBuf I__988 (
            .O(N__4812),
            .I(CLK6_c_g));
    CascadeMux I__987 (
            .O(N__4809),
            .I(\U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_ ));
    InMux I__986 (
            .O(N__4806),
            .I(N__4801));
    InMux I__985 (
            .O(N__4805),
            .I(N__4798));
    InMux I__984 (
            .O(N__4804),
            .I(N__4795));
    LocalMux I__983 (
            .O(N__4801),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__982 (
            .O(N__4798),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__981 (
            .O(N__4795),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    InMux I__980 (
            .O(N__4788),
            .I(N__4784));
    InMux I__979 (
            .O(N__4787),
            .I(N__4781));
    LocalMux I__978 (
            .O(N__4784),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    LocalMux I__977 (
            .O(N__4781),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    InMux I__976 (
            .O(N__4776),
            .I(N__4773));
    LocalMux I__975 (
            .O(N__4773),
            .I(\U409_TRANSFER_ACK.N_49 ));
    CascadeMux I__974 (
            .O(N__4770),
            .I(\U409_TRANSFER_ACK.N_29_cascade_ ));
    InMux I__973 (
            .O(N__4767),
            .I(N__4763));
    InMux I__972 (
            .O(N__4766),
            .I(N__4760));
    LocalMux I__971 (
            .O(N__4763),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__970 (
            .O(N__4760),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__969 (
            .O(N__4755),
            .I(N__4751));
    InMux I__968 (
            .O(N__4754),
            .I(N__4748));
    LocalMux I__967 (
            .O(N__4751),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__966 (
            .O(N__4748),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__965 (
            .O(N__4743),
            .I(N__4739));
    InMux I__964 (
            .O(N__4742),
            .I(N__4736));
    LocalMux I__963 (
            .O(N__4739),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__962 (
            .O(N__4736),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    CascadeMux I__961 (
            .O(N__4731),
            .I(N__4726));
    CascadeMux I__960 (
            .O(N__4730),
            .I(N__4723));
    InMux I__959 (
            .O(N__4729),
            .I(N__4718));
    InMux I__958 (
            .O(N__4726),
            .I(N__4718));
    InMux I__957 (
            .O(N__4723),
            .I(N__4715));
    LocalMux I__956 (
            .O(N__4718),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__955 (
            .O(N__4715),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    IoInMux I__954 (
            .O(N__4710),
            .I(N__4707));
    LocalMux I__953 (
            .O(N__4707),
            .I(N__4703));
    CascadeMux I__952 (
            .O(N__4706),
            .I(N__4700));
    Span12Mux_s10_v I__951 (
            .O(N__4703),
            .I(N__4697));
    InMux I__950 (
            .O(N__4700),
            .I(N__4694));
    Odrv12 I__949 (
            .O(N__4697),
            .I(TICK50_c));
    LocalMux I__948 (
            .O(N__4694),
            .I(TICK50_c));
    InMux I__947 (
            .O(N__4689),
            .I(N__4685));
    InMux I__946 (
            .O(N__4688),
            .I(N__4682));
    LocalMux I__945 (
            .O(N__4685),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__944 (
            .O(N__4682),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__943 (
            .O(N__4677),
            .I(N__4673));
    InMux I__942 (
            .O(N__4676),
            .I(N__4670));
    LocalMux I__941 (
            .O(N__4673),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__940 (
            .O(N__4670),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    CascadeMux I__939 (
            .O(N__4665),
            .I(N__4661));
    InMux I__938 (
            .O(N__4664),
            .I(N__4654));
    InMux I__937 (
            .O(N__4661),
            .I(N__4654));
    InMux I__936 (
            .O(N__4660),
            .I(N__4651));
    InMux I__935 (
            .O(N__4659),
            .I(N__4648));
    LocalMux I__934 (
            .O(N__4654),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__933 (
            .O(N__4651),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__932 (
            .O(N__4648),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__931 (
            .O(N__4641),
            .I(N__4638));
    LocalMux I__930 (
            .O(N__4638),
            .I(\U409_TICK.TICK503_11 ));
    InMux I__929 (
            .O(N__4635),
            .I(N__4631));
    InMux I__928 (
            .O(N__4634),
            .I(N__4628));
    LocalMux I__927 (
            .O(N__4631),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__926 (
            .O(N__4628),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    CascadeMux I__925 (
            .O(N__4623),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    InMux I__924 (
            .O(N__4620),
            .I(N__4616));
    InMux I__923 (
            .O(N__4619),
            .I(N__4613));
    LocalMux I__922 (
            .O(N__4616),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__921 (
            .O(N__4613),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    InMux I__920 (
            .O(N__4608),
            .I(N__4605));
    LocalMux I__919 (
            .O(N__4605),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    CascadeMux I__918 (
            .O(N__4602),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    CascadeMux I__917 (
            .O(N__4599),
            .I(N__4596));
    InMux I__916 (
            .O(N__4596),
            .I(N__4592));
    InMux I__915 (
            .O(N__4595),
            .I(N__4589));
    LocalMux I__914 (
            .O(N__4592),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__913 (
            .O(N__4589),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__912 (
            .O(N__4584),
            .I(N__4581));
    LocalMux I__911 (
            .O(N__4581),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    CascadeMux I__910 (
            .O(N__4578),
            .I(N__4575));
    InMux I__909 (
            .O(N__4575),
            .I(N__4571));
    InMux I__908 (
            .O(N__4574),
            .I(N__4568));
    LocalMux I__907 (
            .O(N__4571),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__906 (
            .O(N__4568),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    CascadeMux I__905 (
            .O(N__4563),
            .I(N__4560));
    InMux I__904 (
            .O(N__4560),
            .I(N__4557));
    LocalMux I__903 (
            .O(N__4557),
            .I(N__4554));
    Odrv4 I__902 (
            .O(N__4554),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__901 (
            .O(N__4551),
            .I(N__4547));
    InMux I__900 (
            .O(N__4550),
            .I(N__4544));
    LocalMux I__899 (
            .O(N__4547),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__898 (
            .O(N__4544),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    CEMux I__897 (
            .O(N__4539),
            .I(N__4536));
    LocalMux I__896 (
            .O(N__4536),
            .I(N__4533));
    Odrv4 I__895 (
            .O(N__4533),
            .I(\U409_TRANSFER_ACK.N_22_0_0 ));
    InMux I__894 (
            .O(N__4530),
            .I(N__4523));
    InMux I__893 (
            .O(N__4529),
            .I(N__4518));
    InMux I__892 (
            .O(N__4528),
            .I(N__4518));
    InMux I__891 (
            .O(N__4527),
            .I(N__4513));
    InMux I__890 (
            .O(N__4526),
            .I(N__4513));
    LocalMux I__889 (
            .O(N__4523),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__888 (
            .O(N__4518),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__887 (
            .O(N__4513),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    InMux I__886 (
            .O(N__4506),
            .I(N__4496));
    InMux I__885 (
            .O(N__4505),
            .I(N__4496));
    InMux I__884 (
            .O(N__4504),
            .I(N__4496));
    InMux I__883 (
            .O(N__4503),
            .I(N__4493));
    LocalMux I__882 (
            .O(N__4496),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__881 (
            .O(N__4493),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__880 (
            .O(N__4488),
            .I(N__4485));
    LocalMux I__879 (
            .O(N__4485),
            .I(\U409_TRANSFER_ACK.N_24 ));
    InMux I__878 (
            .O(N__4482),
            .I(N__4472));
    InMux I__877 (
            .O(N__4481),
            .I(N__4472));
    InMux I__876 (
            .O(N__4480),
            .I(N__4472));
    InMux I__875 (
            .O(N__4479),
            .I(N__4469));
    LocalMux I__874 (
            .O(N__4472),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__873 (
            .O(N__4469),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    CascadeMux I__872 (
            .O(N__4464),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    InMux I__871 (
            .O(N__4461),
            .I(N__4458));
    LocalMux I__870 (
            .O(N__4458),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__869 (
            .O(N__4455),
            .I(N__4451));
    InMux I__868 (
            .O(N__4454),
            .I(N__4448));
    LocalMux I__867 (
            .O(N__4451),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__866 (
            .O(N__4448),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    InMux I__865 (
            .O(N__4443),
            .I(N__4439));
    InMux I__864 (
            .O(N__4442),
            .I(N__4436));
    LocalMux I__863 (
            .O(N__4439),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__862 (
            .O(N__4436),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    InMux I__861 (
            .O(N__4431),
            .I(N__4427));
    InMux I__860 (
            .O(N__4430),
            .I(N__4424));
    LocalMux I__859 (
            .O(N__4427),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__858 (
            .O(N__4424),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    CascadeMux I__857 (
            .O(N__4419),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    InMux I__856 (
            .O(N__4416),
            .I(N__4413));
    LocalMux I__855 (
            .O(N__4413),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__854 (
            .O(N__4410),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__853 (
            .O(N__4407),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__852 (
            .O(N__4404),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__851 (
            .O(N__4401),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__850 (
            .O(N__4398),
            .I(N__4395));
    LocalMux I__849 (
            .O(N__4395),
            .I(N__4391));
    InMux I__848 (
            .O(N__4394),
            .I(N__4388));
    Span4Mux_h I__847 (
            .O(N__4391),
            .I(N__4383));
    LocalMux I__846 (
            .O(N__4388),
            .I(N__4383));
    Odrv4 I__845 (
            .O(N__4383),
            .I(CIA_ENABLEm));
    InMux I__844 (
            .O(N__4380),
            .I(N__4377));
    LocalMux I__843 (
            .O(N__4377),
            .I(N__4374));
    Span4Mux_v I__842 (
            .O(N__4374),
            .I(N__4369));
    InMux I__841 (
            .O(N__4373),
            .I(N__4366));
    InMux I__840 (
            .O(N__4372),
            .I(N__4363));
    Sp12to4 I__839 (
            .O(N__4369),
            .I(N__4358));
    LocalMux I__838 (
            .O(N__4366),
            .I(N__4358));
    LocalMux I__837 (
            .O(N__4363),
            .I(N__4355));
    Span12Mux_h I__836 (
            .O(N__4358),
            .I(N__4350));
    Span12Mux_v I__835 (
            .O(N__4355),
            .I(N__4350));
    Odrv12 I__834 (
            .O(N__4350),
            .I(\U409_CIA.g0Z0Z_14 ));
    CascadeMux I__833 (
            .O(N__4347),
            .I(N__4344));
    InMux I__832 (
            .O(N__4344),
            .I(N__4341));
    LocalMux I__831 (
            .O(N__4341),
            .I(N__4337));
    InMux I__830 (
            .O(N__4340),
            .I(N__4334));
    Span4Mux_h I__829 (
            .O(N__4337),
            .I(N__4328));
    LocalMux I__828 (
            .O(N__4334),
            .I(N__4328));
    CascadeMux I__827 (
            .O(N__4333),
            .I(N__4325));
    Span4Mux_v I__826 (
            .O(N__4328),
            .I(N__4322));
    InMux I__825 (
            .O(N__4325),
            .I(N__4319));
    Span4Mux_h I__824 (
            .O(N__4322),
            .I(N__4316));
    LocalMux I__823 (
            .O(N__4319),
            .I(N__4313));
    Span4Mux_h I__822 (
            .O(N__4316),
            .I(N__4310));
    Span12Mux_v I__821 (
            .O(N__4313),
            .I(N__4307));
    Odrv4 I__820 (
            .O(N__4310),
            .I(\U409_CIA.g0Z0Z_13 ));
    Odrv12 I__819 (
            .O(N__4307),
            .I(\U409_CIA.g0Z0Z_13 ));
    CascadeMux I__818 (
            .O(N__4302),
            .I(N__4299));
    InMux I__817 (
            .O(N__4299),
            .I(N__4295));
    InMux I__816 (
            .O(N__4298),
            .I(N__4292));
    LocalMux I__815 (
            .O(N__4295),
            .I(N__4286));
    LocalMux I__814 (
            .O(N__4292),
            .I(N__4286));
    InMux I__813 (
            .O(N__4291),
            .I(N__4282));
    Span4Mux_v I__812 (
            .O(N__4286),
            .I(N__4279));
    InMux I__811 (
            .O(N__4285),
            .I(N__4276));
    LocalMux I__810 (
            .O(N__4282),
            .I(N__4273));
    Odrv4 I__809 (
            .O(N__4279),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__808 (
            .O(N__4276),
            .I(\U409_CIA.VMAZ0 ));
    Odrv4 I__807 (
            .O(N__4273),
            .I(\U409_CIA.VMAZ0 ));
    InMux I__806 (
            .O(N__4266),
            .I(N__4263));
    LocalMux I__805 (
            .O(N__4263),
            .I(N__4259));
    InMux I__804 (
            .O(N__4262),
            .I(N__4256));
    Span4Mux_v I__803 (
            .O(N__4259),
            .I(N__4250));
    LocalMux I__802 (
            .O(N__4256),
            .I(N__4250));
    InMux I__801 (
            .O(N__4255),
            .I(N__4247));
    Odrv4 I__800 (
            .O(N__4250),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    LocalMux I__799 (
            .O(N__4247),
            .I(\U409_CIA.CIA_HOLDZ0 ));
    IoInMux I__798 (
            .O(N__4242),
            .I(N__4239));
    LocalMux I__797 (
            .O(N__4239),
            .I(N__4236));
    Span4Mux_s1_v I__796 (
            .O(N__4236),
            .I(N__4233));
    Sp12to4 I__795 (
            .O(N__4233),
            .I(N__4229));
    InMux I__794 (
            .O(N__4232),
            .I(N__4226));
    Span12Mux_h I__793 (
            .O(N__4229),
            .I(N__4223));
    LocalMux I__792 (
            .O(N__4226),
            .I(N__4220));
    Span12Mux_v I__791 (
            .O(N__4223),
            .I(N__4216));
    Span4Mux_v I__790 (
            .O(N__4220),
            .I(N__4213));
    InMux I__789 (
            .O(N__4219),
            .I(N__4210));
    Odrv12 I__788 (
            .O(N__4216),
            .I(CLKCIA_c));
    Odrv4 I__787 (
            .O(N__4213),
            .I(CLKCIA_c));
    LocalMux I__786 (
            .O(N__4210),
            .I(CLKCIA_c));
    InMux I__785 (
            .O(N__4203),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__784 (
            .O(N__4200),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    InMux I__783 (
            .O(N__4197),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__782 (
            .O(N__4194),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__781 (
            .O(N__4191),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__780 (
            .O(N__4188),
            .I(bfn_10_6_0_));
    InMux I__779 (
            .O(N__4185),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__778 (
            .O(N__4182),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__777 (
            .O(N__4179),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__776 (
            .O(N__4176),
            .I(N__4172));
    InMux I__775 (
            .O(N__4175),
            .I(N__4169));
    LocalMux I__774 (
            .O(N__4172),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__773 (
            .O(N__4169),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__772 (
            .O(N__4164),
            .I(N__4161));
    LocalMux I__771 (
            .O(N__4161),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__770 (
            .O(N__4158),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__769 (
            .O(N__4155),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__768 (
            .O(N__4152),
            .I(N__4148));
    InMux I__767 (
            .O(N__4151),
            .I(N__4145));
    LocalMux I__766 (
            .O(N__4148),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__765 (
            .O(N__4145),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    CascadeMux I__764 (
            .O(N__4140),
            .I(N__4137));
    InMux I__763 (
            .O(N__4137),
            .I(N__4134));
    LocalMux I__762 (
            .O(N__4134),
            .I(N__4131));
    Odrv12 I__761 (
            .O(N__4131),
            .I(ROMENm));
    CascadeMux I__760 (
            .O(N__4128),
            .I(\U409_TRANSFER_ACK.N_24_cascade_ ));
    InMux I__759 (
            .O(N__4125),
            .I(N__4122));
    LocalMux I__758 (
            .O(N__4122),
            .I(\U409_TRANSFER_ACK.N_22 ));
    InMux I__757 (
            .O(N__4119),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__756 (
            .O(N__4116),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    InMux I__755 (
            .O(N__4113),
            .I(N__4109));
    InMux I__754 (
            .O(N__4112),
            .I(N__4106));
    LocalMux I__753 (
            .O(N__4109),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__752 (
            .O(N__4106),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__751 (
            .O(N__4101),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__750 (
            .O(N__4098),
            .I(N__4094));
    InMux I__749 (
            .O(N__4097),
            .I(N__4091));
    LocalMux I__748 (
            .O(N__4094),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__747 (
            .O(N__4091),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    InMux I__746 (
            .O(N__4086),
            .I(N__4083));
    LocalMux I__745 (
            .O(N__4083),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__744 (
            .O(N__4080),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__743 (
            .O(N__4077),
            .I(N__4073));
    InMux I__742 (
            .O(N__4076),
            .I(N__4070));
    LocalMux I__741 (
            .O(N__4073),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__740 (
            .O(N__4070),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    InMux I__739 (
            .O(N__4065),
            .I(N__4062));
    LocalMux I__738 (
            .O(N__4062),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__737 (
            .O(N__4059),
            .I(bfn_9_8_0_));
    CascadeMux I__736 (
            .O(N__4056),
            .I(N__4053));
    InMux I__735 (
            .O(N__4053),
            .I(N__4049));
    InMux I__734 (
            .O(N__4052),
            .I(N__4046));
    LocalMux I__733 (
            .O(N__4049),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__732 (
            .O(N__4046),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    InMux I__731 (
            .O(N__4041),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__730 (
            .O(N__4038),
            .I(N__4034));
    InMux I__729 (
            .O(N__4037),
            .I(N__4031));
    LocalMux I__728 (
            .O(N__4034),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__727 (
            .O(N__4031),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    InMux I__726 (
            .O(N__4026),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__725 (
            .O(N__4023),
            .I(N__4019));
    InMux I__724 (
            .O(N__4022),
            .I(N__4016));
    LocalMux I__723 (
            .O(N__4019),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__722 (
            .O(N__4016),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__721 (
            .O(N__4011),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__720 (
            .O(N__4008),
            .I(N__4004));
    InMux I__719 (
            .O(N__4007),
            .I(N__4001));
    LocalMux I__718 (
            .O(N__4004),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__717 (
            .O(N__4001),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__716 (
            .O(N__3996),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__715 (
            .O(N__3993),
            .I(N__3989));
    InMux I__714 (
            .O(N__3992),
            .I(N__3986));
    LocalMux I__713 (
            .O(N__3989),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__712 (
            .O(N__3986),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    InMux I__711 (
            .O(N__3981),
            .I(N__3978));
    LocalMux I__710 (
            .O(N__3978),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__709 (
            .O(N__3975),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__708 (
            .O(N__3972),
            .I(N__3969));
    LocalMux I__707 (
            .O(N__3969),
            .I(\U409_TICK.TICK603_11 ));
    InMux I__706 (
            .O(N__3966),
            .I(N__3963));
    LocalMux I__705 (
            .O(N__3963),
            .I(N__3960));
    Span4Mux_v I__704 (
            .O(N__3960),
            .I(N__3957));
    Sp12to4 I__703 (
            .O(N__3957),
            .I(N__3954));
    Span12Mux_h I__702 (
            .O(N__3954),
            .I(N__3951));
    Odrv12 I__701 (
            .O(N__3951),
            .I(A_c_13));
    IoInMux I__700 (
            .O(N__3948),
            .I(N__3945));
    LocalMux I__699 (
            .O(N__3945),
            .I(N__3942));
    IoSpan4Mux I__698 (
            .O(N__3942),
            .I(N__3939));
    Sp12to4 I__697 (
            .O(N__3939),
            .I(N__3936));
    Span12Mux_s7_h I__696 (
            .O(N__3936),
            .I(N__3933));
    Span12Mux_h I__695 (
            .O(N__3933),
            .I(N__3930));
    Odrv12 I__694 (
            .O(N__3930),
            .I(U409_ADDRESS_DECODE_un1_nCIACS1_i));
    InMux I__693 (
            .O(N__3927),
            .I(N__3924));
    LocalMux I__692 (
            .O(N__3924),
            .I(N__3921));
    Span4Mux_v I__691 (
            .O(N__3921),
            .I(N__3918));
    Sp12to4 I__690 (
            .O(N__3918),
            .I(N__3915));
    Odrv12 I__689 (
            .O(N__3915),
            .I(A_c_12));
    IoInMux I__688 (
            .O(N__3912),
            .I(N__3909));
    LocalMux I__687 (
            .O(N__3909),
            .I(N__3906));
    Span4Mux_s0_h I__686 (
            .O(N__3906),
            .I(N__3903));
    Sp12to4 I__685 (
            .O(N__3903),
            .I(N__3900));
    Span12Mux_s11_v I__684 (
            .O(N__3900),
            .I(N__3897));
    Span12Mux_h I__683 (
            .O(N__3897),
            .I(N__3894));
    Odrv12 I__682 (
            .O(N__3894),
            .I(U409_ADDRESS_DECODE_un1_nCIACS0_i));
    InMux I__681 (
            .O(N__3891),
            .I(N__3886));
    InMux I__680 (
            .O(N__3890),
            .I(N__3883));
    InMux I__679 (
            .O(N__3889),
            .I(N__3880));
    LocalMux I__678 (
            .O(N__3886),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__677 (
            .O(N__3883),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__676 (
            .O(N__3880),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    CascadeMux I__675 (
            .O(N__3873),
            .I(N__3867));
    InMux I__674 (
            .O(N__3872),
            .I(N__3862));
    InMux I__673 (
            .O(N__3871),
            .I(N__3862));
    InMux I__672 (
            .O(N__3870),
            .I(N__3859));
    InMux I__671 (
            .O(N__3867),
            .I(N__3856));
    LocalMux I__670 (
            .O(N__3862),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__669 (
            .O(N__3859),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__668 (
            .O(N__3856),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    CascadeMux I__667 (
            .O(N__3849),
            .I(N__3846));
    InMux I__666 (
            .O(N__3846),
            .I(N__3842));
    InMux I__665 (
            .O(N__3845),
            .I(N__3839));
    LocalMux I__664 (
            .O(N__3842),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__663 (
            .O(N__3839),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    InMux I__662 (
            .O(N__3834),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__661 (
            .O(N__3831),
            .I(N__3827));
    InMux I__660 (
            .O(N__3830),
            .I(N__3824));
    LocalMux I__659 (
            .O(N__3827),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__658 (
            .O(N__3824),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    InMux I__657 (
            .O(N__3819),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__656 (
            .O(N__3816),
            .I(N__3812));
    InMux I__655 (
            .O(N__3815),
            .I(N__3809));
    LocalMux I__654 (
            .O(N__3812),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__653 (
            .O(N__3809),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__652 (
            .O(N__3804),
            .I(N__3801));
    LocalMux I__651 (
            .O(N__3801),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__650 (
            .O(N__3798),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__649 (
            .O(N__3795),
            .I(N__3791));
    InMux I__648 (
            .O(N__3794),
            .I(N__3788));
    LocalMux I__647 (
            .O(N__3791),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__646 (
            .O(N__3788),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__645 (
            .O(N__3783),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    CascadeMux I__644 (
            .O(N__3780),
            .I(N__3777));
    InMux I__643 (
            .O(N__3777),
            .I(N__3773));
    InMux I__642 (
            .O(N__3776),
            .I(N__3770));
    LocalMux I__641 (
            .O(N__3773),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__640 (
            .O(N__3770),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    CascadeMux I__639 (
            .O(N__3765),
            .I(N__3762));
    InMux I__638 (
            .O(N__3762),
            .I(N__3759));
    LocalMux I__637 (
            .O(N__3759),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__636 (
            .O(N__3756),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    CascadeMux I__635 (
            .O(N__3753),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    CascadeMux I__634 (
            .O(N__3750),
            .I(\U409_TICK.TICK603_10_cascade_ ));
    CascadeMux I__633 (
            .O(N__3747),
            .I(\U409_TICK.TICK603_8_cascade_ ));
    InMux I__632 (
            .O(N__3744),
            .I(N__3727));
    InMux I__631 (
            .O(N__3743),
            .I(N__3727));
    InMux I__630 (
            .O(N__3742),
            .I(N__3727));
    InMux I__629 (
            .O(N__3741),
            .I(N__3727));
    InMux I__628 (
            .O(N__3740),
            .I(N__3727));
    InMux I__627 (
            .O(N__3739),
            .I(N__3722));
    InMux I__626 (
            .O(N__3738),
            .I(N__3722));
    LocalMux I__625 (
            .O(N__3727),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__624 (
            .O(N__3722),
            .I(\U409_TICK.TICK603_14 ));
    CascadeMux I__623 (
            .O(N__3717),
            .I(N__3714));
    InMux I__622 (
            .O(N__3714),
            .I(N__3709));
    CascadeMux I__621 (
            .O(N__3713),
            .I(N__3706));
    CascadeMux I__620 (
            .O(N__3712),
            .I(N__3700));
    LocalMux I__619 (
            .O(N__3709),
            .I(N__3696));
    InMux I__618 (
            .O(N__3706),
            .I(N__3691));
    InMux I__617 (
            .O(N__3705),
            .I(N__3691));
    InMux I__616 (
            .O(N__3704),
            .I(N__3688));
    InMux I__615 (
            .O(N__3703),
            .I(N__3681));
    InMux I__614 (
            .O(N__3700),
            .I(N__3681));
    InMux I__613 (
            .O(N__3699),
            .I(N__3681));
    Odrv4 I__612 (
            .O(N__3696),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__611 (
            .O(N__3691),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__610 (
            .O(N__3688),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__609 (
            .O(N__3681),
            .I(\U409_TICK.TICK603_9 ));
    CascadeMux I__608 (
            .O(N__3672),
            .I(N__3667));
    InMux I__607 (
            .O(N__3671),
            .I(N__3658));
    InMux I__606 (
            .O(N__3670),
            .I(N__3658));
    InMux I__605 (
            .O(N__3667),
            .I(N__3647));
    InMux I__604 (
            .O(N__3666),
            .I(N__3647));
    InMux I__603 (
            .O(N__3665),
            .I(N__3647));
    InMux I__602 (
            .O(N__3664),
            .I(N__3647));
    InMux I__601 (
            .O(N__3663),
            .I(N__3647));
    LocalMux I__600 (
            .O(N__3658),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__599 (
            .O(N__3647),
            .I(\U409_TICK.TICK603_10 ));
    CascadeMux I__598 (
            .O(N__3642),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    CascadeMux I__597 (
            .O(N__3639),
            .I(\U409_CIA.N_9_cascade_ ));
    InMux I__596 (
            .O(N__3636),
            .I(N__3621));
    InMux I__595 (
            .O(N__3635),
            .I(N__3621));
    InMux I__594 (
            .O(N__3634),
            .I(N__3621));
    InMux I__593 (
            .O(N__3633),
            .I(N__3621));
    InMux I__592 (
            .O(N__3632),
            .I(N__3614));
    InMux I__591 (
            .O(N__3631),
            .I(N__3614));
    InMux I__590 (
            .O(N__3630),
            .I(N__3614));
    LocalMux I__589 (
            .O(N__3621),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__588 (
            .O(N__3614),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    CascadeMux I__587 (
            .O(N__3609),
            .I(\U409_CIA.N_20_cascade_ ));
    InMux I__586 (
            .O(N__3606),
            .I(N__3600));
    InMux I__585 (
            .O(N__3605),
            .I(N__3600));
    LocalMux I__584 (
            .O(N__3600),
            .I(\U409_CIA.CLKCIA8_0_a2_0 ));
    InMux I__583 (
            .O(N__3597),
            .I(N__3594));
    LocalMux I__582 (
            .O(N__3594),
            .I(\U409_CIA.CLKCIA6_0_a2_1 ));
    CascadeMux I__581 (
            .O(N__3591),
            .I(N__3581));
    InMux I__580 (
            .O(N__3590),
            .I(N__3578));
    InMux I__579 (
            .O(N__3589),
            .I(N__3569));
    InMux I__578 (
            .O(N__3588),
            .I(N__3569));
    InMux I__577 (
            .O(N__3587),
            .I(N__3569));
    InMux I__576 (
            .O(N__3586),
            .I(N__3569));
    InMux I__575 (
            .O(N__3585),
            .I(N__3562));
    InMux I__574 (
            .O(N__3584),
            .I(N__3562));
    InMux I__573 (
            .O(N__3581),
            .I(N__3562));
    LocalMux I__572 (
            .O(N__3578),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__571 (
            .O(N__3569),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__570 (
            .O(N__3562),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    CascadeMux I__569 (
            .O(N__3555),
            .I(\U409_CIA.CLKCIAZ0_cascade_ ));
    InMux I__568 (
            .O(N__3552),
            .I(N__3544));
    InMux I__567 (
            .O(N__3551),
            .I(N__3537));
    InMux I__566 (
            .O(N__3550),
            .I(N__3537));
    InMux I__565 (
            .O(N__3549),
            .I(N__3537));
    InMux I__564 (
            .O(N__3548),
            .I(N__3532));
    InMux I__563 (
            .O(N__3547),
            .I(N__3532));
    LocalMux I__562 (
            .O(N__3544),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__561 (
            .O(N__3537),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__560 (
            .O(N__3532),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    ClkMux I__559 (
            .O(N__3525),
            .I(N__3513));
    ClkMux I__558 (
            .O(N__3524),
            .I(N__3513));
    ClkMux I__557 (
            .O(N__3523),
            .I(N__3513));
    ClkMux I__556 (
            .O(N__3522),
            .I(N__3513));
    GlobalMux I__555 (
            .O(N__3513),
            .I(N__3510));
    gio2CtrlBuf I__554 (
            .O(N__3510),
            .I(CLK28_IN_c_g));
    IoInMux I__553 (
            .O(N__3507),
            .I(N__3504));
    LocalMux I__552 (
            .O(N__3504),
            .I(N__3501));
    Span4Mux_s1_v I__551 (
            .O(N__3501),
            .I(N__3498));
    Sp12to4 I__550 (
            .O(N__3498),
            .I(N__3495));
    Span12Mux_h I__549 (
            .O(N__3495),
            .I(N__3491));
    InMux I__548 (
            .O(N__3494),
            .I(N__3488));
    Odrv12 I__547 (
            .O(N__3491),
            .I(TICK60_c));
    LocalMux I__546 (
            .O(N__3488),
            .I(TICK60_c));
    InMux I__545 (
            .O(N__3483),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    CascadeMux I__544 (
            .O(N__3480),
            .I(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ));
    InMux I__543 (
            .O(N__3477),
            .I(N__3474));
    LocalMux I__542 (
            .O(N__3474),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ));
    CascadeMux I__541 (
            .O(N__3471),
            .I(N__3468));
    InMux I__540 (
            .O(N__3468),
            .I(N__3462));
    InMux I__539 (
            .O(N__3467),
            .I(N__3462));
    LocalMux I__538 (
            .O(N__3462),
            .I(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ));
    InMux I__537 (
            .O(N__3459),
            .I(N__3453));
    InMux I__536 (
            .O(N__3458),
            .I(N__3448));
    InMux I__535 (
            .O(N__3457),
            .I(N__3448));
    InMux I__534 (
            .O(N__3456),
            .I(N__3445));
    LocalMux I__533 (
            .O(N__3453),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__532 (
            .O(N__3448),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__531 (
            .O(N__3445),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    InMux I__530 (
            .O(N__3438),
            .I(N__3430));
    InMux I__529 (
            .O(N__3437),
            .I(N__3430));
    InMux I__528 (
            .O(N__3436),
            .I(N__3425));
    InMux I__527 (
            .O(N__3435),
            .I(N__3425));
    LocalMux I__526 (
            .O(N__3430),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__525 (
            .O(N__3425),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    CascadeMux I__524 (
            .O(N__3420),
            .I(N__3416));
    CascadeMux I__523 (
            .O(N__3419),
            .I(N__3412));
    InMux I__522 (
            .O(N__3416),
            .I(N__3406));
    InMux I__521 (
            .O(N__3415),
            .I(N__3406));
    InMux I__520 (
            .O(N__3412),
            .I(N__3401));
    InMux I__519 (
            .O(N__3411),
            .I(N__3401));
    LocalMux I__518 (
            .O(N__3406),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__517 (
            .O(N__3401),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    IoInMux I__516 (
            .O(N__3396),
            .I(N__3393));
    LocalMux I__515 (
            .O(N__3393),
            .I(N__3390));
    Span4Mux_s3_v I__514 (
            .O(N__3390),
            .I(N__3387));
    Span4Mux_h I__513 (
            .O(N__3387),
            .I(N__3384));
    Sp12to4 I__512 (
            .O(N__3384),
            .I(N__3381));
    Span12Mux_v I__511 (
            .O(N__3381),
            .I(N__3378));
    Odrv12 I__510 (
            .O(N__3378),
            .I(U409_ADDRESS_DECODE_un1_nRAMSPACE_i));
    CascadeMux I__509 (
            .O(N__3375),
            .I(N__3370));
    InMux I__508 (
            .O(N__3374),
            .I(N__3361));
    InMux I__507 (
            .O(N__3373),
            .I(N__3361));
    InMux I__506 (
            .O(N__3370),
            .I(N__3361));
    InMux I__505 (
            .O(N__3369),
            .I(N__3358));
    InMux I__504 (
            .O(N__3368),
            .I(N__3355));
    LocalMux I__503 (
            .O(N__3361),
            .I(N__3352));
    LocalMux I__502 (
            .O(N__3358),
            .I(N__3347));
    LocalMux I__501 (
            .O(N__3355),
            .I(N__3344));
    Span4Mux_v I__500 (
            .O(N__3352),
            .I(N__3341));
    InMux I__499 (
            .O(N__3351),
            .I(N__3338));
    InMux I__498 (
            .O(N__3350),
            .I(N__3335));
    Span12Mux_v I__497 (
            .O(N__3347),
            .I(N__3330));
    Span12Mux_v I__496 (
            .O(N__3344),
            .I(N__3330));
    Sp12to4 I__495 (
            .O(N__3341),
            .I(N__3323));
    LocalMux I__494 (
            .O(N__3338),
            .I(N__3323));
    LocalMux I__493 (
            .O(N__3335),
            .I(N__3323));
    Odrv12 I__492 (
            .O(N__3330),
            .I(A_c_21));
    Odrv12 I__491 (
            .O(N__3323),
            .I(A_c_21));
    CascadeMux I__490 (
            .O(N__3318),
            .I(N__3315));
    InMux I__489 (
            .O(N__3315),
            .I(N__3312));
    LocalMux I__488 (
            .O(N__3312),
            .I(N__3308));
    InMux I__487 (
            .O(N__3311),
            .I(N__3305));
    Odrv4 I__486 (
            .O(N__3308),
            .I(\U409_ADDRESS_DECODE.un1_nRAMSPACEZ0Z_2 ));
    LocalMux I__485 (
            .O(N__3305),
            .I(\U409_ADDRESS_DECODE.un1_nRAMSPACEZ0Z_2 ));
    InMux I__484 (
            .O(N__3300),
            .I(N__3297));
    LocalMux I__483 (
            .O(N__3297),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ));
    IoInMux I__482 (
            .O(N__3294),
            .I(N__3291));
    LocalMux I__481 (
            .O(N__3291),
            .I(N__3288));
    IoSpan4Mux I__480 (
            .O(N__3288),
            .I(N__3285));
    Span4Mux_s0_v I__479 (
            .O(N__3285),
            .I(N__3282));
    Sp12to4 I__478 (
            .O(N__3282),
            .I(N__3279));
    Span12Mux_s11_v I__477 (
            .O(N__3279),
            .I(N__3276));
    Span12Mux_h I__476 (
            .O(N__3276),
            .I(N__3273));
    Odrv12 I__475 (
            .O(N__3273),
            .I(nBUFEN_c));
    InMux I__474 (
            .O(N__3270),
            .I(N__3264));
    InMux I__473 (
            .O(N__3269),
            .I(N__3258));
    InMux I__472 (
            .O(N__3268),
            .I(N__3255));
    InMux I__471 (
            .O(N__3267),
            .I(N__3252));
    LocalMux I__470 (
            .O(N__3264),
            .I(N__3249));
    InMux I__469 (
            .O(N__3263),
            .I(N__3244));
    InMux I__468 (
            .O(N__3262),
            .I(N__3244));
    InMux I__467 (
            .O(N__3261),
            .I(N__3241));
    LocalMux I__466 (
            .O(N__3258),
            .I(N__3238));
    LocalMux I__465 (
            .O(N__3255),
            .I(N__3233));
    LocalMux I__464 (
            .O(N__3252),
            .I(N__3233));
    Span4Mux_v I__463 (
            .O(N__3249),
            .I(N__3228));
    LocalMux I__462 (
            .O(N__3244),
            .I(N__3228));
    LocalMux I__461 (
            .O(N__3241),
            .I(N__3225));
    Span4Mux_v I__460 (
            .O(N__3238),
            .I(N__3219));
    Span4Mux_v I__459 (
            .O(N__3233),
            .I(N__3219));
    Span4Mux_v I__458 (
            .O(N__3228),
            .I(N__3214));
    Span4Mux_v I__457 (
            .O(N__3225),
            .I(N__3214));
    InMux I__456 (
            .O(N__3224),
            .I(N__3211));
    Sp12to4 I__455 (
            .O(N__3219),
            .I(N__3204));
    Sp12to4 I__454 (
            .O(N__3214),
            .I(N__3204));
    LocalMux I__453 (
            .O(N__3211),
            .I(N__3204));
    Odrv12 I__452 (
            .O(N__3204),
            .I(A_c_23));
    CascadeMux I__451 (
            .O(N__3201),
            .I(N__3198));
    InMux I__450 (
            .O(N__3198),
            .I(N__3195));
    LocalMux I__449 (
            .O(N__3195),
            .I(N__3192));
    Span4Mux_v I__448 (
            .O(N__3192),
            .I(N__3188));
    InMux I__447 (
            .O(N__3191),
            .I(N__3185));
    Odrv4 I__446 (
            .O(N__3188),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ));
    LocalMux I__445 (
            .O(N__3185),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ));
    IoInMux I__444 (
            .O(N__3180),
            .I(N__3177));
    LocalMux I__443 (
            .O(N__3177),
            .I(N__3174));
    Span4Mux_s3_v I__442 (
            .O(N__3174),
            .I(N__3171));
    Span4Mux_h I__441 (
            .O(N__3171),
            .I(N__3168));
    Span4Mux_h I__440 (
            .O(N__3168),
            .I(N__3165));
    Sp12to4 I__439 (
            .O(N__3165),
            .I(N__3162));
    Span12Mux_s11_v I__438 (
            .O(N__3162),
            .I(N__3159));
    Odrv12 I__437 (
            .O(N__3159),
            .I(U409_ADDRESS_DECODE_un1_nREGSPACE_i));
    InMux I__436 (
            .O(N__3156),
            .I(N__3151));
    InMux I__435 (
            .O(N__3155),
            .I(N__3148));
    InMux I__434 (
            .O(N__3154),
            .I(N__3145));
    LocalMux I__433 (
            .O(N__3151),
            .I(N__3141));
    LocalMux I__432 (
            .O(N__3148),
            .I(N__3138));
    LocalMux I__431 (
            .O(N__3145),
            .I(N__3135));
    InMux I__430 (
            .O(N__3144),
            .I(N__3132));
    Span4Mux_h I__429 (
            .O(N__3141),
            .I(N__3127));
    Span4Mux_h I__428 (
            .O(N__3138),
            .I(N__3122));
    Span4Mux_v I__427 (
            .O(N__3135),
            .I(N__3122));
    LocalMux I__426 (
            .O(N__3132),
            .I(N__3119));
    InMux I__425 (
            .O(N__3131),
            .I(N__3114));
    InMux I__424 (
            .O(N__3130),
            .I(N__3114));
    Odrv4 I__423 (
            .O(N__3127),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ));
    Odrv4 I__422 (
            .O(N__3122),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ));
    Odrv12 I__421 (
            .O(N__3119),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ));
    LocalMux I__420 (
            .O(N__3114),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ));
    InMux I__419 (
            .O(N__3105),
            .I(N__3102));
    LocalMux I__418 (
            .O(N__3102),
            .I(N__3096));
    InMux I__417 (
            .O(N__3101),
            .I(N__3093));
    CascadeMux I__416 (
            .O(N__3100),
            .I(N__3090));
    InMux I__415 (
            .O(N__3099),
            .I(N__3086));
    Span4Mux_v I__414 (
            .O(N__3096),
            .I(N__3081));
    LocalMux I__413 (
            .O(N__3093),
            .I(N__3081));
    InMux I__412 (
            .O(N__3090),
            .I(N__3078));
    CascadeMux I__411 (
            .O(N__3089),
            .I(N__3075));
    LocalMux I__410 (
            .O(N__3086),
            .I(N__3071));
    Span4Mux_h I__409 (
            .O(N__3081),
            .I(N__3068));
    LocalMux I__408 (
            .O(N__3078),
            .I(N__3065));
    InMux I__407 (
            .O(N__3075),
            .I(N__3060));
    InMux I__406 (
            .O(N__3074),
            .I(N__3060));
    Odrv12 I__405 (
            .O(N__3071),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ));
    Odrv4 I__404 (
            .O(N__3068),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ));
    Odrv4 I__403 (
            .O(N__3065),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ));
    LocalMux I__402 (
            .O(N__3060),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ));
    CascadeMux I__401 (
            .O(N__3051),
            .I(N__3047));
    InMux I__400 (
            .O(N__3050),
            .I(N__3044));
    InMux I__399 (
            .O(N__3047),
            .I(N__3041));
    LocalMux I__398 (
            .O(N__3044),
            .I(N__3036));
    LocalMux I__397 (
            .O(N__3041),
            .I(N__3036));
    Span4Mux_v I__396 (
            .O(N__3036),
            .I(N__3033));
    Odrv4 I__395 (
            .O(N__3033),
            .I(\U409_ADDRESS_DECODE.N_23 ));
    IoInMux I__394 (
            .O(N__3030),
            .I(N__3027));
    LocalMux I__393 (
            .O(N__3027),
            .I(N__3024));
    Span4Mux_s2_v I__392 (
            .O(N__3024),
            .I(N__3021));
    Span4Mux_v I__391 (
            .O(N__3021),
            .I(N__3018));
    Span4Mux_v I__390 (
            .O(N__3018),
            .I(N__3015));
    Sp12to4 I__389 (
            .O(N__3015),
            .I(N__3012));
    Odrv12 I__388 (
            .O(N__3012),
            .I(ROMENm_i));
    InMux I__387 (
            .O(N__3009),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__386 (
            .O(N__3006),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__385 (
            .O(N__3003),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__384 (
            .O(N__3000),
            .I(N__2997));
    LocalMux I__383 (
            .O(N__2997),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ));
    CascadeMux I__382 (
            .O(N__2994),
            .I(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0_cascade_ ));
    IoInMux I__381 (
            .O(N__2991),
            .I(N__2988));
    LocalMux I__380 (
            .O(N__2988),
            .I(N__2985));
    Span4Mux_s3_v I__379 (
            .O(N__2985),
            .I(N__2982));
    Span4Mux_v I__378 (
            .O(N__2982),
            .I(N__2979));
    Span4Mux_v I__377 (
            .O(N__2979),
            .I(N__2976));
    Odrv4 I__376 (
            .O(N__2976),
            .I(PORTSIZE_0_i));
    InMux I__375 (
            .O(N__2973),
            .I(N__2963));
    InMux I__374 (
            .O(N__2972),
            .I(N__2963));
    InMux I__373 (
            .O(N__2971),
            .I(N__2963));
    InMux I__372 (
            .O(N__2970),
            .I(N__2960));
    LocalMux I__371 (
            .O(N__2963),
            .I(N__2954));
    LocalMux I__370 (
            .O(N__2960),
            .I(N__2954));
    InMux I__369 (
            .O(N__2959),
            .I(N__2951));
    Span4Mux_v I__368 (
            .O(N__2954),
            .I(N__2945));
    LocalMux I__367 (
            .O(N__2951),
            .I(N__2945));
    InMux I__366 (
            .O(N__2950),
            .I(N__2942));
    Span4Mux_h I__365 (
            .O(N__2945),
            .I(N__2937));
    LocalMux I__364 (
            .O(N__2942),
            .I(N__2937));
    Sp12to4 I__363 (
            .O(N__2937),
            .I(N__2934));
    Span12Mux_v I__362 (
            .O(N__2934),
            .I(N__2931));
    Odrv12 I__361 (
            .O(N__2931),
            .I(A_c_22));
    InMux I__360 (
            .O(N__2928),
            .I(N__2925));
    LocalMux I__359 (
            .O(N__2925),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ));
    CascadeMux I__358 (
            .O(N__2922),
            .I(\U409_CIA.g0Z0Z_2_cascade_ ));
    InMux I__357 (
            .O(N__2919),
            .I(N__2916));
    LocalMux I__356 (
            .O(N__2916),
            .I(\U409_CIA.g0Z0Z_10 ));
    InMux I__355 (
            .O(N__2913),
            .I(N__2907));
    InMux I__354 (
            .O(N__2912),
            .I(N__2907));
    LocalMux I__353 (
            .O(N__2907),
            .I(N__2904));
    Odrv12 I__352 (
            .O(N__2904),
            .I(A_c_27));
    InMux I__351 (
            .O(N__2901),
            .I(N__2895));
    InMux I__350 (
            .O(N__2900),
            .I(N__2895));
    LocalMux I__349 (
            .O(N__2895),
            .I(N__2892));
    Odrv12 I__348 (
            .O(N__2892),
            .I(A_c_25));
    CascadeMux I__347 (
            .O(N__2889),
            .I(N__2885));
    InMux I__346 (
            .O(N__2888),
            .I(N__2880));
    InMux I__345 (
            .O(N__2885),
            .I(N__2880));
    LocalMux I__344 (
            .O(N__2880),
            .I(N__2877));
    Span4Mux_v I__343 (
            .O(N__2877),
            .I(N__2874));
    Span4Mux_v I__342 (
            .O(N__2874),
            .I(N__2871));
    Span4Mux_h I__341 (
            .O(N__2871),
            .I(N__2868));
    Odrv4 I__340 (
            .O(N__2868),
            .I(A_c_26));
    CascadeMux I__339 (
            .O(N__2865),
            .I(N__2862));
    InMux I__338 (
            .O(N__2862),
            .I(N__2856));
    InMux I__337 (
            .O(N__2861),
            .I(N__2856));
    LocalMux I__336 (
            .O(N__2856),
            .I(N__2853));
    Span4Mux_v I__335 (
            .O(N__2853),
            .I(N__2850));
    Span4Mux_v I__334 (
            .O(N__2850),
            .I(N__2847));
    Span4Mux_h I__333 (
            .O(N__2847),
            .I(N__2844));
    Odrv4 I__332 (
            .O(N__2844),
            .I(A_c_24));
    InMux I__331 (
            .O(N__2841),
            .I(N__2835));
    InMux I__330 (
            .O(N__2840),
            .I(N__2835));
    LocalMux I__329 (
            .O(N__2835),
            .I(N__2832));
    Span4Mux_v I__328 (
            .O(N__2832),
            .I(N__2829));
    Sp12to4 I__327 (
            .O(N__2829),
            .I(N__2826));
    Odrv12 I__326 (
            .O(N__2826),
            .I(A_c_31));
    InMux I__325 (
            .O(N__2823),
            .I(N__2817));
    InMux I__324 (
            .O(N__2822),
            .I(N__2817));
    LocalMux I__323 (
            .O(N__2817),
            .I(N__2814));
    Sp12to4 I__322 (
            .O(N__2814),
            .I(N__2811));
    Span12Mux_v I__321 (
            .O(N__2811),
            .I(N__2808));
    Odrv12 I__320 (
            .O(N__2808),
            .I(A_c_29));
    InMux I__319 (
            .O(N__2805),
            .I(N__2802));
    LocalMux I__318 (
            .O(N__2802),
            .I(N__2798));
    CascadeMux I__317 (
            .O(N__2801),
            .I(N__2795));
    Span4Mux_v I__316 (
            .O(N__2798),
            .I(N__2792));
    InMux I__315 (
            .O(N__2795),
            .I(N__2789));
    Span4Mux_h I__314 (
            .O(N__2792),
            .I(N__2784));
    LocalMux I__313 (
            .O(N__2789),
            .I(N__2784));
    Span4Mux_v I__312 (
            .O(N__2784),
            .I(N__2781));
    Span4Mux_h I__311 (
            .O(N__2781),
            .I(N__2778));
    Odrv4 I__310 (
            .O(N__2778),
            .I(A_c_30));
    InMux I__309 (
            .O(N__2775),
            .I(N__2771));
    InMux I__308 (
            .O(N__2774),
            .I(N__2768));
    LocalMux I__307 (
            .O(N__2771),
            .I(N__2763));
    LocalMux I__306 (
            .O(N__2768),
            .I(N__2763));
    Span4Mux_h I__305 (
            .O(N__2763),
            .I(N__2760));
    Span4Mux_v I__304 (
            .O(N__2760),
            .I(N__2757));
    Span4Mux_v I__303 (
            .O(N__2757),
            .I(N__2754));
    Odrv4 I__302 (
            .O(N__2754),
            .I(A_c_28));
    InMux I__301 (
            .O(N__2751),
            .I(N__2745));
    InMux I__300 (
            .O(N__2750),
            .I(N__2745));
    LocalMux I__299 (
            .O(N__2745),
            .I(N__2742));
    Span4Mux_v I__298 (
            .O(N__2742),
            .I(N__2739));
    Span4Mux_h I__297 (
            .O(N__2739),
            .I(N__2736));
    Span4Mux_v I__296 (
            .O(N__2736),
            .I(N__2733));
    Span4Mux_v I__295 (
            .O(N__2733),
            .I(N__2730));
    Odrv4 I__294 (
            .O(N__2730),
            .I(A_c_18));
    CascadeMux I__293 (
            .O(N__2727),
            .I(N__2723));
    CascadeMux I__292 (
            .O(N__2726),
            .I(N__2720));
    InMux I__291 (
            .O(N__2723),
            .I(N__2717));
    InMux I__290 (
            .O(N__2720),
            .I(N__2714));
    LocalMux I__289 (
            .O(N__2717),
            .I(N__2709));
    LocalMux I__288 (
            .O(N__2714),
            .I(N__2709));
    Span4Mux_h I__287 (
            .O(N__2709),
            .I(N__2706));
    Sp12to4 I__286 (
            .O(N__2706),
            .I(N__2703));
    Span12Mux_v I__285 (
            .O(N__2703),
            .I(N__2700));
    Odrv12 I__284 (
            .O(N__2700),
            .I(A_c_16));
    InMux I__283 (
            .O(N__2697),
            .I(N__2691));
    InMux I__282 (
            .O(N__2696),
            .I(N__2691));
    LocalMux I__281 (
            .O(N__2691),
            .I(N__2688));
    Sp12to4 I__280 (
            .O(N__2688),
            .I(N__2685));
    Span12Mux_v I__279 (
            .O(N__2685),
            .I(N__2682));
    Odrv12 I__278 (
            .O(N__2682),
            .I(A_c_17));
    CascadeMux I__277 (
            .O(N__2679),
            .I(\U409_CIA.g0Z0Z_11_cascade_ ));
    InMux I__276 (
            .O(N__2676),
            .I(N__2673));
    LocalMux I__275 (
            .O(N__2673),
            .I(N__2670));
    Odrv4 I__274 (
            .O(N__2670),
            .I(\U409_CIA.g0Z0Z_8 ));
    InMux I__273 (
            .O(N__2667),
            .I(N__2664));
    LocalMux I__272 (
            .O(N__2664),
            .I(N__2659));
    InMux I__271 (
            .O(N__2663),
            .I(N__2654));
    InMux I__270 (
            .O(N__2662),
            .I(N__2654));
    Span4Mux_v I__269 (
            .O(N__2659),
            .I(N__2651));
    LocalMux I__268 (
            .O(N__2654),
            .I(N__2648));
    Sp12to4 I__267 (
            .O(N__2651),
            .I(N__2645));
    Span4Mux_h I__266 (
            .O(N__2648),
            .I(N__2642));
    Span12Mux_s3_h I__265 (
            .O(N__2645),
            .I(N__2637));
    Sp12to4 I__264 (
            .O(N__2642),
            .I(N__2637));
    Span12Mux_v I__263 (
            .O(N__2637),
            .I(N__2634));
    Odrv12 I__262 (
            .O(N__2634),
            .I(A_c_19));
    CascadeMux I__261 (
            .O(N__2631),
            .I(\U409_ADDRESS_DECODE.ROMEN_0_a2_0Z0Z_2_cascade_ ));
    InMux I__260 (
            .O(N__2628),
            .I(N__2625));
    LocalMux I__259 (
            .O(N__2625),
            .I(\U409_ADDRESS_DECODE.N_58 ));
    InMux I__258 (
            .O(N__2622),
            .I(N__2618));
    InMux I__257 (
            .O(N__2621),
            .I(N__2615));
    LocalMux I__256 (
            .O(N__2618),
            .I(N__2610));
    LocalMux I__255 (
            .O(N__2615),
            .I(N__2610));
    Span4Mux_v I__254 (
            .O(N__2610),
            .I(N__2607));
    Sp12to4 I__253 (
            .O(N__2607),
            .I(N__2604));
    Span12Mux_h I__252 (
            .O(N__2604),
            .I(N__2601));
    Span12Mux_v I__251 (
            .O(N__2601),
            .I(N__2598));
    Span12Mux_h I__250 (
            .O(N__2598),
            .I(N__2595));
    Odrv12 I__249 (
            .O(N__2595),
            .I(OVL_c));
    CascadeMux I__248 (
            .O(N__2592),
            .I(N__2589));
    InMux I__247 (
            .O(N__2589),
            .I(N__2583));
    InMux I__246 (
            .O(N__2588),
            .I(N__2583));
    LocalMux I__245 (
            .O(N__2583),
            .I(N__2580));
    Odrv12 I__244 (
            .O(N__2580),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEm_6 ));
    CascadeMux I__243 (
            .O(N__2577),
            .I(N__2572));
    InMux I__242 (
            .O(N__2576),
            .I(N__2569));
    InMux I__241 (
            .O(N__2575),
            .I(N__2564));
    InMux I__240 (
            .O(N__2572),
            .I(N__2564));
    LocalMux I__239 (
            .O(N__2569),
            .I(N__2561));
    LocalMux I__238 (
            .O(N__2564),
            .I(N__2558));
    Span4Mux_v I__237 (
            .O(N__2561),
            .I(N__2552));
    Span4Mux_v I__236 (
            .O(N__2558),
            .I(N__2552));
    InMux I__235 (
            .O(N__2557),
            .I(N__2549));
    Sp12to4 I__234 (
            .O(N__2552),
            .I(N__2544));
    LocalMux I__233 (
            .O(N__2549),
            .I(N__2544));
    Odrv12 I__232 (
            .O(N__2544),
            .I(A_c_20));
    ClkMux I__231 (
            .O(N__2541),
            .I(N__2505));
    ClkMux I__230 (
            .O(N__2540),
            .I(N__2505));
    ClkMux I__229 (
            .O(N__2539),
            .I(N__2505));
    ClkMux I__228 (
            .O(N__2538),
            .I(N__2505));
    ClkMux I__227 (
            .O(N__2537),
            .I(N__2505));
    ClkMux I__226 (
            .O(N__2536),
            .I(N__2505));
    ClkMux I__225 (
            .O(N__2535),
            .I(N__2505));
    ClkMux I__224 (
            .O(N__2534),
            .I(N__2505));
    ClkMux I__223 (
            .O(N__2533),
            .I(N__2505));
    ClkMux I__222 (
            .O(N__2532),
            .I(N__2505));
    ClkMux I__221 (
            .O(N__2531),
            .I(N__2505));
    ClkMux I__220 (
            .O(N__2530),
            .I(N__2505));
    GlobalMux I__219 (
            .O(N__2505),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .I(N__2541));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .I(N__2540));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .I(N__2539));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .I(N__2534));
    INV \INVU409_TRANSFER_ACK.TACK_EN_iC  (
            .O(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .I(N__2537));
    INV \INVU409_TRANSFER_ACK.TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .I(N__2535));
    INV \INVU409_TRANSFER_ACK.CIA_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .I(N__2533));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__2532));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .I(N__2530));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .I(N__2538));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_EN_nesrC  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_EN_nesrC_net ),
            .I(N__2536));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .I(N__2531));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_10_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_5_0_));
    defparam IN_MUX_bfv_10_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_6_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_10_6_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_6_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_9_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_9_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_1_9_0  (
            .in0(N__2662),
            .in1(N__2750),
            .in2(N__2726),
            .in3(N__2696),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEm_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_11_LC_1_9_1 .C_ON=1'b0;
    defparam \U409_CIA.g0_11_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_11_LC_1_9_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.g0_11_LC_1_9_1  (
            .in0(N__2751),
            .in1(N__3270),
            .in2(N__2727),
            .in3(N__2663),
            .lcout(),
            .ltout(\U409_CIA.g0Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_14_LC_1_9_2 .C_ON=1'b0;
    defparam \U409_CIA.g0_14_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_14_LC_1_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.g0_14_LC_1_9_2  (
            .in0(N__2576),
            .in1(N__2697),
            .in2(N__2679),
            .in3(N__2676),
            .lcout(\U409_CIA.g0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_8_LC_1_12_1 .C_ON=1'b0;
    defparam \U409_CIA.g0_8_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_8_LC_1_12_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_CIA.g0_8_LC_1_12_1  (
            .in0(N__2973),
            .in1(N__3374),
            .in2(_gnd_net_),
            .in3(N__2805),
            .lcout(\U409_CIA.g0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_0_2_LC_1_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_0_2_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_0_2_LC_1_12_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a2_0_2_LC_1_12_2  (
            .in0(N__2557),
            .in1(N__2971),
            .in2(_gnd_net_),
            .in3(N__3262),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.ROMEN_0_a2_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_o2_LC_1_12_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_o2_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_o2_LC_1_12_3 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_o2_LC_1_12_3  (
            .in0(N__2667),
            .in1(N__3373),
            .in2(N__2631),
            .in3(N__2628),
            .lcout(\U409_ADDRESS_DECODE.N_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_1_LC_1_12_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_1_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_1_LC_1_12_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a2_1_LC_1_12_6  (
            .in0(N__2621),
            .in1(N__2972),
            .in2(N__3375),
            .in3(N__3263),
            .lcout(\U409_ADDRESS_DECODE.N_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_2_LC_1_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_2_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_2_LC_1_13_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nRAMSPACE_2_LC_1_13_4  (
            .in0(N__2970),
            .in1(N__3144),
            .in2(N__3100),
            .in3(N__2622),
            .lcout(\U409_ADDRESS_DECODE.un1_nRAMSPACEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_1_14_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_1_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_1_14_4  (
            .in0(N__3224),
            .in1(N__3350),
            .in2(N__2577),
            .in3(N__2588),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_1_14_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_1_14_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_1_14_7  (
            .in0(N__2959),
            .in1(N__3351),
            .in2(N__2592),
            .in3(N__2575),
            .lcout(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_1_15_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_1_15_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_1_15_1  (
            .in0(N__3131),
            .in1(N__3261),
            .in2(N__3089),
            .in3(N__3191),
            .lcout(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0 ),
            .ltout(\U409_ADDRESS_DECODE.un1_nREGSPACEZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_1_15_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_1_15_2 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_1_15_2  (
            .in0(N__3000),
            .in1(_gnd_net_),
            .in2(N__2994),
            .in3(N__2928),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_15_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_15_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_1_15_6  (
            .in0(N__2950),
            .in1(N__3130),
            .in2(N__5865),
            .in3(N__3074),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_2_LC_1_16_1 .C_ON=1'b0;
    defparam \U409_CIA.g0_2_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_2_LC_1_16_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_CIA.g0_2_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__2823),
            .in2(_gnd_net_),
            .in3(N__5874),
            .lcout(),
            .ltout(\U409_CIA.g0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_13_LC_1_16_2 .C_ON=1'b0;
    defparam \U409_CIA.g0_13_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_13_LC_1_16_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_CIA.g0_13_LC_1_16_2  (
            .in0(N__2919),
            .in1(N__2841),
            .in2(N__2922),
            .in3(N__2775),
            .lcout(\U409_CIA.g0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.g0_10_LC_1_16_3 .C_ON=1'b0;
    defparam \U409_CIA.g0_10_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.g0_10_LC_1_16_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.g0_10_LC_1_16_3  (
            .in0(N__2901),
            .in1(N__2913),
            .in2(N__2865),
            .in3(N__2888),
            .lcout(\U409_CIA.g0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_16_4  (
            .in0(N__2912),
            .in1(N__2900),
            .in2(N__2889),
            .in3(N__2861),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_16_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_16_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_16_7  (
            .in0(N__2840),
            .in1(N__2822),
            .in2(N__2801),
            .in3(N__2774),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_2_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_2_12_2 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_2_12_2  (
            .in0(N__3369),
            .in1(N__3269),
            .in2(_gnd_net_),
            .in3(N__3311),
            .lcout(U409_ADDRESS_DECODE_un1_nRAMSPACE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_2_15_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_2_15_7 .LUT_INIT=16'b0000000011101111;
    LogicCell40 \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_2_15_7  (
            .in0(N__3267),
            .in1(N__3368),
            .in2(N__3318),
            .in3(N__3300),
            .lcout(nBUFEN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_3_15_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_3_15_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_3_15_4  (
            .in0(N__3154),
            .in1(N__3268),
            .in2(N__3201),
            .in3(N__3101),
            .lcout(U409_ADDRESS_DECODE_un1_nREGSPACE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_5_13_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_5_13_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_5_13_7  (
            .in0(N__3105),
            .in1(N__3156),
            .in2(N__3051),
            .in3(N__5866),
            .lcout(ROMENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_5_16_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_5_16_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMENm_i_LC_5_16_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_ADDRESS_DECODE.ROMENm_i_LC_5_16_6  (
            .in0(N__3155),
            .in1(N__3099),
            .in2(N__5873),
            .in3(N__3050),
            .lcout(ROMENm_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_7_6_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_7_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__3547),
            .in2(N__3591),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_6_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_7_6_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_7_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__3435),
            .in2(_gnd_net_),
            .in3(N__3009),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__3525),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_7_6_2 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_7_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__3630),
            .in2(_gnd_net_),
            .in3(N__3006),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_7_6_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_7_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__3457),
            .in2(_gnd_net_),
            .in3(N__3003),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__3525),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_7_6_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_7_6_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(N__3415),
            .in2(_gnd_net_),
            .in3(N__3483),
            .lcout(),
            .ltout(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_7_6_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_7_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_7_6_5 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_7_6_5  (
            .in0(N__3632),
            .in1(N__3467),
            .in2(N__3480),
            .in3(N__3584),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3525),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_7_6_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_7_6_6 .LUT_INIT=16'b0011001101001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_7_6_6  (
            .in0(N__3585),
            .in1(N__3477),
            .in2(N__3471),
            .in3(N__3631),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3525),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_7_6_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_7_6_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_7_6_7  (
            .in0(N__3548),
            .in1(N__3458),
            .in2(N__3420),
            .in3(N__3436),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_7_7_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_7_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__3590),
            .in2(_gnd_net_),
            .in3(N__3552),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3523),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_HOLD_LC_7_8_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_HOLD_LC_7_8_0 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U409_CIA.CIA_HOLD_LC_7_8_0  (
            .in0(N__4372),
            .in1(N__4291),
            .in2(N__4333),
            .in3(N__4255),
            .lcout(\U409_CIA.CIA_HOLDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3522),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_8_6_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_8_6_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_8_6_0  (
            .in0(N__3411),
            .in1(N__3437),
            .in2(_gnd_net_),
            .in3(N__3456),
            .lcout(\U409_CIA.CLKCIA8_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_8_6_1 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_8_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3588),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3524),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_1_LC_8_6_2 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_1_LC_8_6_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CLKCIA_RNO_1_LC_8_6_2  (
            .in0(N__3459),
            .in1(N__3438),
            .in2(N__3419),
            .in3(N__3635),
            .lcout(\U409_CIA.CLKCIA6_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_8_6_3 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_8_6_3 .LUT_INIT=16'b0100010000100010;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_8_6_3  (
            .in0(N__3634),
            .in1(N__3587),
            .in2(_gnd_net_),
            .in3(N__3550),
            .lcout(),
            .ltout(\U409_CIA.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_8_6_4 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_8_6_4 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \U409_CIA.VMA_LC_8_6_4  (
            .in0(N__4285),
            .in1(N__3636),
            .in2(N__3639),
            .in3(N__3606),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3524),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_2_LC_8_6_5 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_2_LC_8_6_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_CIA.CLKCIA_RNO_2_LC_8_6_5  (
            .in0(N__3633),
            .in1(N__3586),
            .in2(_gnd_net_),
            .in3(N__3549),
            .lcout(),
            .ltout(\U409_CIA.N_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_RNO_0_LC_8_6_6 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLKCIA_RNO_0_LC_8_6_6 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \U409_CIA.CLKCIA_RNO_0_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(N__4219),
            .in2(N__3609),
            .in3(N__3605),
            .lcout(),
            .ltout(\U409_CIA.CLKCIAZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLKCIA_LC_8_6_7 .C_ON=1'b0;
    defparam \U409_CIA.CLKCIA_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLKCIA_LC_8_6_7 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \U409_CIA.CLKCIA_LC_8_6_7  (
            .in0(N__3597),
            .in1(N__3589),
            .in2(N__3555),
            .in3(N__3551),
            .lcout(CLKCIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3524),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_8_7_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_8_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__3871),
            .in2(_gnd_net_),
            .in3(N__3891),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4837),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_8_7_1 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_8_7_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \U409_TICK.TICK60_LC_8_7_1  (
            .in0(N__3741),
            .in1(N__3666),
            .in2(N__3717),
            .in3(N__3494),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4837),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_8_7_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_8_7_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_8_7_2  (
            .in0(N__3664),
            .in1(N__3744),
            .in2(N__3712),
            .in3(N__4086),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4837),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_8_7_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_8_7_3 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_8_7_3  (
            .in0(N__3740),
            .in1(N__3665),
            .in2(N__3765),
            .in3(N__3703),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4837),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_8_7_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_8_7_4 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_8_7_4  (
            .in0(N__3699),
            .in1(N__3742),
            .in2(N__3672),
            .in3(N__3872),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4837),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_8_7_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_8_7_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_8_7_5  (
            .in0(N__4077),
            .in1(N__4098),
            .in2(N__3780),
            .in3(N__3993),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_8_7_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_8_7_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_8_7_6  (
            .in0(N__3663),
            .in1(N__3743),
            .in2(N__3753),
            .in3(N__3804),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4837),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_8_8_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_8_8_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_8_8_0  (
            .in0(N__3738),
            .in1(N__3671),
            .in2(N__3713),
            .in3(N__4065),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4839),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_8_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_8_8_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_8_8_2  (
            .in0(N__4113),
            .in1(N__4008),
            .in2(N__4056),
            .in3(N__4176),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(\U409_TICK.TICK603_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_8_8_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_8_8_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_8_8_3  (
            .in0(N__3704),
            .in1(N__3739),
            .in2(N__3750),
            .in3(N__4164),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4839),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_8_8_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_8_8_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_8_8_4  (
            .in0(N__3795),
            .in1(N__3816),
            .in2(_gnd_net_),
            .in3(N__3870),
            .lcout(),
            .ltout(\U409_TICK.TICK603_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_8_8_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_8_8_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_8_8_5  (
            .in0(N__3972),
            .in1(N__4038),
            .in2(N__3747),
            .in3(N__3831),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_8_8_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_8_8_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_8_8_6  (
            .in0(N__3705),
            .in1(N__3670),
            .in2(N__3642),
            .in3(N__3981),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4839),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_8_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_8_8_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_8_8_7  (
            .in0(N__4023),
            .in1(N__3890),
            .in2(N__3849),
            .in3(N__4151),
            .lcout(\U409_TICK.TICK603_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_9_4_3  (
            .in0(N__4398),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3966),
            .lcout(U409_ADDRESS_DECODE_un1_nCIACS1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_6_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_6_1 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_9_6_1  (
            .in0(N__3927),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4394),
            .lcout(U409_ADDRESS_DECODE_un1_nCIACS0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_9_7_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_9_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__3889),
            .in2(N__3873),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_9_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_9_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__3845),
            .in2(_gnd_net_),
            .in3(N__3834),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__4836),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_9_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_9_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__3830),
            .in2(_gnd_net_),
            .in3(N__3819),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__4836),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_9_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_9_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(N__3815),
            .in2(_gnd_net_),
            .in3(N__3798),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_9_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_9_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__3794),
            .in2(_gnd_net_),
            .in3(N__3783),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__4836),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_9_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_9_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__3776),
            .in2(_gnd_net_),
            .in3(N__3756),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_9_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_9_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(N__4112),
            .in2(_gnd_net_),
            .in3(N__4101),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__4836),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_9_7_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_9_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(N__4097),
            .in2(_gnd_net_),
            .in3(N__4080),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_9_8_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_9_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__4076),
            .in2(_gnd_net_),
            .in3(N__4059),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_9_8_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_9_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__4052),
            .in2(_gnd_net_),
            .in3(N__4041),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__4838),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_9_8_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_9_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__4037),
            .in2(_gnd_net_),
            .in3(N__4026),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__4838),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_9_8_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_9_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__4022),
            .in2(_gnd_net_),
            .in3(N__4011),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__4838),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_9_8_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_9_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__4007),
            .in2(_gnd_net_),
            .in3(N__3996),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__4838),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_9_8_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_9_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__3992),
            .in2(_gnd_net_),
            .in3(N__3975),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_9_8_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_9_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__4175),
            .in2(_gnd_net_),
            .in3(N__4158),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_9_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_9_8_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__4152),
            .in2(_gnd_net_),
            .in3(N__4155),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4838),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_9_11_3.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_9_11_3.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_9_11_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_9_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5855),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNO_LC_9_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNO_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNO_LC_9_12_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNO_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__5023),
            .in2(_gnd_net_),
            .in3(N__4125),
            .lcout(\U409_TRANSFER_ACK.N_22_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI8GRM5_2_LC_9_13_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI8GRM5_2_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI8GRM5_2_LC_9_13_4 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI8GRM5_2_LC_9_13_4  (
            .in0(N__5471),
            .in1(N__5432),
            .in2(N__4140),
            .in3(N__4526),
            .lcout(\U409_TRANSFER_ACK.N_24 ),
            .ltout(\U409_TRANSFER_ACK.N_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNO_0_LC_9_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNO_0_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNO_0_LC_9_13_5 .LUT_INIT=16'b1101110111111100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNO_0_LC_9_13_5  (
            .in0(N__4527),
            .in1(N__4503),
            .in2(N__4128),
            .in3(N__4479),
            .lcout(\U409_TRANSFER_ACK.N_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_10_5_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_10_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_10_5_0  (
            .in0(_gnd_net_),
            .in1(N__4659),
            .in2(N__4730),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_5_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_10_5_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_10_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_10_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_10_5_1  (
            .in0(_gnd_net_),
            .in1(N__4754),
            .in2(_gnd_net_),
            .in3(N__4119),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__4833),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_10_5_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_10_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_10_5_2  (
            .in0(_gnd_net_),
            .in1(N__4676),
            .in2(_gnd_net_),
            .in3(N__4116),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__4833),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_10_5_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_10_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_10_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_10_5_3  (
            .in0(_gnd_net_),
            .in1(N__4430),
            .in2(_gnd_net_),
            .in3(N__4203),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__4833),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_10_5_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_10_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_10_5_4  (
            .in0(_gnd_net_),
            .in1(N__4688),
            .in2(_gnd_net_),
            .in3(N__4200),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_10_5_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_10_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_10_5_5  (
            .in0(_gnd_net_),
            .in1(N__4454),
            .in2(_gnd_net_),
            .in3(N__4197),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_10_5_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_10_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_10_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_10_5_6  (
            .in0(_gnd_net_),
            .in1(N__4442),
            .in2(_gnd_net_),
            .in3(N__4194),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__4833),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_10_5_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_10_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_10_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_10_5_7  (
            .in0(_gnd_net_),
            .in1(N__4766),
            .in2(_gnd_net_),
            .in3(N__4191),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__4833),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_10_6_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_10_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_10_6_0  (
            .in0(_gnd_net_),
            .in1(N__4850),
            .in2(_gnd_net_),
            .in3(N__4188),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_10_6_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_10_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_10_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_10_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_10_6_1  (
            .in0(_gnd_net_),
            .in1(N__4619),
            .in2(_gnd_net_),
            .in3(N__4185),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__4835),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_10_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_10_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(N__4595),
            .in2(_gnd_net_),
            .in3(N__4182),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_10_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_10_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_10_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_10_6_3  (
            .in0(_gnd_net_),
            .in1(N__4634),
            .in2(_gnd_net_),
            .in3(N__4179),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__4835),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_10_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_10_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_10_6_4  (
            .in0(_gnd_net_),
            .in1(N__4550),
            .in2(_gnd_net_),
            .in3(N__4410),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_10_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_10_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_10_6_5  (
            .in0(_gnd_net_),
            .in1(N__4574),
            .in2(_gnd_net_),
            .in3(N__4407),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_10_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_10_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_10_6_6  (
            .in0(_gnd_net_),
            .in1(N__4979),
            .in2(_gnd_net_),
            .in3(N__4404),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_10_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_10_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_10_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_10_6_7  (
            .in0(_gnd_net_),
            .in1(N__4743),
            .in2(_gnd_net_),
            .in3(N__4401),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4835),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_10_8_3 .C_ON=1'b0;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_10_8_3 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_10_8_3  (
            .in0(N__4298),
            .in1(N__4380),
            .in2(N__4347),
            .in3(N__4262),
            .lcout(CIA_ENABLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_9_0 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_10_9_0  (
            .in0(N__4373),
            .in1(N__4340),
            .in2(N__4302),
            .in3(N__4266),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__5051));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_10_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_10_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_10_9_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_10_9_2  (
            .in0(N__4232),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__5051));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_10_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_10_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4806),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__5051));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_10_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_10_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_10_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5214),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__5051));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_LC_10_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_LC_10_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4530),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_EN_nesrC_net ),
            .ce(N__4539),
            .sr(N__5044));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_10_13_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_10_13_1 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_10_13_1  (
            .in0(N__4505),
            .in1(N__4481),
            .in2(_gnd_net_),
            .in3(N__4529),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__5055));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_10_13_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_10_13_3 .LUT_INIT=16'b0010001001100110;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_10_13_3  (
            .in0(N__4504),
            .in1(N__4480),
            .in2(_gnd_net_),
            .in3(N__4528),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__5055));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_10_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_10_13_5 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_10_13_5  (
            .in0(N__4506),
            .in1(N__4488),
            .in2(_gnd_net_),
            .in3(N__4482),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__5055));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_11_5_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_11_5_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_11_5_0  (
            .in0(N__4551),
            .in1(N__4851),
            .in2(N__4599),
            .in3(N__4455),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_11_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_11_5_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_11_5_1  (
            .in0(N__4875),
            .in1(N__4934),
            .in2(N__4464),
            .in3(N__4461),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4832),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_11_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_11_5_2 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_11_5_2  (
            .in0(N__4961),
            .in1(N__4930),
            .in2(N__4665),
            .in3(N__4874),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4832),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_11_5_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_11_5_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_11_5_3  (
            .in0(N__4980),
            .in1(N__4443),
            .in2(N__4578),
            .in3(N__4431),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_11_5_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_11_5_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_11_5_4  (
            .in0(N__4962),
            .in1(N__4931),
            .in2(N__4419),
            .in3(N__4416),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4832),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_5_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_5_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_11_5_5  (
            .in0(N__4767),
            .in1(N__4755),
            .in2(N__4731),
            .in3(N__4742),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_11_5_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_11_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_11_5_6  (
            .in0(N__4664),
            .in1(N__4729),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4832),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_11_5_7 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_11_5_7 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \U409_TICK.TICK50_LC_11_5_7  (
            .in0(N__4876),
            .in1(N__4963),
            .in2(N__4706),
            .in3(N__4935),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4832),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_11_6_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_11_6_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_11_6_0  (
            .in0(N__4689),
            .in1(N__4677),
            .in2(_gnd_net_),
            .in3(N__4660),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_11_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_11_6_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_11_6_1  (
            .in0(N__4641),
            .in1(N__4635),
            .in2(N__4623),
            .in3(N__4620),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_11_6_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_11_6_2 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_11_6_2  (
            .in0(N__4608),
            .in1(N__4877),
            .in2(N__4602),
            .in3(N__4964),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4834),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_11_6_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_11_6_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_11_6_3  (
            .in0(N__4879),
            .in1(N__4966),
            .in2(N__4932),
            .in3(N__4584),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4834),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_11_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_11_6_4 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_11_6_4  (
            .in0(N__4965),
            .in1(N__4923),
            .in2(N__4563),
            .in3(N__4878),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4834),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_11_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_11_6_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_11_6_5  (
            .in0(N__4880),
            .in1(N__4967),
            .in2(N__4933),
            .in3(N__4986),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4834),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_11_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_11_6_6 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_11_6_6  (
            .in0(N__4968),
            .in1(N__4924),
            .in2(N__4893),
            .in3(N__4881),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4834),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_0_LC_11_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_0_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_0_LC_11_9_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_0_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__5179),
            .in2(_gnd_net_),
            .in3(N__5099),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_2_LC_11_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_2_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_2_LC_11_9_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_2_LC_11_9_2  (
            .in0(N__5160),
            .in1(N__5211),
            .in2(N__4809),
            .in3(N__5441),
            .lcout(\U409_TRANSFER_ACK.N_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m12_0_a4_LC_11_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m12_0_a4_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m12_0_a4_LC_11_9_3 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m12_0_a4_LC_11_9_3  (
            .in0(N__5210),
            .in1(N__5183),
            .in2(N__5159),
            .in3(N__5101),
            .lcout(\U409_TRANSFER_ACK.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_1_LC_11_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_1_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_1_LC_11_9_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_1_LC_11_9_4  (
            .in0(N__5100),
            .in1(N__4788),
            .in2(N__5187),
            .in3(N__4805),
            .lcout(\U409_TRANSFER_ACK.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_o2_0_LC_11_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_o2_0_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_o2_0_LC_11_9_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_o2_0_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__4804),
            .in2(_gnd_net_),
            .in3(N__4787),
            .lcout(\U409_TRANSFER_ACK.N_29 ),
            .ltout(\U409_TRANSFER_ACK.N_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_9_6 .LUT_INIT=16'b0010000000100010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_9_6  (
            .in0(N__5833),
            .in1(N__4776),
            .in2(N__4770),
            .in3(N__5082),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_LC_11_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_LC_11_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__5185),
            .in2(_gnd_net_),
            .in3(N__5102),
            .lcout(\U409_TRANSFER_ACK.N_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_10_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_10_2  (
            .in0(N__5433),
            .in1(N__5212),
            .in2(N__5157),
            .in3(N__5186),
            .lcout(\U409_TRANSFER_ACK.N_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_0_LC_11_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_0_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_0_LC_11_10_4 .LUT_INIT=16'b0001001100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a4_0_LC_11_10_4  (
            .in0(N__5213),
            .in1(N__5184),
            .in2(N__5158),
            .in3(N__5103),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.N_52_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_1_LC_11_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_1_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_1_LC_11_10_5 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_1_LC_11_10_5  (
            .in0(N__5077),
            .in1(N__5127),
            .in2(N__5121),
            .in3(N__5118),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.m9_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_10_6 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_10_6  (
            .in0(N__5834),
            .in1(_gnd_net_),
            .in2(N__5112),
            .in3(N__5109),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_11_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_11_0  (
            .in0(N__5078),
            .in1(N__5061),
            .in2(_gnd_net_),
            .in3(N__5001),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__5043));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_11_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_11_12_0 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_11_12_0  (
            .in0(N__5330),
            .in1(N__5840),
            .in2(_gnd_net_),
            .in3(N__5314),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNIUBID_LC_11_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNIUBID_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNIUBID_LC_11_12_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_nesr_RNIUBID_LC_11_12_2  (
            .in0(N__5007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5000),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNILJA71_LC_11_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNILJA71_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNILJA71_LC_11_12_3 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNILJA71_LC_11_12_3  (
            .in0(N__5315),
            .in1(N__5329),
            .in2(N__4989),
            .in3(N__5234),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_12_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_12_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5334),
            .in3(N__5838),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_12_5  (
            .in0(N__5839),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5331),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_12_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_12_6 .LUT_INIT=16'b0010001011101010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_11_12_6  (
            .in0(N__5285),
            .in1(N__5841),
            .in2(N__5319),
            .in3(N__5274),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_11_13_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_11_13_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_LC_11_13_1  (
            .in0(N__5842),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5273),
            .lcout(TACK_EN_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .ce(N__5262),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_13_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_13_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_13_7 .LUT_INIT=16'b0010001011111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_13_7  (
            .in0(N__5235),
            .in1(N__5223),
            .in2(_gnd_net_),
            .in3(N__5993),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .ce(),
            .sr(N__5754));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNO_0_LC_13_13_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNO_0_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNO_0_LC_13_13_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNO_0_LC_13_13_2  (
            .in0(N__5514),
            .in1(N__5346),
            .in2(N__5364),
            .in3(N__5618),
            .lcout(\U409_TRANSFER_ACK.N_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIT7KM1_4_LC_13_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIT7KM1_4_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIT7KM1_4_LC_13_13_6 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIT7KM1_4_LC_13_13_6  (
            .in0(N__5513),
            .in1(N__6034),
            .in2(N__5619),
            .in3(N__5552),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CJV2_7_LC_13_13_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CJV2_7_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CJV2_7_LC_13_13_7 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CJV2_7_LC_13_13_7  (
            .in0(N__5923),
            .in1(N__5583),
            .in2(N__5217),
            .in3(N__5652),
            .lcout(\U409_TRANSFER_ACK.N_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_13_14_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_13_14_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_13_14_0 .LUT_INIT=16'b1101110011101100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_13_14_0  (
            .in0(N__5681),
            .in1(N__5951),
            .in2(N__6003),
            .in3(N__5666),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5745));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_0_LC_13_14_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_0_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_0_LC_13_14_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_0_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(N__5680),
            .in2(_gnd_net_),
            .in3(N__5580),
            .lcout(\U409_TRANSFER_ACK.N_41_4 ),
            .ltout(\U409_TRANSFER_ACK.N_41_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIGDB12_2_LC_13_14_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIGDB12_2_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIGDB12_2_LC_13_14_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIGDB12_2_LC_13_14_2  (
            .in0(N__5478),
            .in1(N__5617),
            .in2(N__5451),
            .in3(N__5515),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a4_0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI772Q3_2_LC_13_14_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI772Q3_2_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI772Q3_2_LC_13_14_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI772Q3_2_LC_13_14_3  (
            .in0(N__5363),
            .in1(_gnd_net_),
            .in2(N__5448),
            .in3(N__5437),
            .lcout(\U409_TRANSFER_ACK.N_44 ),
            .ltout(\U409_TRANSFER_ACK.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_13_14_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_13_14_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_13_14_4 .LUT_INIT=16'b0000010000001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_13_14_4  (
            .in0(N__5581),
            .in1(N__6001),
            .in2(N__5367),
            .in3(N__5562),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5745));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_13_14_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_13_14_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_13_14_5 .LUT_INIT=16'b0000010000001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_13_14_5  (
            .in0(N__5516),
            .in1(N__5997),
            .in2(N__5960),
            .in3(N__5487),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5745));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_13_14_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_13_14_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_13_14_6 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_13_14_6  (
            .in0(N__5998),
            .in1(N__5955),
            .in2(N__6039),
            .in3(N__6012),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5745));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIU8KM1_7_LC_14_13_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIU8KM1_7_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIU8KM1_7_LC_14_13_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIU8KM1_7_LC_14_13_4  (
            .in0(N__5550),
            .in1(N__5649),
            .in2(N__5924),
            .in3(N__6033),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_2_LC_14_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_2_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_2_LC_14_13_5 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_2_LC_14_13_5  (
            .in0(N__5612),
            .in1(N__5512),
            .in2(N__5349),
            .in3(N__5345),
            .lcout(\U409_TRANSFER_ACK.N_41_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_14_13_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_14_13_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_14_13_6 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_14_13_6  (
            .in0(N__5999),
            .in1(N__5956),
            .in2(N__5631),
            .in3(N__5650),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__5750));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_14_13_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_14_13_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_14_13_7 .LUT_INIT=16'b0000010000001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_14_13_7  (
            .in0(N__5553),
            .in1(N__6000),
            .in2(N__5961),
            .in3(N__5529),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__5750));
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_c_LC_14_14_0 .C_ON=1'b1;
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_c_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_c_LC_14_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_c_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__5682),
            .in2(N__5667),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_THRU_LUT4_0_LC_14_14_1 .C_ON=1'b1;
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_THRU_LUT4_0_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_THRU_LUT4_0_LC_14_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_THRU_LUT4_0_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__5651),
            .in2(_gnd_net_),
            .in3(N__5622),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_0 ),
            .carryout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_14_14_2 .C_ON=1'b1;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_14_14_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_14_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__5613),
            .in2(_gnd_net_),
            .in3(N__5586),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_1 ),
            .carryout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2 ),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__5749));
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2_THRU_LUT4_0_LC_14_14_3 .C_ON=1'b1;
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2_THRU_LUT4_0_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2_THRU_LUT4_0_LC_14_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2_THRU_LUT4_0_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__5582),
            .in2(_gnd_net_),
            .in3(N__5556),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_2 ),
            .carryout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3_THRU_LUT4_0_LC_14_14_4 .C_ON=1'b1;
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3_THRU_LUT4_0_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3_THRU_LUT4_0_LC_14_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3_THRU_LUT4_0_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__5551),
            .in2(_gnd_net_),
            .in3(N__5523),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_3 ),
            .carryout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4_THRU_LUT4_0_LC_14_14_5 .C_ON=1'b1;
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4_THRU_LUT4_0_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4_THRU_LUT4_0_LC_14_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4_THRU_LUT4_0_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5520),
            .in3(N__5481),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_4 ),
            .carryout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5_THRU_LUT4_0_LC_14_14_6 .C_ON=1'b1;
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5_THRU_LUT4_0_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5_THRU_LUT4_0_LC_14_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5_THRU_LUT4_0_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__6035),
            .in2(_gnd_net_),
            .in3(N__6006),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_5 ),
            .carryout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_14_14_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_14_14_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_14_14_7 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_14_14_7  (
            .in0(N__6002),
            .in1(N__5950),
            .in2(N__5925),
            .in3(N__5928),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__5749));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_14_15_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_14_15_4 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_14_15_4  (
            .in0(N__5895),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5832),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_iobuf_RNO_LC_19_19_5.C_ON=1'b0;
    defparam TACKn_iobuf_RNO_LC_19_19_5.SEQ_MODE=4'b0000;
    defparam TACKn_iobuf_RNO_LC_19_19_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_iobuf_RNO_LC_19_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5718),
            .lcout(N_391_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

module U110_BUFFERS (

    output IDELENn, IDEHRENn, IDEHWENn, IDELATCH

);

//ATA BUFFERS
//DISABLE EVERYTHING FORT NOW

assign IDELENn = 1;
assign IDEHRENn = 1;
assign IDEHWENn = 1;
assign IDELATCH = 1;


endmodule

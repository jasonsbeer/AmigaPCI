// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 25 2024 14:30:47

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    CMA,
    DRA,
    A,
    TSn,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    VBENn,
    CUMBEn,
    CLKRAM,
    C3,
    ASn,
    LDSn,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    DBRn,
    CLK40C,
    CLK40_IN,
    REGSPACEn,
    RAMENn,
    RASn,
    TACKn,
    C1);

    input [1:0] SIZ;
    output [10:0] CMA;
    input [9:0] DRA;
    input [20:0] A;
    input TSn;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    input C3;
    output ASn;
    output LDSn;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    input DBRn;
    output CLK40C;
    input CLK40_IN;
    input REGSPACEn;
    output RAMENn;
    output RASn;
    output TACKn;
    input C1;

    wire N__10026;
    wire N__10025;
    wire N__10024;
    wire N__10017;
    wire N__10016;
    wire N__10015;
    wire N__10008;
    wire N__10007;
    wire N__10006;
    wire N__9999;
    wire N__9998;
    wire N__9997;
    wire N__9990;
    wire N__9989;
    wire N__9988;
    wire N__9981;
    wire N__9980;
    wire N__9979;
    wire N__9972;
    wire N__9971;
    wire N__9970;
    wire N__9963;
    wire N__9962;
    wire N__9961;
    wire N__9954;
    wire N__9953;
    wire N__9952;
    wire N__9945;
    wire N__9944;
    wire N__9943;
    wire N__9936;
    wire N__9935;
    wire N__9934;
    wire N__9927;
    wire N__9926;
    wire N__9925;
    wire N__9918;
    wire N__9917;
    wire N__9916;
    wire N__9909;
    wire N__9908;
    wire N__9907;
    wire N__9900;
    wire N__9899;
    wire N__9898;
    wire N__9891;
    wire N__9890;
    wire N__9889;
    wire N__9882;
    wire N__9881;
    wire N__9880;
    wire N__9873;
    wire N__9872;
    wire N__9871;
    wire N__9864;
    wire N__9863;
    wire N__9862;
    wire N__9855;
    wire N__9854;
    wire N__9853;
    wire N__9846;
    wire N__9845;
    wire N__9844;
    wire N__9837;
    wire N__9836;
    wire N__9835;
    wire N__9828;
    wire N__9827;
    wire N__9826;
    wire N__9819;
    wire N__9818;
    wire N__9817;
    wire N__9810;
    wire N__9809;
    wire N__9808;
    wire N__9801;
    wire N__9800;
    wire N__9799;
    wire N__9792;
    wire N__9791;
    wire N__9790;
    wire N__9783;
    wire N__9782;
    wire N__9781;
    wire N__9774;
    wire N__9773;
    wire N__9772;
    wire N__9765;
    wire N__9764;
    wire N__9763;
    wire N__9756;
    wire N__9755;
    wire N__9754;
    wire N__9747;
    wire N__9746;
    wire N__9745;
    wire N__9738;
    wire N__9737;
    wire N__9736;
    wire N__9729;
    wire N__9728;
    wire N__9727;
    wire N__9720;
    wire N__9719;
    wire N__9718;
    wire N__9711;
    wire N__9710;
    wire N__9709;
    wire N__9702;
    wire N__9701;
    wire N__9700;
    wire N__9693;
    wire N__9692;
    wire N__9691;
    wire N__9684;
    wire N__9683;
    wire N__9682;
    wire N__9675;
    wire N__9674;
    wire N__9673;
    wire N__9666;
    wire N__9665;
    wire N__9664;
    wire N__9657;
    wire N__9656;
    wire N__9655;
    wire N__9648;
    wire N__9647;
    wire N__9646;
    wire N__9639;
    wire N__9638;
    wire N__9637;
    wire N__9630;
    wire N__9629;
    wire N__9628;
    wire N__9621;
    wire N__9620;
    wire N__9619;
    wire N__9612;
    wire N__9611;
    wire N__9610;
    wire N__9603;
    wire N__9602;
    wire N__9601;
    wire N__9594;
    wire N__9593;
    wire N__9592;
    wire N__9585;
    wire N__9584;
    wire N__9583;
    wire N__9576;
    wire N__9575;
    wire N__9574;
    wire N__9567;
    wire N__9566;
    wire N__9565;
    wire N__9558;
    wire N__9557;
    wire N__9556;
    wire N__9549;
    wire N__9548;
    wire N__9547;
    wire N__9540;
    wire N__9539;
    wire N__9538;
    wire N__9531;
    wire N__9530;
    wire N__9529;
    wire N__9522;
    wire N__9521;
    wire N__9520;
    wire N__9513;
    wire N__9512;
    wire N__9511;
    wire N__9504;
    wire N__9503;
    wire N__9502;
    wire N__9495;
    wire N__9494;
    wire N__9493;
    wire N__9486;
    wire N__9485;
    wire N__9484;
    wire N__9477;
    wire N__9476;
    wire N__9475;
    wire N__9468;
    wire N__9467;
    wire N__9466;
    wire N__9459;
    wire N__9458;
    wire N__9457;
    wire N__9450;
    wire N__9449;
    wire N__9448;
    wire N__9441;
    wire N__9440;
    wire N__9439;
    wire N__9432;
    wire N__9431;
    wire N__9430;
    wire N__9423;
    wire N__9422;
    wire N__9421;
    wire N__9414;
    wire N__9413;
    wire N__9412;
    wire N__9405;
    wire N__9404;
    wire N__9403;
    wire N__9396;
    wire N__9395;
    wire N__9394;
    wire N__9387;
    wire N__9386;
    wire N__9385;
    wire N__9378;
    wire N__9377;
    wire N__9376;
    wire N__9369;
    wire N__9368;
    wire N__9367;
    wire N__9360;
    wire N__9359;
    wire N__9358;
    wire N__9351;
    wire N__9350;
    wire N__9349;
    wire N__9342;
    wire N__9341;
    wire N__9340;
    wire N__9333;
    wire N__9332;
    wire N__9331;
    wire N__9324;
    wire N__9323;
    wire N__9322;
    wire N__9315;
    wire N__9314;
    wire N__9313;
    wire N__9296;
    wire N__9295;
    wire N__9292;
    wire N__9289;
    wire N__9286;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9274;
    wire N__9271;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9244;
    wire N__9243;
    wire N__9242;
    wire N__9241;
    wire N__9240;
    wire N__9239;
    wire N__9238;
    wire N__9237;
    wire N__9236;
    wire N__9235;
    wire N__9234;
    wire N__9233;
    wire N__9232;
    wire N__9231;
    wire N__9230;
    wire N__9229;
    wire N__9228;
    wire N__9227;
    wire N__9226;
    wire N__9225;
    wire N__9224;
    wire N__9223;
    wire N__9222;
    wire N__9219;
    wire N__9218;
    wire N__9217;
    wire N__9216;
    wire N__9215;
    wire N__9214;
    wire N__9213;
    wire N__9212;
    wire N__9211;
    wire N__9210;
    wire N__9209;
    wire N__9208;
    wire N__9207;
    wire N__9206;
    wire N__9205;
    wire N__9204;
    wire N__9203;
    wire N__9202;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9112;
    wire N__9109;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9089;
    wire N__9088;
    wire N__9087;
    wire N__9086;
    wire N__9085;
    wire N__9084;
    wire N__9083;
    wire N__9082;
    wire N__9081;
    wire N__9080;
    wire N__9077;
    wire N__9072;
    wire N__9069;
    wire N__9066;
    wire N__9063;
    wire N__9060;
    wire N__9057;
    wire N__9054;
    wire N__9051;
    wire N__9050;
    wire N__9047;
    wire N__9046;
    wire N__9043;
    wire N__9040;
    wire N__9037;
    wire N__9036;
    wire N__9033;
    wire N__9032;
    wire N__9031;
    wire N__9030;
    wire N__9029;
    wire N__9028;
    wire N__9027;
    wire N__9026;
    wire N__9025;
    wire N__9024;
    wire N__9023;
    wire N__9022;
    wire N__9021;
    wire N__9020;
    wire N__9019;
    wire N__9018;
    wire N__9015;
    wire N__9014;
    wire N__9013;
    wire N__9012;
    wire N__9009;
    wire N__9008;
    wire N__9007;
    wire N__9006;
    wire N__9005;
    wire N__9004;
    wire N__9003;
    wire N__9000;
    wire N__8999;
    wire N__8998;
    wire N__8995;
    wire N__8994;
    wire N__8993;
    wire N__8992;
    wire N__8991;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8893;
    wire N__8892;
    wire N__8889;
    wire N__8886;
    wire N__8883;
    wire N__8878;
    wire N__8875;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8858;
    wire N__8857;
    wire N__8854;
    wire N__8853;
    wire N__8850;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8827;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8806;
    wire N__8803;
    wire N__8802;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8779;
    wire N__8776;
    wire N__8773;
    wire N__8768;
    wire N__8767;
    wire N__8764;
    wire N__8761;
    wire N__8760;
    wire N__8759;
    wire N__8758;
    wire N__8757;
    wire N__8756;
    wire N__8755;
    wire N__8754;
    wire N__8753;
    wire N__8750;
    wire N__8749;
    wire N__8744;
    wire N__8741;
    wire N__8736;
    wire N__8731;
    wire N__8728;
    wire N__8725;
    wire N__8722;
    wire N__8719;
    wire N__8718;
    wire N__8717;
    wire N__8714;
    wire N__8709;
    wire N__8706;
    wire N__8697;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8679;
    wire N__8676;
    wire N__8673;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8641;
    wire N__8640;
    wire N__8639;
    wire N__8638;
    wire N__8635;
    wire N__8632;
    wire N__8631;
    wire N__8628;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8620;
    wire N__8619;
    wire N__8616;
    wire N__8615;
    wire N__8614;
    wire N__8609;
    wire N__8604;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8586;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8570;
    wire N__8569;
    wire N__8568;
    wire N__8563;
    wire N__8560;
    wire N__8557;
    wire N__8552;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8521;
    wire N__8520;
    wire N__8519;
    wire N__8518;
    wire N__8515;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8507;
    wire N__8506;
    wire N__8505;
    wire N__8504;
    wire N__8503;
    wire N__8502;
    wire N__8497;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8480;
    wire N__8477;
    wire N__8472;
    wire N__8471;
    wire N__8470;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8446;
    wire N__8443;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8420;
    wire N__8417;
    wire N__8410;
    wire N__8407;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8315;
    wire N__8312;
    wire N__8309;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8219;
    wire N__8216;
    wire N__8213;
    wire N__8210;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8173;
    wire N__8170;
    wire N__8169;
    wire N__8168;
    wire N__8167;
    wire N__8166;
    wire N__8163;
    wire N__8162;
    wire N__8159;
    wire N__8158;
    wire N__8155;
    wire N__8152;
    wire N__8151;
    wire N__8150;
    wire N__8149;
    wire N__8148;
    wire N__8147;
    wire N__8146;
    wire N__8141;
    wire N__8138;
    wire N__8137;
    wire N__8136;
    wire N__8135;
    wire N__8134;
    wire N__8133;
    wire N__8132;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8115;
    wire N__8108;
    wire N__8107;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8099;
    wire N__8094;
    wire N__8093;
    wire N__8092;
    wire N__8089;
    wire N__8086;
    wire N__8081;
    wire N__8080;
    wire N__8077;
    wire N__8076;
    wire N__8073;
    wire N__8064;
    wire N__8063;
    wire N__8062;
    wire N__8061;
    wire N__8056;
    wire N__8051;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8035;
    wire N__8028;
    wire N__8021;
    wire N__8016;
    wire N__8009;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7966;
    wire N__7965;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7951;
    wire N__7948;
    wire N__7945;
    wire N__7942;
    wire N__7939;
    wire N__7936;
    wire N__7931;
    wire N__7928;
    wire N__7923;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7906;
    wire N__7903;
    wire N__7900;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7871;
    wire N__7868;
    wire N__7867;
    wire N__7864;
    wire N__7861;
    wire N__7856;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7844;
    wire N__7841;
    wire N__7838;
    wire N__7837;
    wire N__7834;
    wire N__7833;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7809;
    wire N__7804;
    wire N__7801;
    wire N__7796;
    wire N__7795;
    wire N__7794;
    wire N__7791;
    wire N__7786;
    wire N__7781;
    wire N__7778;
    wire N__7777;
    wire N__7774;
    wire N__7771;
    wire N__7766;
    wire N__7763;
    wire N__7762;
    wire N__7759;
    wire N__7756;
    wire N__7751;
    wire N__7748;
    wire N__7745;
    wire N__7744;
    wire N__7743;
    wire N__7740;
    wire N__7735;
    wire N__7730;
    wire N__7727;
    wire N__7724;
    wire N__7721;
    wire N__7718;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7708;
    wire N__7703;
    wire N__7702;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7691;
    wire N__7686;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7650;
    wire N__7647;
    wire N__7644;
    wire N__7641;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7618;
    wire N__7615;
    wire N__7612;
    wire N__7609;
    wire N__7606;
    wire N__7601;
    wire N__7598;
    wire N__7595;
    wire N__7592;
    wire N__7589;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7564;
    wire N__7561;
    wire N__7558;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7526;
    wire N__7525;
    wire N__7522;
    wire N__7519;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7505;
    wire N__7502;
    wire N__7499;
    wire N__7496;
    wire N__7493;
    wire N__7490;
    wire N__7489;
    wire N__7486;
    wire N__7483;
    wire N__7480;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7453;
    wire N__7450;
    wire N__7447;
    wire N__7444;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7421;
    wire N__7418;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7382;
    wire N__7379;
    wire N__7376;
    wire N__7373;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7363;
    wire N__7362;
    wire N__7359;
    wire N__7354;
    wire N__7349;
    wire N__7346;
    wire N__7345;
    wire N__7342;
    wire N__7341;
    wire N__7338;
    wire N__7333;
    wire N__7328;
    wire N__7325;
    wire N__7322;
    wire N__7319;
    wire N__7316;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7244;
    wire N__7241;
    wire N__7238;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7216;
    wire N__7213;
    wire N__7210;
    wire N__7205;
    wire N__7204;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7194;
    wire N__7193;
    wire N__7190;
    wire N__7189;
    wire N__7188;
    wire N__7185;
    wire N__7182;
    wire N__7181;
    wire N__7180;
    wire N__7179;
    wire N__7178;
    wire N__7177;
    wire N__7174;
    wire N__7171;
    wire N__7168;
    wire N__7165;
    wire N__7160;
    wire N__7155;
    wire N__7150;
    wire N__7147;
    wire N__7130;
    wire N__7129;
    wire N__7128;
    wire N__7127;
    wire N__7126;
    wire N__7125;
    wire N__7118;
    wire N__7115;
    wire N__7114;
    wire N__7113;
    wire N__7112;
    wire N__7109;
    wire N__7108;
    wire N__7105;
    wire N__7102;
    wire N__7099;
    wire N__7098;
    wire N__7097;
    wire N__7092;
    wire N__7085;
    wire N__7078;
    wire N__7073;
    wire N__7070;
    wire N__7061;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7044;
    wire N__7043;
    wire N__7038;
    wire N__7035;
    wire N__7032;
    wire N__7025;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6989;
    wire N__6986;
    wire N__6983;
    wire N__6980;
    wire N__6977;
    wire N__6976;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6965;
    wire N__6964;
    wire N__6963;
    wire N__6962;
    wire N__6959;
    wire N__6956;
    wire N__6955;
    wire N__6954;
    wire N__6951;
    wire N__6946;
    wire N__6943;
    wire N__6940;
    wire N__6935;
    wire N__6930;
    wire N__6925;
    wire N__6914;
    wire N__6913;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6898;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6865;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6800;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6755;
    wire N__6752;
    wire N__6749;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6710;
    wire N__6707;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6646;
    wire N__6645;
    wire N__6644;
    wire N__6641;
    wire N__6640;
    wire N__6639;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6626;
    wire N__6619;
    wire N__6608;
    wire N__6607;
    wire N__6606;
    wire N__6605;
    wire N__6604;
    wire N__6603;
    wire N__6600;
    wire N__6597;
    wire N__6590;
    wire N__6587;
    wire N__6578;
    wire N__6577;
    wire N__6576;
    wire N__6575;
    wire N__6574;
    wire N__6571;
    wire N__6568;
    wire N__6561;
    wire N__6554;
    wire N__6553;
    wire N__6552;
    wire N__6551;
    wire N__6548;
    wire N__6543;
    wire N__6540;
    wire N__6533;
    wire N__6532;
    wire N__6531;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6523;
    wire N__6520;
    wire N__6519;
    wire N__6516;
    wire N__6511;
    wire N__6504;
    wire N__6497;
    wire N__6494;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6467;
    wire N__6464;
    wire N__6461;
    wire N__6458;
    wire N__6455;
    wire N__6452;
    wire N__6449;
    wire N__6446;
    wire N__6443;
    wire N__6440;
    wire N__6437;
    wire N__6434;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6419;
    wire N__6416;
    wire N__6413;
    wire N__6410;
    wire N__6407;
    wire N__6406;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6389;
    wire N__6388;
    wire N__6387;
    wire N__6384;
    wire N__6379;
    wire N__6374;
    wire N__6373;
    wire N__6372;
    wire N__6371;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6357;
    wire N__6350;
    wire N__6349;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6326;
    wire N__6323;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6305;
    wire N__6304;
    wire N__6301;
    wire N__6300;
    wire N__6295;
    wire N__6292;
    wire N__6287;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6265;
    wire N__6264;
    wire N__6263;
    wire N__6258;
    wire N__6253;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6236;
    wire N__6233;
    wire N__6232;
    wire N__6231;
    wire N__6230;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6205;
    wire N__6204;
    wire N__6203;
    wire N__6198;
    wire N__6193;
    wire N__6190;
    wire N__6187;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6173;
    wire N__6170;
    wire N__6169;
    wire N__6166;
    wire N__6163;
    wire N__6160;
    wire N__6157;
    wire N__6154;
    wire N__6151;
    wire N__6146;
    wire N__6143;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6124;
    wire N__6121;
    wire N__6118;
    wire N__6113;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6080;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6065;
    wire N__6062;
    wire N__6059;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6047;
    wire N__6044;
    wire N__6041;
    wire N__6038;
    wire N__6035;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6025;
    wire N__6024;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6014;
    wire N__6011;
    wire N__6006;
    wire N__6003;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5984;
    wire N__5983;
    wire N__5982;
    wire N__5979;
    wire N__5974;
    wire N__5973;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5959;
    wire N__5958;
    wire N__5957;
    wire N__5948;
    wire N__5941;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5915;
    wire N__5914;
    wire N__5913;
    wire N__5912;
    wire N__5907;
    wire N__5902;
    wire N__5897;
    wire N__5894;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5851;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5838;
    wire N__5835;
    wire N__5828;
    wire N__5825;
    wire N__5822;
    wire N__5819;
    wire N__5818;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5801;
    wire N__5800;
    wire N__5799;
    wire N__5798;
    wire N__5795;
    wire N__5794;
    wire N__5793;
    wire N__5792;
    wire N__5791;
    wire N__5790;
    wire N__5789;
    wire N__5788;
    wire N__5787;
    wire N__5784;
    wire N__5783;
    wire N__5782;
    wire N__5781;
    wire N__5778;
    wire N__5775;
    wire N__5772;
    wire N__5765;
    wire N__5758;
    wire N__5753;
    wire N__5750;
    wire N__5747;
    wire N__5746;
    wire N__5743;
    wire N__5742;
    wire N__5741;
    wire N__5738;
    wire N__5737;
    wire N__5736;
    wire N__5735;
    wire N__5734;
    wire N__5733;
    wire N__5732;
    wire N__5731;
    wire N__5728;
    wire N__5723;
    wire N__5720;
    wire N__5713;
    wire N__5706;
    wire N__5701;
    wire N__5696;
    wire N__5693;
    wire N__5686;
    wire N__5681;
    wire N__5660;
    wire N__5659;
    wire N__5658;
    wire N__5657;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5646;
    wire N__5643;
    wire N__5642;
    wire N__5639;
    wire N__5638;
    wire N__5637;
    wire N__5634;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5616;
    wire N__5615;
    wire N__5614;
    wire N__5613;
    wire N__5612;
    wire N__5611;
    wire N__5608;
    wire N__5607;
    wire N__5606;
    wire N__5605;
    wire N__5602;
    wire N__5597;
    wire N__5592;
    wire N__5587;
    wire N__5582;
    wire N__5579;
    wire N__5572;
    wire N__5567;
    wire N__5562;
    wire N__5543;
    wire N__5542;
    wire N__5541;
    wire N__5536;
    wire N__5535;
    wire N__5532;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5520;
    wire N__5513;
    wire N__5510;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5498;
    wire N__5495;
    wire N__5494;
    wire N__5493;
    wire N__5492;
    wire N__5487;
    wire N__5482;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5446;
    wire N__5443;
    wire N__5442;
    wire N__5439;
    wire N__5438;
    wire N__5435;
    wire N__5428;
    wire N__5423;
    wire N__5420;
    wire N__5419;
    wire N__5416;
    wire N__5413;
    wire N__5408;
    wire N__5407;
    wire N__5406;
    wire N__5403;
    wire N__5402;
    wire N__5401;
    wire N__5398;
    wire N__5397;
    wire N__5396;
    wire N__5395;
    wire N__5392;
    wire N__5391;
    wire N__5388;
    wire N__5385;
    wire N__5376;
    wire N__5373;
    wire N__5370;
    wire N__5367;
    wire N__5354;
    wire N__5353;
    wire N__5350;
    wire N__5349;
    wire N__5346;
    wire N__5343;
    wire N__5340;
    wire N__5339;
    wire N__5338;
    wire N__5335;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5327;
    wire N__5326;
    wire N__5325;
    wire N__5324;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5314;
    wire N__5311;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5292;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5263;
    wire N__5262;
    wire N__5261;
    wire N__5260;
    wire N__5259;
    wire N__5258;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5247;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5233;
    wire N__5228;
    wire N__5225;
    wire N__5220;
    wire N__5207;
    wire N__5204;
    wire N__5203;
    wire N__5202;
    wire N__5197;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5187;
    wire N__5182;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5162;
    wire N__5161;
    wire N__5160;
    wire N__5155;
    wire N__5152;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5111;
    wire N__5110;
    wire N__5109;
    wire N__5106;
    wire N__5101;
    wire N__5096;
    wire N__5095;
    wire N__5092;
    wire N__5091;
    wire N__5090;
    wire N__5089;
    wire N__5086;
    wire N__5085;
    wire N__5082;
    wire N__5081;
    wire N__5078;
    wire N__5077;
    wire N__5076;
    wire N__5075;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5053;
    wire N__5048;
    wire N__5043;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5014;
    wire N__5011;
    wire N__5008;
    wire N__5003;
    wire N__5000;
    wire N__4999;
    wire N__4998;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4978;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4945;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4921;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4903;
    wire N__4898;
    wire N__4895;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4882;
    wire N__4879;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4864;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4834;
    wire N__4833;
    wire N__4832;
    wire N__4829;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4811;
    wire N__4808;
    wire N__4807;
    wire N__4804;
    wire N__4801;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4784;
    wire N__4783;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4766;
    wire N__4765;
    wire N__4760;
    wire N__4757;
    wire N__4756;
    wire N__4755;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4738;
    wire N__4737;
    wire N__4736;
    wire N__4733;
    wire N__4726;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4691;
    wire N__4690;
    wire N__4687;
    wire N__4684;
    wire N__4679;
    wire N__4678;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4657;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4621;
    wire N__4618;
    wire N__4615;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4558;
    wire N__4557;
    wire N__4554;
    wire N__4549;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4537;
    wire N__4534;
    wire N__4533;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4521;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4489;
    wire N__4486;
    wire N__4483;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4456;
    wire N__4455;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4439;
    wire N__4436;
    wire N__4433;
    wire N__4432;
    wire N__4429;
    wire N__4428;
    wire N__4425;
    wire N__4424;
    wire N__4421;
    wire N__4414;
    wire N__4411;
    wire N__4406;
    wire N__4403;
    wire N__4402;
    wire N__4401;
    wire N__4398;
    wire N__4393;
    wire N__4388;
    wire N__4387;
    wire N__4384;
    wire N__4381;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4366;
    wire N__4365;
    wire N__4364;
    wire N__4363;
    wire N__4360;
    wire N__4357;
    wire N__4350;
    wire N__4343;
    wire N__4342;
    wire N__4339;
    wire N__4336;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4303;
    wire N__4300;
    wire N__4297;
    wire N__4292;
    wire N__4291;
    wire N__4288;
    wire N__4285;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4223;
    wire N__4222;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4212;
    wire N__4209;
    wire N__4202;
    wire N__4201;
    wire N__4200;
    wire N__4197;
    wire N__4192;
    wire N__4189;
    wire N__4184;
    wire N__4181;
    wire N__4180;
    wire N__4179;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4157;
    wire N__4154;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4142;
    wire N__4139;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4090;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4037;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4025;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4012;
    wire N__4011;
    wire N__4006;
    wire N__4003;
    wire N__3998;
    wire N__3997;
    wire N__3994;
    wire N__3991;
    wire N__3986;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3976;
    wire N__3975;
    wire N__3972;
    wire N__3967;
    wire N__3962;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3938;
    wire N__3935;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3914;
    wire N__3911;
    wire N__3908;
    wire N__3905;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3892;
    wire N__3891;
    wire N__3890;
    wire N__3883;
    wire N__3880;
    wire N__3877;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3850;
    wire N__3847;
    wire N__3844;
    wire N__3839;
    wire N__3838;
    wire N__3837;
    wire N__3836;
    wire N__3827;
    wire N__3824;
    wire N__3823;
    wire N__3820;
    wire N__3817;
    wire N__3812;
    wire N__3809;
    wire N__3808;
    wire N__3805;
    wire N__3802;
    wire N__3797;
    wire N__3794;
    wire N__3791;
    wire N__3788;
    wire N__3785;
    wire N__3782;
    wire N__3779;
    wire N__3776;
    wire N__3773;
    wire N__3770;
    wire N__3767;
    wire N__3764;
    wire N__3761;
    wire N__3758;
    wire N__3755;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3680;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3668;
    wire N__3665;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3629;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3617;
    wire N__3614;
    wire N__3611;
    wire N__3608;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_OUT_i_i;
    wire N_839_i;
    wire A_c_13;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4_cascade_ ;
    wire A_c_6;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.N_319 ;
    wire CMA_c_4;
    wire A_c_12;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_ ;
    wire A_c_5;
    wire \U712_CHIP_RAM.N_318 ;
    wire CLK40_OUT_i_i;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_0_a2_i_0_cascade_ ;
    wire \U712_CHIP_RAM.N_181 ;
    wire CLK40_OUT_i;
    wire TACK_OUTn;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire CPU_TACKm;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0_cascade_ ;
    wire \U712_CYCLE_TERM.N_307_i_0_en_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire TACK_EN_i_ess;
    wire \U712_CYCLE_TERM.N_307_i_0_en_0 ;
    wire VBENn_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_ ;
    wire RAMSPACEn_c;
    wire DBRn_c;
    wire \U712_CHIP_RAM.N_287_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_1_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ;
    wire REG_TACK;
    wire TSn_c;
    wire REGSPACEn_c;
    wire \U712_REG_SM.REG_CYCLE_GOZ0 ;
    wire \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1 ;
    wire \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_ ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire \U712_REG_SM.LDS_OUT_2_0_a2Z0Z_0 ;
    wire \U712_REG_SM.N_342 ;
    wire \U712_REG_SM.LDS_OUTZ0 ;
    wire U712_REG_SM_un1_LDSn_i;
    wire \U712_REG_SM.UDS_OUTZ0 ;
    wire \U712_REG_SM.DS_ENZ0 ;
    wire U712_REG_SM_un1_UDSn_i;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.N_287 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_1_0_cascade_ ;
    wire \U712_CHIP_RAM.N_273_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_0 ;
    wire \U712_CHIP_RAM.N_347_cascade_ ;
    wire \U712_CHIP_RAM.N_378_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_tz ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_0_a2_0_a2_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER50_cascade_ ;
    wire AWEn_c;
    wire \U712_CHIP_RAM.N_296_i ;
    wire \U712_CHIP_RAM.SDRAM_CMD_e_1_2_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_0_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0 ;
    wire DBDIR_c;
    wire N_188;
    wire U712_REG_SM_DBR_SYNC_1;
    wire \U712_REG_SM.N_288_cascade_ ;
    wire U712_REG_SM_DBR_SYNC_0;
    wire \U712_REG_SM.STATE_COUNTZ0Z_5 ;
    wire \U712_REG_SM.N_301_cascade_ ;
    wire \U712_REG_SM.N_288 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.N_301 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire REG_CYCLEm;
    wire DRDENn_c;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.N_341 ;
    wire \U712_REG_SM.N_294_cascade_ ;
    wire \U712_REG_SM.N_373 ;
    wire \U712_REG_SM.N_292_cascade_ ;
    wire \U712_REG_SM.N_507 ;
    wire RnW_c;
    wire \U712_REG_SM.N_104 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_REG_SM.N_372 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_6 ;
    wire ASn_c;
    wire \U712_REG_SM.N_186_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_0_a2_2_cascade_ ;
    wire \U712_CHIP_RAM.N_393 ;
    wire \U712_CHIP_RAM.N_310 ;
    wire \U712_CHIP_RAM.N_310_cascade_ ;
    wire \U712_CHIP_RAM.N_46 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_3_0_a2_i_0_cascade_ ;
    wire \U712_CHIP_RAM.N_179_cascade_ ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.REFRESH_CYCLEZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.N_438_cascade_ ;
    wire \U712_CHIP_RAM.N_289 ;
    wire \U712_CHIP_RAM.N_425_cascade_ ;
    wire \U712_CHIP_RAM.N_424 ;
    wire \U712_CHIP_RAM.N_302 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.REFRESH_CYCLE_START_2_0_a2_1_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_438 ;
    wire \U712_CHIP_RAM.N_284 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_1_cascade_ ;
    wire \U712_CHIP_RAM.N_272 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_cascade_ ;
    wire \U712_CHIP_RAM.DBENn_7_0_a2_0 ;
    wire \U712_CHIP_RAM.N_347 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_3_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_2_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER50 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_273 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_1_0_cascade_ ;
    wire \U712_CHIP_RAM.N_305 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ;
    wire \U712_CHIP_RAM.REFRESH_RST_cascade_ ;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0_cascade_ ;
    wire N_192_i;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0 ;
    wire N_194_i;
    wire SIZ_c_0;
    wire DBENn_c;
    wire RAMENn_c;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_cascade_ ;
    wire N_196_i;
    wire \U712_BYTE_ENABLE.N_404 ;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0 ;
    wire \U712_BYTE_ENABLE.N_411_cascade_ ;
    wire N_198_i;
    wire \U712_BYTE_ENABLE.N_405 ;
    wire \U712_REG_SM.N_292 ;
    wire \U712_REG_SM.N_298 ;
    wire \U712_REG_SM.N_294 ;
    wire \U712_REG_SM.N_309 ;
    wire \U712_REG_SM.N_282 ;
    wire \U712_REG_SM.N_282_cascade_ ;
    wire \U712_REG_SM.N_306 ;
    wire SIZ_c_1;
    wire \U712_BYTE_ENABLE.N_407 ;
    wire A_c_1;
    wire A_c_0;
    wire \U712_BYTE_ENABLE.N_409 ;
    wire C1_c;
    wire C3_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_2 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_2 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire CMA_c_2;
    wire CMA_c_1;
    wire CMA_c_10;
    wire A_c_11;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_ ;
    wire A_c_4;
    wire \U712_CHIP_RAM.N_317 ;
    wire A_c_14;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5_cascade_ ;
    wire A_c_7;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire A_c_15;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6_cascade_ ;
    wire A_c_8;
    wire A_c_9;
    wire A_c_2;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0_cascade_ ;
    wire \U712_CHIP_RAM.N_315_cascade_ ;
    wire CMA_c_0;
    wire A_c_3;
    wire A_c_10;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_ ;
    wire \U712_CHIP_RAM.N_316 ;
    wire \U712_CHIP_RAM.N_425 ;
    wire \U712_CHIP_RAM.N_276 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_a2_0 ;
    wire \U712_CHIP_RAM.N_314 ;
    wire \U712_CHIP_RAM.N_293 ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.un1_CMA31_0_i ;
    wire \U712_CHIP_RAM.REFRESH_RNO_0Z0Z_0_cascade_ ;
    wire \U712_CHIP_RAM.REFRESHZ0Z_0 ;
    wire \U712_CHIP_RAM.REFRESH9lt7_cascade_ ;
    wire \U712_CHIP_RAM.REFRESHZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH9lto7_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.N_321 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.N_320 ;
    wire CMA_c_5;
    wire A_c_17;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire CONSTANT_ONE_NET;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ;
    wire bfn_12_8_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH9lto2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire RESETn_c;
    wire RESETn_c_i;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire A_c_18;
    wire \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_ ;
    wire A_c_16;
    wire \U712_CHIP_RAM.N_322_cascade_ ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.CMA_5_i_0_8 ;
    wire A_c_19;
    wire \U712_CHIP_RAM.CMA_5_i_0_8_cascade_ ;
    wire CPU_CYCLEm;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.un1_CMA31_0_i_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ;
    wire CASLn_c;
    wire CASUn_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire WEn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CASn_c;
    wire RAS0n_c;
    wire RAS1n_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire _gnd_net_;
    wire CLK80_OUT;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ;
    wire RESETn_c_i_g;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_OUT_i),
            .REFERENCECLK(N__3617),
            .RESETB(N__7409),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_OUT),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__10026),
            .DIN(N__10025),
            .DOUT(N__10024),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__10026),
            .PADOUT(N__10025),
            .PADIN(N__10024),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6038),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__10017),
            .DIN(N__10016),
            .DOUT(N__10015),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__10017),
            .PADOUT(N__10016),
            .PADIN(N__10015),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__10008),
            .DIN(N__10007),
            .DOUT(N__10006),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__10008),
            .PADOUT(N__10007),
            .PADIN(N__10006),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8396),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__9999),
            .DIN(N__9998),
            .DOUT(N__9997),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__9999),
            .PADOUT(N__9998),
            .PADIN(N__9997),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4589),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__9990),
            .DIN(N__9989),
            .DOUT(N__9988),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__9990),
            .PADOUT(N__9989),
            .PADIN(N__9988),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__9981),
            .DIN(N__9980),
            .DOUT(N__9979),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__9981),
            .PADOUT(N__9980),
            .PADIN(N__9979),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__9972),
            .DIN(N__9971),
            .DOUT(N__9970),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__9972),
            .PADOUT(N__9971),
            .PADIN(N__9970),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__9963),
            .DIN(N__9962),
            .DOUT(N__9961),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__9963),
            .PADOUT(N__9962),
            .PADIN(N__9961),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__9954),
            .DIN(N__9953),
            .DOUT(N__9952),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__9954),
            .PADOUT(N__9953),
            .PADIN(N__9952),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__9945),
            .DIN(N__9944),
            .DOUT(N__9943),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__9945),
            .PADOUT(N__9944),
            .PADIN(N__9943),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__9936),
            .DIN(N__9935),
            .DOUT(N__9934),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__9936),
            .PADOUT(N__9935),
            .PADIN(N__9934),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8225),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__9927),
            .DIN(N__9926),
            .DOUT(N__9925),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__9927),
            .PADOUT(N__9926),
            .PADIN(N__9925),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5996),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__9918),
            .DIN(N__9917),
            .DOUT(N__9916),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__9918),
            .PADOUT(N__9917),
            .PADIN(N__9916),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__9909),
            .DIN(N__9908),
            .DOUT(N__9907),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__9909),
            .PADOUT(N__9908),
            .PADIN(N__9907),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__9900),
            .DIN(N__9899),
            .DOUT(N__9898),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__9900),
            .PADOUT(N__9899),
            .PADIN(N__9898),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3917),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__9891),
            .DIN(N__9890),
            .DOUT(N__9889),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__9891),
            .PADOUT(N__9890),
            .PADIN(N__9889),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__9882),
            .DIN(N__9881),
            .DOUT(N__9880),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__9882),
            .PADOUT(N__9881),
            .PADIN(N__9880),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__9873),
            .DIN(N__9872),
            .DOUT(N__9871),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__9873),
            .PADOUT(N__9872),
            .PADIN(N__9871),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6719),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__9864),
            .DIN(N__9863),
            .DOUT(N__9862),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__9864),
            .PADOUT(N__9863),
            .PADIN(N__9862),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__9855),
            .DIN(N__9854),
            .DOUT(N__9853),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__9855),
            .PADOUT(N__9854),
            .PADIN(N__9853),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7025),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__9846),
            .DIN(N__9845),
            .DOUT(N__9844),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__9846),
            .PADOUT(N__9845),
            .PADIN(N__9844),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__9837),
            .DIN(N__9836),
            .DOUT(N__9835),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__9837),
            .PADOUT(N__9836),
            .PADIN(N__9835),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__9828),
            .DIN(N__9827),
            .DOUT(N__9826),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__9828),
            .PADOUT(N__9827),
            .PADIN(N__9826),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__9819),
            .DIN(N__9818),
            .DOUT(N__9817),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__9819),
            .PADOUT(N__9818),
            .PADIN(N__9817),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__9810),
            .DIN(N__9809),
            .DOUT(N__9808),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__9810),
            .PADOUT(N__9809),
            .PADIN(N__9808),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__9801),
            .DIN(N__9800),
            .DOUT(N__9799),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__9801),
            .PADOUT(N__9800),
            .PADIN(N__9799),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5141),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__9792),
            .DIN(N__9791),
            .DOUT(N__9790),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__9792),
            .PADOUT(N__9791),
            .PADIN(N__9790),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__9783),
            .DIN(N__9782),
            .DOUT(N__9781),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__9783),
            .PADOUT(N__9782),
            .PADIN(N__9781),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__9774),
            .DIN(N__9773),
            .DOUT(N__9772),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__9774),
            .PADOUT(N__9773),
            .PADIN(N__9772),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__9765),
            .DIN(N__9764),
            .DOUT(N__9763),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__9765),
            .PADOUT(N__9764),
            .PADIN(N__9763),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__9756),
            .DIN(N__9755),
            .DOUT(N__9754),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__9756),
            .PADOUT(N__9755),
            .PADIN(N__9754),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__9747),
            .DIN(N__9746),
            .DOUT(N__9745),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__9747),
            .PADOUT(N__9746),
            .PADIN(N__9745),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7313),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__9738),
            .DIN(N__9737),
            .DOUT(N__9736),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__9738),
            .PADOUT(N__9737),
            .PADIN(N__9736),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__9729),
            .DIN(N__9728),
            .DOUT(N__9727),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__9729),
            .PADOUT(N__9728),
            .PADIN(N__9727),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__9720),
            .DIN(N__9719),
            .DOUT(N__9718),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__9720),
            .PADOUT(N__9719),
            .PADIN(N__9718),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__9711),
            .DIN(N__9710),
            .DOUT(N__9709),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__9711),
            .PADOUT(N__9710),
            .PADIN(N__9709),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__9702),
            .DIN(N__9701),
            .DOUT(N__9700),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__9702),
            .PADOUT(N__9701),
            .PADIN(N__9700),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3674),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__9693),
            .DIN(N__9692),
            .DOUT(N__9691),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__9693),
            .PADOUT(N__9692),
            .PADIN(N__9691),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4331),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__9684),
            .DIN(N__9683),
            .DOUT(N__9682),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__9684),
            .PADOUT(N__9683),
            .PADIN(N__9682),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__9675),
            .DIN(N__9674),
            .DOUT(N__9673),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__9675),
            .PADOUT(N__9674),
            .PADIN(N__9673),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8660),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__9666),
            .DIN(N__9665),
            .DOUT(N__9664),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__9666),
            .PADOUT(N__9665),
            .PADIN(N__9664),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__9657),
            .DIN(N__9656),
            .DOUT(N__9655),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__9657),
            .PADOUT(N__9656),
            .PADIN(N__9655),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__9648),
            .DIN(N__9647),
            .DOUT(N__9646),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__9648),
            .PADOUT(N__9647),
            .PADIN(N__9646),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3653),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__9639),
            .DIN(N__9638),
            .DOUT(N__9637),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__9639),
            .PADOUT(N__9638),
            .PADIN(N__9637),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__9630),
            .DIN(N__9629),
            .DOUT(N__9628),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__9630),
            .PADOUT(N__9629),
            .PADIN(N__9628),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4898),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__9621),
            .DIN(N__9620),
            .DOUT(N__9619),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__9621),
            .PADOUT(N__9620),
            .PADIN(N__9619),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3758),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__9612),
            .DIN(N__9611),
            .DOUT(N__9610),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__9612),
            .PADOUT(N__9611),
            .PADIN(N__9610),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__9603),
            .DIN(N__9602),
            .DOUT(N__9601),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__9603),
            .PADOUT(N__9602),
            .PADIN(N__9601),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_0_iopad (
            .OE(N__9594),
            .DIN(N__9593),
            .DOUT(N__9592),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__9594),
            .PADOUT(N__9593),
            .PADIN(N__9592),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__9585),
            .DIN(N__9584),
            .DOUT(N__9583),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__9585),
            .PADOUT(N__9584),
            .PADIN(N__9583),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6476),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__9576),
            .DIN(N__9575),
            .DOUT(N__9574),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__9576),
            .PADOUT(N__9575),
            .PADIN(N__9574),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__9567),
            .DIN(N__9566),
            .DOUT(N__9565),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__9567),
            .PADOUT(N__9566),
            .PADIN(N__9565),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3737),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__9558),
            .DIN(N__9557),
            .DOUT(N__9556),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__9558),
            .PADOUT(N__9557),
            .PADIN(N__9556),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4721),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__9549),
            .DIN(N__9548),
            .DOUT(N__9547),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__9549),
            .PADOUT(N__9548),
            .PADIN(N__9547),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5888),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__9540),
            .DIN(N__9539),
            .DOUT(N__9538),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__9540),
            .PADOUT(N__9539),
            .PADIN(N__9538),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7988),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__9531),
            .DIN(N__9530),
            .DOUT(N__9529),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__9531),
            .PADOUT(N__9530),
            .PADIN(N__9529),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4894),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__9522),
            .DIN(N__9521),
            .DOUT(N__9520),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__9522),
            .PADOUT(N__9521),
            .PADIN(N__9520),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__9513),
            .DIN(N__9512),
            .DOUT(N__9511),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__9513),
            .PADOUT(N__9512),
            .PADIN(N__9511),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__9504),
            .DIN(N__9503),
            .DOUT(N__9502),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__9504),
            .PADOUT(N__9503),
            .PADIN(N__9502),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5933),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__9495),
            .DIN(N__9494),
            .DOUT(N__9493),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__9495),
            .PADOUT(N__9494),
            .PADIN(N__9493),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8543),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__9486),
            .DIN(N__9485),
            .DOUT(N__9484),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__9486),
            .PADOUT(N__9485),
            .PADIN(N__9484),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4628),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__9477),
            .DIN(N__9476),
            .DOUT(N__9475),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__9477),
            .PADOUT(N__9476),
            .PADIN(N__9475),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6083),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__9468),
            .DIN(N__9467),
            .DOUT(N__9466),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__9468),
            .PADOUT(N__9467),
            .PADIN(N__9466),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__9459),
            .DIN(N__9458),
            .DOUT(N__9457),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__9459),
            .PADOUT(N__9458),
            .PADIN(N__9457),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__9450),
            .DIN(N__9449),
            .DOUT(N__9448),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__9450),
            .PADOUT(N__9449),
            .PADIN(N__9448),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__9441),
            .DIN(N__9440),
            .DOUT(N__9439),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__9441),
            .PADOUT(N__9440),
            .PADIN(N__9439),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__9432),
            .DIN(N__9431),
            .DOUT(N__9430),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__9432),
            .PADOUT(N__9431),
            .PADIN(N__9430),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6488),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__9423),
            .DIN(N__9422),
            .DOUT(N__9421),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__9423),
            .PADOUT(N__9422),
            .PADIN(N__9421),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__9414),
            .DIN(N__9413),
            .DOUT(N__9412),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__9414),
            .PADOUT(N__9413),
            .PADIN(N__9412),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6110),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__9405),
            .DIN(N__9404),
            .DOUT(N__9403),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__9405),
            .PADOUT(N__9404),
            .PADIN(N__9403),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3635),
            .DIN0(),
            .DOUT0(N__3860),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__9396),
            .DIN(N__9395),
            .DOUT(N__9394),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__9396),
            .PADOUT(N__9395),
            .PADIN(N__9394),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6497),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__9387),
            .DIN(N__9386),
            .DOUT(N__9385),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__9387),
            .PADOUT(N__9386),
            .PADIN(N__9385),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__9378),
            .DIN(N__9377),
            .DOUT(N__9376),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__9378),
            .PADOUT(N__9377),
            .PADIN(N__9376),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__9369),
            .DIN(N__9368),
            .DOUT(N__9367),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__9369),
            .PADOUT(N__9368),
            .PADIN(N__9367),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7256),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__9360),
            .DIN(N__9359),
            .DOUT(N__9358),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__9360),
            .PADOUT(N__9359),
            .PADIN(N__9358),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__9351),
            .DIN(N__9350),
            .DOUT(N__9349),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__9351),
            .PADOUT(N__9350),
            .PADIN(N__9349),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__9342),
            .DIN(N__9341),
            .DOUT(N__9340),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__9342),
            .PADOUT(N__9341),
            .PADIN(N__9340),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__9333),
            .DIN(N__9332),
            .DOUT(N__9331),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__9333),
            .PADOUT(N__9332),
            .PADIN(N__9331),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__9324),
            .DIN(N__9323),
            .DOUT(N__9322),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__9324),
            .PADOUT(N__9323),
            .PADIN(N__9322),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7286),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__9315),
            .DIN(N__9314),
            .DOUT(N__9313),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__9315),
            .PADOUT(N__9314),
            .PADIN(N__9313),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4268),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2203 (
            .O(N__9296),
            .I(N__9292));
    InMux I__2202 (
            .O(N__9295),
            .I(N__9289));
    LocalMux I__2201 (
            .O(N__9292),
            .I(N__9286));
    LocalMux I__2200 (
            .O(N__9289),
            .I(N__9283));
    Span4Mux_v I__2199 (
            .O(N__9286),
            .I(N__9280));
    Span4Mux_h I__2198 (
            .O(N__9283),
            .I(N__9277));
    Span4Mux_v I__2197 (
            .O(N__9280),
            .I(N__9274));
    Span4Mux_v I__2196 (
            .O(N__9277),
            .I(N__9271));
    Sp12to4 I__2195 (
            .O(N__9274),
            .I(N__9266));
    Sp12to4 I__2194 (
            .O(N__9271),
            .I(N__9266));
    Span12Mux_h I__2193 (
            .O(N__9266),
            .I(N__9263));
    Span12Mux_v I__2192 (
            .O(N__9263),
            .I(N__9260));
    Odrv12 I__2191 (
            .O(N__9260),
            .I(DRA_c_0));
    InMux I__2190 (
            .O(N__9257),
            .I(N__9254));
    LocalMux I__2189 (
            .O(N__9254),
            .I(N__9251));
    Odrv4 I__2188 (
            .O(N__9251),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__2187 (
            .O(N__9248),
            .I(N__9245));
    LocalMux I__2186 (
            .O(N__9245),
            .I(N__9219));
    ClkMux I__2185 (
            .O(N__9244),
            .I(N__9119));
    ClkMux I__2184 (
            .O(N__9243),
            .I(N__9119));
    ClkMux I__2183 (
            .O(N__9242),
            .I(N__9119));
    ClkMux I__2182 (
            .O(N__9241),
            .I(N__9119));
    ClkMux I__2181 (
            .O(N__9240),
            .I(N__9119));
    ClkMux I__2180 (
            .O(N__9239),
            .I(N__9119));
    ClkMux I__2179 (
            .O(N__9238),
            .I(N__9119));
    ClkMux I__2178 (
            .O(N__9237),
            .I(N__9119));
    ClkMux I__2177 (
            .O(N__9236),
            .I(N__9119));
    ClkMux I__2176 (
            .O(N__9235),
            .I(N__9119));
    ClkMux I__2175 (
            .O(N__9234),
            .I(N__9119));
    ClkMux I__2174 (
            .O(N__9233),
            .I(N__9119));
    ClkMux I__2173 (
            .O(N__9232),
            .I(N__9119));
    ClkMux I__2172 (
            .O(N__9231),
            .I(N__9119));
    ClkMux I__2171 (
            .O(N__9230),
            .I(N__9119));
    ClkMux I__2170 (
            .O(N__9229),
            .I(N__9119));
    ClkMux I__2169 (
            .O(N__9228),
            .I(N__9119));
    ClkMux I__2168 (
            .O(N__9227),
            .I(N__9119));
    ClkMux I__2167 (
            .O(N__9226),
            .I(N__9119));
    ClkMux I__2166 (
            .O(N__9225),
            .I(N__9119));
    ClkMux I__2165 (
            .O(N__9224),
            .I(N__9119));
    ClkMux I__2164 (
            .O(N__9223),
            .I(N__9119));
    ClkMux I__2163 (
            .O(N__9222),
            .I(N__9119));
    Glb2LocalMux I__2162 (
            .O(N__9219),
            .I(N__9119));
    ClkMux I__2161 (
            .O(N__9218),
            .I(N__9119));
    ClkMux I__2160 (
            .O(N__9217),
            .I(N__9119));
    ClkMux I__2159 (
            .O(N__9216),
            .I(N__9119));
    ClkMux I__2158 (
            .O(N__9215),
            .I(N__9119));
    ClkMux I__2157 (
            .O(N__9214),
            .I(N__9119));
    ClkMux I__2156 (
            .O(N__9213),
            .I(N__9119));
    ClkMux I__2155 (
            .O(N__9212),
            .I(N__9119));
    ClkMux I__2154 (
            .O(N__9211),
            .I(N__9119));
    ClkMux I__2153 (
            .O(N__9210),
            .I(N__9119));
    ClkMux I__2152 (
            .O(N__9209),
            .I(N__9119));
    ClkMux I__2151 (
            .O(N__9208),
            .I(N__9119));
    ClkMux I__2150 (
            .O(N__9207),
            .I(N__9119));
    ClkMux I__2149 (
            .O(N__9206),
            .I(N__9119));
    ClkMux I__2148 (
            .O(N__9205),
            .I(N__9119));
    ClkMux I__2147 (
            .O(N__9204),
            .I(N__9119));
    ClkMux I__2146 (
            .O(N__9203),
            .I(N__9119));
    ClkMux I__2145 (
            .O(N__9202),
            .I(N__9119));
    GlobalMux I__2144 (
            .O(N__9119),
            .I(CLK80_OUT));
    CEMux I__2143 (
            .O(N__9116),
            .I(N__9113));
    LocalMux I__2142 (
            .O(N__9113),
            .I(N__9109));
    CEMux I__2141 (
            .O(N__9112),
            .I(N__9105));
    Span4Mux_h I__2140 (
            .O(N__9109),
            .I(N__9102));
    CEMux I__2139 (
            .O(N__9108),
            .I(N__9099));
    LocalMux I__2138 (
            .O(N__9105),
            .I(N__9096));
    Odrv4 I__2137 (
            .O(N__9102),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    LocalMux I__2136 (
            .O(N__9099),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    Odrv12 I__2135 (
            .O(N__9096),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    InMux I__2134 (
            .O(N__9089),
            .I(N__9077));
    InMux I__2133 (
            .O(N__9088),
            .I(N__9072));
    InMux I__2132 (
            .O(N__9087),
            .I(N__9072));
    InMux I__2131 (
            .O(N__9086),
            .I(N__9069));
    InMux I__2130 (
            .O(N__9085),
            .I(N__9066));
    InMux I__2129 (
            .O(N__9084),
            .I(N__9063));
    InMux I__2128 (
            .O(N__9083),
            .I(N__9060));
    InMux I__2127 (
            .O(N__9082),
            .I(N__9057));
    InMux I__2126 (
            .O(N__9081),
            .I(N__9054));
    InMux I__2125 (
            .O(N__9080),
            .I(N__9051));
    LocalMux I__2124 (
            .O(N__9077),
            .I(N__9047));
    LocalMux I__2123 (
            .O(N__9072),
            .I(N__9043));
    LocalMux I__2122 (
            .O(N__9069),
            .I(N__9040));
    LocalMux I__2121 (
            .O(N__9066),
            .I(N__9037));
    LocalMux I__2120 (
            .O(N__9063),
            .I(N__9033));
    LocalMux I__2119 (
            .O(N__9060),
            .I(N__9015));
    LocalMux I__2118 (
            .O(N__9057),
            .I(N__9009));
    LocalMux I__2117 (
            .O(N__9054),
            .I(N__9000));
    LocalMux I__2116 (
            .O(N__9051),
            .I(N__8995));
    SRMux I__2115 (
            .O(N__9050),
            .I(N__8906));
    Glb2LocalMux I__2114 (
            .O(N__9047),
            .I(N__8906));
    SRMux I__2113 (
            .O(N__9046),
            .I(N__8906));
    Glb2LocalMux I__2112 (
            .O(N__9043),
            .I(N__8906));
    Glb2LocalMux I__2111 (
            .O(N__9040),
            .I(N__8906));
    Glb2LocalMux I__2110 (
            .O(N__9037),
            .I(N__8906));
    SRMux I__2109 (
            .O(N__9036),
            .I(N__8906));
    Glb2LocalMux I__2108 (
            .O(N__9033),
            .I(N__8906));
    SRMux I__2107 (
            .O(N__9032),
            .I(N__8906));
    SRMux I__2106 (
            .O(N__9031),
            .I(N__8906));
    SRMux I__2105 (
            .O(N__9030),
            .I(N__8906));
    SRMux I__2104 (
            .O(N__9029),
            .I(N__8906));
    SRMux I__2103 (
            .O(N__9028),
            .I(N__8906));
    SRMux I__2102 (
            .O(N__9027),
            .I(N__8906));
    SRMux I__2101 (
            .O(N__9026),
            .I(N__8906));
    SRMux I__2100 (
            .O(N__9025),
            .I(N__8906));
    SRMux I__2099 (
            .O(N__9024),
            .I(N__8906));
    SRMux I__2098 (
            .O(N__9023),
            .I(N__8906));
    SRMux I__2097 (
            .O(N__9022),
            .I(N__8906));
    SRMux I__2096 (
            .O(N__9021),
            .I(N__8906));
    SRMux I__2095 (
            .O(N__9020),
            .I(N__8906));
    SRMux I__2094 (
            .O(N__9019),
            .I(N__8906));
    SRMux I__2093 (
            .O(N__9018),
            .I(N__8906));
    Glb2LocalMux I__2092 (
            .O(N__9015),
            .I(N__8906));
    SRMux I__2091 (
            .O(N__9014),
            .I(N__8906));
    SRMux I__2090 (
            .O(N__9013),
            .I(N__8906));
    SRMux I__2089 (
            .O(N__9012),
            .I(N__8906));
    Glb2LocalMux I__2088 (
            .O(N__9009),
            .I(N__8906));
    SRMux I__2087 (
            .O(N__9008),
            .I(N__8906));
    SRMux I__2086 (
            .O(N__9007),
            .I(N__8906));
    SRMux I__2085 (
            .O(N__9006),
            .I(N__8906));
    SRMux I__2084 (
            .O(N__9005),
            .I(N__8906));
    SRMux I__2083 (
            .O(N__9004),
            .I(N__8906));
    SRMux I__2082 (
            .O(N__9003),
            .I(N__8906));
    Glb2LocalMux I__2081 (
            .O(N__9000),
            .I(N__8906));
    SRMux I__2080 (
            .O(N__8999),
            .I(N__8906));
    SRMux I__2079 (
            .O(N__8998),
            .I(N__8906));
    Glb2LocalMux I__2078 (
            .O(N__8995),
            .I(N__8906));
    SRMux I__2077 (
            .O(N__8994),
            .I(N__8906));
    SRMux I__2076 (
            .O(N__8993),
            .I(N__8906));
    SRMux I__2075 (
            .O(N__8992),
            .I(N__8906));
    SRMux I__2074 (
            .O(N__8991),
            .I(N__8906));
    GlobalMux I__2073 (
            .O(N__8906),
            .I(N__8903));
    gio2CtrlBuf I__2072 (
            .O(N__8903),
            .I(RESETn_c_i_g));
    CascadeMux I__2071 (
            .O(N__8900),
            .I(N__8897));
    InMux I__2070 (
            .O(N__8897),
            .I(N__8894));
    LocalMux I__2069 (
            .O(N__8894),
            .I(N__8889));
    InMux I__2068 (
            .O(N__8893),
            .I(N__8886));
    InMux I__2067 (
            .O(N__8892),
            .I(N__8883));
    Span4Mux_v I__2066 (
            .O(N__8889),
            .I(N__8878));
    LocalMux I__2065 (
            .O(N__8886),
            .I(N__8878));
    LocalMux I__2064 (
            .O(N__8883),
            .I(N__8875));
    Span4Mux_h I__2063 (
            .O(N__8878),
            .I(N__8870));
    Span4Mux_v I__2062 (
            .O(N__8875),
            .I(N__8870));
    Sp12to4 I__2061 (
            .O(N__8870),
            .I(N__8867));
    Span12Mux_v I__2060 (
            .O(N__8867),
            .I(N__8864));
    Span12Mux_h I__2059 (
            .O(N__8864),
            .I(N__8861));
    Odrv12 I__2058 (
            .O(N__8861),
            .I(CASLn_c));
    InMux I__2057 (
            .O(N__8858),
            .I(N__8854));
    InMux I__2056 (
            .O(N__8857),
            .I(N__8850));
    LocalMux I__2055 (
            .O(N__8854),
            .I(N__8847));
    InMux I__2054 (
            .O(N__8853),
            .I(N__8844));
    LocalMux I__2053 (
            .O(N__8850),
            .I(N__8841));
    Span4Mux_h I__2052 (
            .O(N__8847),
            .I(N__8836));
    LocalMux I__2051 (
            .O(N__8844),
            .I(N__8836));
    Span4Mux_v I__2050 (
            .O(N__8841),
            .I(N__8833));
    Span4Mux_v I__2049 (
            .O(N__8836),
            .I(N__8830));
    Span4Mux_v I__2048 (
            .O(N__8833),
            .I(N__8827));
    Sp12to4 I__2047 (
            .O(N__8830),
            .I(N__8822));
    Sp12to4 I__2046 (
            .O(N__8827),
            .I(N__8822));
    Span12Mux_h I__2045 (
            .O(N__8822),
            .I(N__8819));
    Span12Mux_v I__2044 (
            .O(N__8819),
            .I(N__8816));
    Odrv12 I__2043 (
            .O(N__8816),
            .I(CASUn_c));
    CascadeMux I__2042 (
            .O(N__8813),
            .I(N__8810));
    InMux I__2041 (
            .O(N__8810),
            .I(N__8807));
    LocalMux I__2040 (
            .O(N__8807),
            .I(N__8803));
    InMux I__2039 (
            .O(N__8806),
            .I(N__8799));
    Span4Mux_v I__2038 (
            .O(N__8803),
            .I(N__8796));
    InMux I__2037 (
            .O(N__8802),
            .I(N__8793));
    LocalMux I__2036 (
            .O(N__8799),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    Odrv4 I__2035 (
            .O(N__8796),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    LocalMux I__2034 (
            .O(N__8793),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__2033 (
            .O(N__8786),
            .I(N__8783));
    LocalMux I__2032 (
            .O(N__8783),
            .I(N__8780));
    Span4Mux_h I__2031 (
            .O(N__8780),
            .I(N__8776));
    InMux I__2030 (
            .O(N__8779),
            .I(N__8773));
    Odrv4 I__2029 (
            .O(N__8776),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__2028 (
            .O(N__8773),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__2027 (
            .O(N__8768),
            .I(N__8764));
    CascadeMux I__2026 (
            .O(N__8767),
            .I(N__8761));
    LocalMux I__2025 (
            .O(N__8764),
            .I(N__8750));
    InMux I__2024 (
            .O(N__8761),
            .I(N__8744));
    InMux I__2023 (
            .O(N__8760),
            .I(N__8744));
    InMux I__2022 (
            .O(N__8759),
            .I(N__8741));
    InMux I__2021 (
            .O(N__8758),
            .I(N__8736));
    InMux I__2020 (
            .O(N__8757),
            .I(N__8736));
    InMux I__2019 (
            .O(N__8756),
            .I(N__8731));
    InMux I__2018 (
            .O(N__8755),
            .I(N__8731));
    InMux I__2017 (
            .O(N__8754),
            .I(N__8728));
    InMux I__2016 (
            .O(N__8753),
            .I(N__8725));
    Span4Mux_h I__2015 (
            .O(N__8750),
            .I(N__8722));
    InMux I__2014 (
            .O(N__8749),
            .I(N__8719));
    LocalMux I__2013 (
            .O(N__8744),
            .I(N__8714));
    LocalMux I__2012 (
            .O(N__8741),
            .I(N__8709));
    LocalMux I__2011 (
            .O(N__8736),
            .I(N__8709));
    LocalMux I__2010 (
            .O(N__8731),
            .I(N__8706));
    LocalMux I__2009 (
            .O(N__8728),
            .I(N__8697));
    LocalMux I__2008 (
            .O(N__8725),
            .I(N__8697));
    Span4Mux_v I__2007 (
            .O(N__8722),
            .I(N__8697));
    LocalMux I__2006 (
            .O(N__8719),
            .I(N__8697));
    InMux I__2005 (
            .O(N__8718),
            .I(N__8693));
    InMux I__2004 (
            .O(N__8717),
            .I(N__8690));
    Span4Mux_v I__2003 (
            .O(N__8714),
            .I(N__8687));
    Span12Mux_h I__2002 (
            .O(N__8709),
            .I(N__8684));
    Span4Mux_h I__2001 (
            .O(N__8706),
            .I(N__8679));
    Span4Mux_h I__2000 (
            .O(N__8697),
            .I(N__8679));
    InMux I__1999 (
            .O(N__8696),
            .I(N__8676));
    LocalMux I__1998 (
            .O(N__8693),
            .I(N__8673));
    LocalMux I__1997 (
            .O(N__8690),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1996 (
            .O(N__8687),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv12 I__1995 (
            .O(N__8684),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1994 (
            .O(N__8679),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1993 (
            .O(N__8676),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1992 (
            .O(N__8673),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__1991 (
            .O(N__8660),
            .I(N__8657));
    LocalMux I__1990 (
            .O(N__8657),
            .I(N__8654));
    Span4Mux_s2_v I__1989 (
            .O(N__8654),
            .I(N__8651));
    Span4Mux_v I__1988 (
            .O(N__8651),
            .I(N__8648));
    Span4Mux_h I__1987 (
            .O(N__8648),
            .I(N__8645));
    Odrv4 I__1986 (
            .O(N__8645),
            .I(RASn_c));
    InMux I__1985 (
            .O(N__8642),
            .I(N__8635));
    CascadeMux I__1984 (
            .O(N__8641),
            .I(N__8632));
    CascadeMux I__1983 (
            .O(N__8640),
            .I(N__8628));
    CascadeMux I__1982 (
            .O(N__8639),
            .I(N__8624));
    CascadeMux I__1981 (
            .O(N__8638),
            .I(N__8621));
    LocalMux I__1980 (
            .O(N__8635),
            .I(N__8616));
    InMux I__1979 (
            .O(N__8632),
            .I(N__8609));
    InMux I__1978 (
            .O(N__8631),
            .I(N__8609));
    InMux I__1977 (
            .O(N__8628),
            .I(N__8604));
    InMux I__1976 (
            .O(N__8627),
            .I(N__8604));
    InMux I__1975 (
            .O(N__8624),
            .I(N__8597));
    InMux I__1974 (
            .O(N__8621),
            .I(N__8597));
    InMux I__1973 (
            .O(N__8620),
            .I(N__8597));
    InMux I__1972 (
            .O(N__8619),
            .I(N__8594));
    Span4Mux_h I__1971 (
            .O(N__8616),
            .I(N__8591));
    InMux I__1970 (
            .O(N__8615),
            .I(N__8586));
    InMux I__1969 (
            .O(N__8614),
            .I(N__8586));
    LocalMux I__1968 (
            .O(N__8609),
            .I(N__8583));
    LocalMux I__1967 (
            .O(N__8604),
            .I(N__8580));
    LocalMux I__1966 (
            .O(N__8597),
            .I(N__8577));
    LocalMux I__1965 (
            .O(N__8594),
            .I(N__8570));
    Span4Mux_v I__1964 (
            .O(N__8591),
            .I(N__8570));
    LocalMux I__1963 (
            .O(N__8586),
            .I(N__8570));
    Span4Mux_v I__1962 (
            .O(N__8583),
            .I(N__8563));
    Span4Mux_v I__1961 (
            .O(N__8580),
            .I(N__8563));
    Span4Mux_v I__1960 (
            .O(N__8577),
            .I(N__8560));
    Span4Mux_h I__1959 (
            .O(N__8570),
            .I(N__8557));
    InMux I__1958 (
            .O(N__8569),
            .I(N__8552));
    InMux I__1957 (
            .O(N__8568),
            .I(N__8552));
    Odrv4 I__1956 (
            .O(N__8563),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1955 (
            .O(N__8560),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1954 (
            .O(N__8557),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1953 (
            .O(N__8552),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1952 (
            .O(N__8543),
            .I(N__8540));
    LocalMux I__1951 (
            .O(N__8540),
            .I(N__8537));
    IoSpan4Mux I__1950 (
            .O(N__8537),
            .I(N__8534));
    IoSpan4Mux I__1949 (
            .O(N__8534),
            .I(N__8531));
    Span4Mux_s1_h I__1948 (
            .O(N__8531),
            .I(N__8528));
    Sp12to4 I__1947 (
            .O(N__8528),
            .I(N__8525));
    Odrv12 I__1946 (
            .O(N__8525),
            .I(WEn_c));
    InMux I__1945 (
            .O(N__8522),
            .I(N__8515));
    CascadeMux I__1944 (
            .O(N__8521),
            .I(N__8511));
    InMux I__1943 (
            .O(N__8520),
            .I(N__8508));
    InMux I__1942 (
            .O(N__8519),
            .I(N__8497));
    InMux I__1941 (
            .O(N__8518),
            .I(N__8497));
    LocalMux I__1940 (
            .O(N__8515),
            .I(N__8493));
    CascadeMux I__1939 (
            .O(N__8514),
            .I(N__8490));
    InMux I__1938 (
            .O(N__8511),
            .I(N__8487));
    LocalMux I__1937 (
            .O(N__8508),
            .I(N__8484));
    InMux I__1936 (
            .O(N__8507),
            .I(N__8481));
    InMux I__1935 (
            .O(N__8506),
            .I(N__8477));
    InMux I__1934 (
            .O(N__8505),
            .I(N__8472));
    InMux I__1933 (
            .O(N__8504),
            .I(N__8472));
    InMux I__1932 (
            .O(N__8503),
            .I(N__8465));
    InMux I__1931 (
            .O(N__8502),
            .I(N__8465));
    LocalMux I__1930 (
            .O(N__8497),
            .I(N__8462));
    InMux I__1929 (
            .O(N__8496),
            .I(N__8459));
    Span4Mux_v I__1928 (
            .O(N__8493),
            .I(N__8456));
    InMux I__1927 (
            .O(N__8490),
            .I(N__8453));
    LocalMux I__1926 (
            .O(N__8487),
            .I(N__8446));
    Span4Mux_h I__1925 (
            .O(N__8484),
            .I(N__8446));
    LocalMux I__1924 (
            .O(N__8481),
            .I(N__8446));
    InMux I__1923 (
            .O(N__8480),
            .I(N__8443));
    LocalMux I__1922 (
            .O(N__8477),
            .I(N__8438));
    LocalMux I__1921 (
            .O(N__8472),
            .I(N__8438));
    InMux I__1920 (
            .O(N__8471),
            .I(N__8435));
    CascadeMux I__1919 (
            .O(N__8470),
            .I(N__8432));
    LocalMux I__1918 (
            .O(N__8465),
            .I(N__8429));
    Span4Mux_v I__1917 (
            .O(N__8462),
            .I(N__8420));
    LocalMux I__1916 (
            .O(N__8459),
            .I(N__8420));
    Span4Mux_h I__1915 (
            .O(N__8456),
            .I(N__8420));
    LocalMux I__1914 (
            .O(N__8453),
            .I(N__8420));
    Span4Mux_v I__1913 (
            .O(N__8446),
            .I(N__8417));
    LocalMux I__1912 (
            .O(N__8443),
            .I(N__8410));
    Span4Mux_v I__1911 (
            .O(N__8438),
            .I(N__8410));
    LocalMux I__1910 (
            .O(N__8435),
            .I(N__8410));
    InMux I__1909 (
            .O(N__8432),
            .I(N__8407));
    Odrv4 I__1908 (
            .O(N__8429),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1907 (
            .O(N__8420),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1906 (
            .O(N__8417),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1905 (
            .O(N__8410),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1904 (
            .O(N__8407),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    IoInMux I__1903 (
            .O(N__8396),
            .I(N__8393));
    LocalMux I__1902 (
            .O(N__8393),
            .I(N__8390));
    Span4Mux_s1_v I__1901 (
            .O(N__8390),
            .I(N__8387));
    Sp12to4 I__1900 (
            .O(N__8387),
            .I(N__8384));
    Span12Mux_h I__1899 (
            .O(N__8384),
            .I(N__8381));
    Odrv12 I__1898 (
            .O(N__8381),
            .I(CASn_c));
    InMux I__1897 (
            .O(N__8378),
            .I(N__8374));
    InMux I__1896 (
            .O(N__8377),
            .I(N__8371));
    LocalMux I__1895 (
            .O(N__8374),
            .I(N__8368));
    LocalMux I__1894 (
            .O(N__8371),
            .I(N__8365));
    Span4Mux_v I__1893 (
            .O(N__8368),
            .I(N__8362));
    Span4Mux_h I__1892 (
            .O(N__8365),
            .I(N__8359));
    Span4Mux_v I__1891 (
            .O(N__8362),
            .I(N__8356));
    Span4Mux_v I__1890 (
            .O(N__8359),
            .I(N__8353));
    Sp12to4 I__1889 (
            .O(N__8356),
            .I(N__8348));
    Sp12to4 I__1888 (
            .O(N__8353),
            .I(N__8348));
    Span12Mux_h I__1887 (
            .O(N__8348),
            .I(N__8345));
    Odrv12 I__1886 (
            .O(N__8345),
            .I(RAS0n_c));
    InMux I__1885 (
            .O(N__8342),
            .I(N__8339));
    LocalMux I__1884 (
            .O(N__8339),
            .I(N__8336));
    Span12Mux_v I__1883 (
            .O(N__8336),
            .I(N__8333));
    Span12Mux_h I__1882 (
            .O(N__8333),
            .I(N__8330));
    Odrv12 I__1881 (
            .O(N__8330),
            .I(RAS1n_c));
    InMux I__1880 (
            .O(N__8327),
            .I(N__8323));
    InMux I__1879 (
            .O(N__8326),
            .I(N__8320));
    LocalMux I__1878 (
            .O(N__8323),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    LocalMux I__1877 (
            .O(N__8320),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__1876 (
            .O(N__8315),
            .I(N__8312));
    LocalMux I__1875 (
            .O(N__8312),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    InMux I__1874 (
            .O(N__8309),
            .I(N__8305));
    InMux I__1873 (
            .O(N__8308),
            .I(N__8302));
    LocalMux I__1872 (
            .O(N__8305),
            .I(N__8299));
    LocalMux I__1871 (
            .O(N__8302),
            .I(N__8296));
    Span4Mux_v I__1870 (
            .O(N__8299),
            .I(N__8293));
    Span4Mux_v I__1869 (
            .O(N__8296),
            .I(N__8290));
    Span4Mux_v I__1868 (
            .O(N__8293),
            .I(N__8287));
    Span4Mux_v I__1867 (
            .O(N__8290),
            .I(N__8284));
    Sp12to4 I__1866 (
            .O(N__8287),
            .I(N__8279));
    Sp12to4 I__1865 (
            .O(N__8284),
            .I(N__8279));
    Span12Mux_h I__1864 (
            .O(N__8279),
            .I(N__8276));
    Odrv12 I__1863 (
            .O(N__8276),
            .I(DRA_c_7));
    InMux I__1862 (
            .O(N__8273),
            .I(N__8270));
    LocalMux I__1861 (
            .O(N__8270),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__1860 (
            .O(N__8267),
            .I(N__8264));
    LocalMux I__1859 (
            .O(N__8264),
            .I(N__8261));
    Sp12to4 I__1858 (
            .O(N__8261),
            .I(N__8258));
    Span12Mux_v I__1857 (
            .O(N__8258),
            .I(N__8255));
    Span12Mux_h I__1856 (
            .O(N__8255),
            .I(N__8252));
    Odrv12 I__1855 (
            .O(N__8252),
            .I(A_c_18));
    CascadeMux I__1854 (
            .O(N__8249),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_ ));
    InMux I__1853 (
            .O(N__8246),
            .I(N__8243));
    LocalMux I__1852 (
            .O(N__8243),
            .I(N__8240));
    Sp12to4 I__1851 (
            .O(N__8240),
            .I(N__8237));
    Span12Mux_v I__1850 (
            .O(N__8237),
            .I(N__8234));
    Span12Mux_h I__1849 (
            .O(N__8234),
            .I(N__8231));
    Odrv12 I__1848 (
            .O(N__8231),
            .I(A_c_16));
    CascadeMux I__1847 (
            .O(N__8228),
            .I(\U712_CHIP_RAM.N_322_cascade_ ));
    IoInMux I__1846 (
            .O(N__8225),
            .I(N__8222));
    LocalMux I__1845 (
            .O(N__8222),
            .I(N__8219));
    Span4Mux_s2_h I__1844 (
            .O(N__8219),
            .I(N__8216));
    Span4Mux_v I__1843 (
            .O(N__8216),
            .I(N__8213));
    Sp12to4 I__1842 (
            .O(N__8213),
            .I(N__8210));
    Span12Mux_h I__1841 (
            .O(N__8210),
            .I(N__8207));
    Odrv12 I__1840 (
            .O(N__8207),
            .I(CMA_c_7));
    InMux I__1839 (
            .O(N__8204),
            .I(N__8201));
    LocalMux I__1838 (
            .O(N__8201),
            .I(\U712_CHIP_RAM.CMA_5_i_0_8 ));
    InMux I__1837 (
            .O(N__8198),
            .I(N__8195));
    LocalMux I__1836 (
            .O(N__8195),
            .I(N__8192));
    Span4Mux_v I__1835 (
            .O(N__8192),
            .I(N__8189));
    Span4Mux_v I__1834 (
            .O(N__8189),
            .I(N__8186));
    Sp12to4 I__1833 (
            .O(N__8186),
            .I(N__8183));
    Span12Mux_h I__1832 (
            .O(N__8183),
            .I(N__8180));
    Odrv12 I__1831 (
            .O(N__8180),
            .I(A_c_19));
    CascadeMux I__1830 (
            .O(N__8177),
            .I(\U712_CHIP_RAM.CMA_5_i_0_8_cascade_ ));
    CascadeMux I__1829 (
            .O(N__8174),
            .I(N__8170));
    CascadeMux I__1828 (
            .O(N__8173),
            .I(N__8163));
    InMux I__1827 (
            .O(N__8170),
            .I(N__8159));
    CascadeMux I__1826 (
            .O(N__8169),
            .I(N__8155));
    CascadeMux I__1825 (
            .O(N__8168),
            .I(N__8152));
    InMux I__1824 (
            .O(N__8167),
            .I(N__8141));
    InMux I__1823 (
            .O(N__8166),
            .I(N__8141));
    InMux I__1822 (
            .O(N__8163),
            .I(N__8138));
    InMux I__1821 (
            .O(N__8162),
            .I(N__8129));
    LocalMux I__1820 (
            .O(N__8159),
            .I(N__8126));
    InMux I__1819 (
            .O(N__8158),
            .I(N__8123));
    InMux I__1818 (
            .O(N__8155),
            .I(N__8120));
    InMux I__1817 (
            .O(N__8152),
            .I(N__8115));
    InMux I__1816 (
            .O(N__8151),
            .I(N__8115));
    InMux I__1815 (
            .O(N__8150),
            .I(N__8108));
    InMux I__1814 (
            .O(N__8149),
            .I(N__8108));
    InMux I__1813 (
            .O(N__8148),
            .I(N__8108));
    CascadeMux I__1812 (
            .O(N__8147),
            .I(N__8103));
    CascadeMux I__1811 (
            .O(N__8146),
            .I(N__8100));
    LocalMux I__1810 (
            .O(N__8141),
            .I(N__8094));
    LocalMux I__1809 (
            .O(N__8138),
            .I(N__8094));
    InMux I__1808 (
            .O(N__8137),
            .I(N__8089));
    InMux I__1807 (
            .O(N__8136),
            .I(N__8086));
    InMux I__1806 (
            .O(N__8135),
            .I(N__8081));
    InMux I__1805 (
            .O(N__8134),
            .I(N__8081));
    CascadeMux I__1804 (
            .O(N__8133),
            .I(N__8077));
    InMux I__1803 (
            .O(N__8132),
            .I(N__8073));
    LocalMux I__1802 (
            .O(N__8129),
            .I(N__8064));
    Span4Mux_v I__1801 (
            .O(N__8126),
            .I(N__8064));
    LocalMux I__1800 (
            .O(N__8123),
            .I(N__8064));
    LocalMux I__1799 (
            .O(N__8120),
            .I(N__8064));
    LocalMux I__1798 (
            .O(N__8115),
            .I(N__8056));
    LocalMux I__1797 (
            .O(N__8108),
            .I(N__8056));
    InMux I__1796 (
            .O(N__8107),
            .I(N__8051));
    InMux I__1795 (
            .O(N__8106),
            .I(N__8051));
    InMux I__1794 (
            .O(N__8103),
            .I(N__8046));
    InMux I__1793 (
            .O(N__8100),
            .I(N__8046));
    InMux I__1792 (
            .O(N__8099),
            .I(N__8043));
    Span4Mux_h I__1791 (
            .O(N__8094),
            .I(N__8040));
    InMux I__1790 (
            .O(N__8093),
            .I(N__8035));
    InMux I__1789 (
            .O(N__8092),
            .I(N__8035));
    LocalMux I__1788 (
            .O(N__8089),
            .I(N__8028));
    LocalMux I__1787 (
            .O(N__8086),
            .I(N__8028));
    LocalMux I__1786 (
            .O(N__8081),
            .I(N__8028));
    InMux I__1785 (
            .O(N__8080),
            .I(N__8021));
    InMux I__1784 (
            .O(N__8077),
            .I(N__8021));
    InMux I__1783 (
            .O(N__8076),
            .I(N__8021));
    LocalMux I__1782 (
            .O(N__8073),
            .I(N__8016));
    Span4Mux_h I__1781 (
            .O(N__8064),
            .I(N__8016));
    InMux I__1780 (
            .O(N__8063),
            .I(N__8009));
    InMux I__1779 (
            .O(N__8062),
            .I(N__8009));
    InMux I__1778 (
            .O(N__8061),
            .I(N__8009));
    Odrv12 I__1777 (
            .O(N__8056),
            .I(CPU_CYCLEm));
    LocalMux I__1776 (
            .O(N__8051),
            .I(CPU_CYCLEm));
    LocalMux I__1775 (
            .O(N__8046),
            .I(CPU_CYCLEm));
    LocalMux I__1774 (
            .O(N__8043),
            .I(CPU_CYCLEm));
    Odrv4 I__1773 (
            .O(N__8040),
            .I(CPU_CYCLEm));
    LocalMux I__1772 (
            .O(N__8035),
            .I(CPU_CYCLEm));
    Odrv12 I__1771 (
            .O(N__8028),
            .I(CPU_CYCLEm));
    LocalMux I__1770 (
            .O(N__8021),
            .I(CPU_CYCLEm));
    Odrv4 I__1769 (
            .O(N__8016),
            .I(CPU_CYCLEm));
    LocalMux I__1768 (
            .O(N__8009),
            .I(CPU_CYCLEm));
    IoInMux I__1767 (
            .O(N__7988),
            .I(N__7985));
    LocalMux I__1766 (
            .O(N__7985),
            .I(N__7982));
    IoSpan4Mux I__1765 (
            .O(N__7982),
            .I(N__7979));
    Span4Mux_s2_h I__1764 (
            .O(N__7979),
            .I(N__7976));
    Sp12to4 I__1763 (
            .O(N__7976),
            .I(N__7973));
    Span12Mux_h I__1762 (
            .O(N__7973),
            .I(N__7970));
    Odrv12 I__1761 (
            .O(N__7970),
            .I(CMA_c_9));
    CEMux I__1760 (
            .O(N__7967),
            .I(N__7961));
    CEMux I__1759 (
            .O(N__7966),
            .I(N__7958));
    CEMux I__1758 (
            .O(N__7965),
            .I(N__7955));
    CEMux I__1757 (
            .O(N__7964),
            .I(N__7952));
    LocalMux I__1756 (
            .O(N__7961),
            .I(N__7948));
    LocalMux I__1755 (
            .O(N__7958),
            .I(N__7945));
    LocalMux I__1754 (
            .O(N__7955),
            .I(N__7942));
    LocalMux I__1753 (
            .O(N__7952),
            .I(N__7939));
    CEMux I__1752 (
            .O(N__7951),
            .I(N__7936));
    Span4Mux_h I__1751 (
            .O(N__7948),
            .I(N__7931));
    Span4Mux_h I__1750 (
            .O(N__7945),
            .I(N__7931));
    Span4Mux_v I__1749 (
            .O(N__7942),
            .I(N__7928));
    Span4Mux_v I__1748 (
            .O(N__7939),
            .I(N__7923));
    LocalMux I__1747 (
            .O(N__7936),
            .I(N__7923));
    Odrv4 I__1746 (
            .O(N__7931),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv4 I__1745 (
            .O(N__7928),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv4 I__1744 (
            .O(N__7923),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    InMux I__1743 (
            .O(N__7916),
            .I(N__7913));
    LocalMux I__1742 (
            .O(N__7913),
            .I(N__7910));
    Odrv12 I__1741 (
            .O(N__7910),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1740 (
            .O(N__7907),
            .I(N__7903));
    InMux I__1739 (
            .O(N__7906),
            .I(N__7900));
    LocalMux I__1738 (
            .O(N__7903),
            .I(N__7895));
    LocalMux I__1737 (
            .O(N__7900),
            .I(N__7895));
    Span4Mux_v I__1736 (
            .O(N__7895),
            .I(N__7892));
    Sp12to4 I__1735 (
            .O(N__7892),
            .I(N__7889));
    Span12Mux_h I__1734 (
            .O(N__7889),
            .I(N__7886));
    Span12Mux_v I__1733 (
            .O(N__7886),
            .I(N__7883));
    Odrv12 I__1732 (
            .O(N__7883),
            .I(DRA_c_4));
    InMux I__1731 (
            .O(N__7880),
            .I(N__7877));
    LocalMux I__1730 (
            .O(N__7877),
            .I(N__7874));
    Odrv12 I__1729 (
            .O(N__7874),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__1728 (
            .O(N__7871),
            .I(N__7868));
    LocalMux I__1727 (
            .O(N__7868),
            .I(N__7864));
    InMux I__1726 (
            .O(N__7867),
            .I(N__7861));
    Span4Mux_v I__1725 (
            .O(N__7864),
            .I(N__7856));
    LocalMux I__1724 (
            .O(N__7861),
            .I(N__7856));
    Span4Mux_v I__1723 (
            .O(N__7856),
            .I(N__7853));
    Sp12to4 I__1722 (
            .O(N__7853),
            .I(N__7850));
    Span12Mux_h I__1721 (
            .O(N__7850),
            .I(N__7847));
    Odrv12 I__1720 (
            .O(N__7847),
            .I(DRA_c_8));
    InMux I__1719 (
            .O(N__7844),
            .I(N__7841));
    LocalMux I__1718 (
            .O(N__7841),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    CEMux I__1717 (
            .O(N__7838),
            .I(N__7834));
    CEMux I__1716 (
            .O(N__7837),
            .I(N__7829));
    LocalMux I__1715 (
            .O(N__7834),
            .I(N__7826));
    CEMux I__1714 (
            .O(N__7833),
            .I(N__7823));
    CEMux I__1713 (
            .O(N__7832),
            .I(N__7820));
    LocalMux I__1712 (
            .O(N__7829),
            .I(N__7817));
    Span4Mux_v I__1711 (
            .O(N__7826),
            .I(N__7814));
    LocalMux I__1710 (
            .O(N__7823),
            .I(N__7809));
    LocalMux I__1709 (
            .O(N__7820),
            .I(N__7809));
    Span4Mux_h I__1708 (
            .O(N__7817),
            .I(N__7804));
    Span4Mux_h I__1707 (
            .O(N__7814),
            .I(N__7804));
    Span4Mux_v I__1706 (
            .O(N__7809),
            .I(N__7801));
    Odrv4 I__1705 (
            .O(N__7804),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    Odrv4 I__1704 (
            .O(N__7801),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    InMux I__1703 (
            .O(N__7796),
            .I(N__7791));
    InMux I__1702 (
            .O(N__7795),
            .I(N__7786));
    InMux I__1701 (
            .O(N__7794),
            .I(N__7786));
    LocalMux I__1700 (
            .O(N__7791),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__1699 (
            .O(N__7786),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__1698 (
            .O(N__7781),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__1697 (
            .O(N__7778),
            .I(N__7774));
    InMux I__1696 (
            .O(N__7777),
            .I(N__7771));
    LocalMux I__1695 (
            .O(N__7774),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__1694 (
            .O(N__7771),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__1693 (
            .O(N__7766),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__1692 (
            .O(N__7763),
            .I(N__7759));
    InMux I__1691 (
            .O(N__7762),
            .I(N__7756));
    LocalMux I__1690 (
            .O(N__7759),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__1689 (
            .O(N__7756),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__1688 (
            .O(N__7751),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__1687 (
            .O(N__7748),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    InMux I__1686 (
            .O(N__7745),
            .I(N__7740));
    InMux I__1685 (
            .O(N__7744),
            .I(N__7735));
    InMux I__1684 (
            .O(N__7743),
            .I(N__7735));
    LocalMux I__1683 (
            .O(N__7740),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__1682 (
            .O(N__7735),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    ClkMux I__1681 (
            .O(N__7730),
            .I(N__7727));
    GlobalMux I__1680 (
            .O(N__7727),
            .I(N__7724));
    gio2CtrlBuf I__1679 (
            .O(N__7724),
            .I(C1_c_g));
    SRMux I__1678 (
            .O(N__7721),
            .I(N__7718));
    LocalMux I__1677 (
            .O(N__7718),
            .I(N__7715));
    Span4Mux_h I__1676 (
            .O(N__7715),
            .I(N__7712));
    Odrv4 I__1675 (
            .O(N__7712),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__1674 (
            .O(N__7709),
            .I(N__7703));
    InMux I__1673 (
            .O(N__7708),
            .I(N__7703));
    LocalMux I__1672 (
            .O(N__7703),
            .I(N__7698));
    InMux I__1671 (
            .O(N__7702),
            .I(N__7695));
    InMux I__1670 (
            .O(N__7701),
            .I(N__7692));
    Span4Mux_v I__1669 (
            .O(N__7698),
            .I(N__7686));
    LocalMux I__1668 (
            .O(N__7695),
            .I(N__7686));
    LocalMux I__1667 (
            .O(N__7692),
            .I(N__7682));
    InMux I__1666 (
            .O(N__7691),
            .I(N__7679));
    Span4Mux_h I__1665 (
            .O(N__7686),
            .I(N__7676));
    InMux I__1664 (
            .O(N__7685),
            .I(N__7673));
    Span4Mux_v I__1663 (
            .O(N__7682),
            .I(N__7670));
    LocalMux I__1662 (
            .O(N__7679),
            .I(N__7667));
    Span4Mux_v I__1661 (
            .O(N__7676),
            .I(N__7664));
    LocalMux I__1660 (
            .O(N__7673),
            .I(N__7661));
    Sp12to4 I__1659 (
            .O(N__7670),
            .I(N__7658));
    Span12Mux_h I__1658 (
            .O(N__7667),
            .I(N__7655));
    Sp12to4 I__1657 (
            .O(N__7664),
            .I(N__7650));
    Span12Mux_v I__1656 (
            .O(N__7661),
            .I(N__7650));
    Span12Mux_h I__1655 (
            .O(N__7658),
            .I(N__7647));
    Span12Mux_h I__1654 (
            .O(N__7655),
            .I(N__7644));
    Span12Mux_h I__1653 (
            .O(N__7650),
            .I(N__7641));
    Odrv12 I__1652 (
            .O(N__7647),
            .I(RESETn_c));
    Odrv12 I__1651 (
            .O(N__7644),
            .I(RESETn_c));
    Odrv12 I__1650 (
            .O(N__7641),
            .I(RESETn_c));
    IoInMux I__1649 (
            .O(N__7634),
            .I(N__7631));
    LocalMux I__1648 (
            .O(N__7631),
            .I(N__7628));
    Span12Mux_s7_v I__1647 (
            .O(N__7628),
            .I(N__7625));
    Odrv12 I__1646 (
            .O(N__7625),
            .I(RESETn_c_i));
    InMux I__1645 (
            .O(N__7622),
            .I(N__7619));
    LocalMux I__1644 (
            .O(N__7619),
            .I(N__7615));
    InMux I__1643 (
            .O(N__7618),
            .I(N__7612));
    Span4Mux_h I__1642 (
            .O(N__7615),
            .I(N__7609));
    LocalMux I__1641 (
            .O(N__7612),
            .I(N__7606));
    Sp12to4 I__1640 (
            .O(N__7609),
            .I(N__7601));
    Sp12to4 I__1639 (
            .O(N__7606),
            .I(N__7601));
    Span12Mux_v I__1638 (
            .O(N__7601),
            .I(N__7598));
    Span12Mux_h I__1637 (
            .O(N__7598),
            .I(N__7595));
    Odrv12 I__1636 (
            .O(N__7595),
            .I(DRA_c_5));
    InMux I__1635 (
            .O(N__7592),
            .I(N__7589));
    LocalMux I__1634 (
            .O(N__7589),
            .I(N__7586));
    Odrv4 I__1633 (
            .O(N__7586),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1632 (
            .O(N__7583),
            .I(N__7580));
    LocalMux I__1631 (
            .O(N__7580),
            .I(N__7577));
    Odrv12 I__1630 (
            .O(N__7577),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    CascadeMux I__1629 (
            .O(N__7574),
            .I(N__7571));
    InMux I__1628 (
            .O(N__7571),
            .I(N__7568));
    LocalMux I__1627 (
            .O(N__7568),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__1626 (
            .O(N__7565),
            .I(N__7561));
    InMux I__1625 (
            .O(N__7564),
            .I(N__7558));
    LocalMux I__1624 (
            .O(N__7561),
            .I(N__7553));
    LocalMux I__1623 (
            .O(N__7558),
            .I(N__7553));
    Span4Mux_v I__1622 (
            .O(N__7553),
            .I(N__7550));
    Sp12to4 I__1621 (
            .O(N__7550),
            .I(N__7547));
    Span12Mux_h I__1620 (
            .O(N__7547),
            .I(N__7544));
    Span12Mux_v I__1619 (
            .O(N__7544),
            .I(N__7541));
    Odrv12 I__1618 (
            .O(N__7541),
            .I(DRA_c_6));
    InMux I__1617 (
            .O(N__7538),
            .I(N__7535));
    LocalMux I__1616 (
            .O(N__7535),
            .I(N__7532));
    Odrv4 I__1615 (
            .O(N__7532),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__1614 (
            .O(N__7529),
            .I(N__7526));
    LocalMux I__1613 (
            .O(N__7526),
            .I(N__7522));
    InMux I__1612 (
            .O(N__7525),
            .I(N__7519));
    Span4Mux_h I__1611 (
            .O(N__7522),
            .I(N__7514));
    LocalMux I__1610 (
            .O(N__7519),
            .I(N__7514));
    Span4Mux_v I__1609 (
            .O(N__7514),
            .I(N__7511));
    Sp12to4 I__1608 (
            .O(N__7511),
            .I(N__7508));
    Span12Mux_h I__1607 (
            .O(N__7508),
            .I(N__7505));
    Span12Mux_v I__1606 (
            .O(N__7505),
            .I(N__7502));
    Odrv12 I__1605 (
            .O(N__7502),
            .I(DRA_c_1));
    InMux I__1604 (
            .O(N__7499),
            .I(N__7496));
    LocalMux I__1603 (
            .O(N__7496),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__1602 (
            .O(N__7493),
            .I(N__7490));
    LocalMux I__1601 (
            .O(N__7490),
            .I(N__7486));
    InMux I__1600 (
            .O(N__7489),
            .I(N__7483));
    Span4Mux_v I__1599 (
            .O(N__7486),
            .I(N__7480));
    LocalMux I__1598 (
            .O(N__7483),
            .I(N__7475));
    Sp12to4 I__1597 (
            .O(N__7480),
            .I(N__7475));
    Span12Mux_h I__1596 (
            .O(N__7475),
            .I(N__7472));
    Span12Mux_v I__1595 (
            .O(N__7472),
            .I(N__7469));
    Odrv12 I__1594 (
            .O(N__7469),
            .I(DRA_c_3));
    InMux I__1593 (
            .O(N__7466),
            .I(N__7463));
    LocalMux I__1592 (
            .O(N__7463),
            .I(N__7460));
    Odrv12 I__1591 (
            .O(N__7460),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__1590 (
            .O(N__7457),
            .I(N__7454));
    LocalMux I__1589 (
            .O(N__7454),
            .I(N__7450));
    InMux I__1588 (
            .O(N__7453),
            .I(N__7447));
    Span4Mux_v I__1587 (
            .O(N__7450),
            .I(N__7444));
    LocalMux I__1586 (
            .O(N__7447),
            .I(N__7441));
    Sp12to4 I__1585 (
            .O(N__7444),
            .I(N__7438));
    Span12Mux_h I__1584 (
            .O(N__7441),
            .I(N__7435));
    Span12Mux_h I__1583 (
            .O(N__7438),
            .I(N__7432));
    Span12Mux_v I__1582 (
            .O(N__7435),
            .I(N__7429));
    Span12Mux_v I__1581 (
            .O(N__7432),
            .I(N__7426));
    Odrv12 I__1580 (
            .O(N__7429),
            .I(DRA_c_2));
    Odrv12 I__1579 (
            .O(N__7426),
            .I(DRA_c_2));
    CascadeMux I__1578 (
            .O(N__7421),
            .I(N__7418));
    InMux I__1577 (
            .O(N__7418),
            .I(N__7415));
    LocalMux I__1576 (
            .O(N__7415),
            .I(N__7412));
    Odrv4 I__1575 (
            .O(N__7412),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    IoInMux I__1574 (
            .O(N__7409),
            .I(N__7406));
    LocalMux I__1573 (
            .O(N__7406),
            .I(N__7403));
    Span4Mux_s3_v I__1572 (
            .O(N__7403),
            .I(N__7400));
    Span4Mux_v I__1571 (
            .O(N__7400),
            .I(N__7397));
    Span4Mux_v I__1570 (
            .O(N__7397),
            .I(N__7394));
    Span4Mux_h I__1569 (
            .O(N__7394),
            .I(N__7390));
    InMux I__1568 (
            .O(N__7393),
            .I(N__7387));
    Odrv4 I__1567 (
            .O(N__7390),
            .I(CONSTANT_ONE_NET));
    LocalMux I__1566 (
            .O(N__7387),
            .I(CONSTANT_ONE_NET));
    InMux I__1565 (
            .O(N__7382),
            .I(N__7379));
    LocalMux I__1564 (
            .O(N__7379),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ));
    InMux I__1563 (
            .O(N__7376),
            .I(bfn_12_8_0_));
    InMux I__1562 (
            .O(N__7373),
            .I(N__7370));
    LocalMux I__1561 (
            .O(N__7370),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__1560 (
            .O(N__7367),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__1559 (
            .O(N__7364),
            .I(N__7359));
    InMux I__1558 (
            .O(N__7363),
            .I(N__7354));
    InMux I__1557 (
            .O(N__7362),
            .I(N__7354));
    LocalMux I__1556 (
            .O(N__7359),
            .I(\U712_CHIP_RAM.REFRESH9lto2 ));
    LocalMux I__1555 (
            .O(N__7354),
            .I(\U712_CHIP_RAM.REFRESH9lto2 ));
    InMux I__1554 (
            .O(N__7349),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    CascadeMux I__1553 (
            .O(N__7346),
            .I(N__7342));
    InMux I__1552 (
            .O(N__7345),
            .I(N__7338));
    InMux I__1551 (
            .O(N__7342),
            .I(N__7333));
    InMux I__1550 (
            .O(N__7341),
            .I(N__7333));
    LocalMux I__1549 (
            .O(N__7338),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__1548 (
            .O(N__7333),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__1547 (
            .O(N__7328),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__1546 (
            .O(N__7325),
            .I(N__7322));
    LocalMux I__1545 (
            .O(N__7322),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1544 (
            .O(N__7319),
            .I(N__7316));
    LocalMux I__1543 (
            .O(N__7316),
            .I(\U712_CHIP_RAM.N_321 ));
    IoInMux I__1542 (
            .O(N__7313),
            .I(N__7310));
    LocalMux I__1541 (
            .O(N__7310),
            .I(N__7307));
    Span4Mux_s0_h I__1540 (
            .O(N__7307),
            .I(N__7304));
    Sp12to4 I__1539 (
            .O(N__7304),
            .I(N__7301));
    Span12Mux_s9_v I__1538 (
            .O(N__7301),
            .I(N__7298));
    Span12Mux_h I__1537 (
            .O(N__7298),
            .I(N__7295));
    Odrv12 I__1536 (
            .O(N__7295),
            .I(CMA_c_6));
    InMux I__1535 (
            .O(N__7292),
            .I(N__7289));
    LocalMux I__1534 (
            .O(N__7289),
            .I(\U712_CHIP_RAM.N_320 ));
    IoInMux I__1533 (
            .O(N__7286),
            .I(N__7283));
    LocalMux I__1532 (
            .O(N__7283),
            .I(N__7280));
    Span12Mux_s4_h I__1531 (
            .O(N__7280),
            .I(N__7277));
    Span12Mux_h I__1530 (
            .O(N__7277),
            .I(N__7274));
    Odrv12 I__1529 (
            .O(N__7274),
            .I(CMA_c_5));
    InMux I__1528 (
            .O(N__7271),
            .I(N__7268));
    LocalMux I__1527 (
            .O(N__7268),
            .I(N__7265));
    Span12Mux_v I__1526 (
            .O(N__7265),
            .I(N__7262));
    Span12Mux_h I__1525 (
            .O(N__7262),
            .I(N__7259));
    Odrv12 I__1524 (
            .O(N__7259),
            .I(A_c_17));
    IoInMux I__1523 (
            .O(N__7256),
            .I(N__7253));
    LocalMux I__1522 (
            .O(N__7253),
            .I(N__7250));
    Span12Mux_s4_h I__1521 (
            .O(N__7250),
            .I(N__7247));
    Span12Mux_h I__1520 (
            .O(N__7247),
            .I(N__7244));
    Odrv12 I__1519 (
            .O(N__7244),
            .I(CMA_c_8));
    InMux I__1518 (
            .O(N__7241),
            .I(N__7238));
    LocalMux I__1517 (
            .O(N__7238),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__1516 (
            .O(N__7235),
            .I(N__7232));
    LocalMux I__1515 (
            .O(N__7232),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__1514 (
            .O(N__7229),
            .I(N__7226));
    LocalMux I__1513 (
            .O(N__7226),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1512 (
            .O(N__7223),
            .I(N__7220));
    LocalMux I__1511 (
            .O(N__7220),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__1510 (
            .O(N__7217),
            .I(N__7213));
    InMux I__1509 (
            .O(N__7216),
            .I(N__7210));
    LocalMux I__1508 (
            .O(N__7213),
            .I(\U712_CHIP_RAM.N_425 ));
    LocalMux I__1507 (
            .O(N__7210),
            .I(\U712_CHIP_RAM.N_425 ));
    InMux I__1506 (
            .O(N__7205),
            .I(N__7200));
    InMux I__1505 (
            .O(N__7204),
            .I(N__7197));
    InMux I__1504 (
            .O(N__7203),
            .I(N__7194));
    LocalMux I__1503 (
            .O(N__7200),
            .I(N__7190));
    LocalMux I__1502 (
            .O(N__7197),
            .I(N__7185));
    LocalMux I__1501 (
            .O(N__7194),
            .I(N__7182));
    InMux I__1500 (
            .O(N__7193),
            .I(N__7174));
    Span4Mux_v I__1499 (
            .O(N__7190),
            .I(N__7171));
    InMux I__1498 (
            .O(N__7189),
            .I(N__7168));
    InMux I__1497 (
            .O(N__7188),
            .I(N__7165));
    Span4Mux_v I__1496 (
            .O(N__7185),
            .I(N__7160));
    Span4Mux_v I__1495 (
            .O(N__7182),
            .I(N__7160));
    InMux I__1494 (
            .O(N__7181),
            .I(N__7155));
    InMux I__1493 (
            .O(N__7180),
            .I(N__7155));
    InMux I__1492 (
            .O(N__7179),
            .I(N__7150));
    InMux I__1491 (
            .O(N__7178),
            .I(N__7150));
    InMux I__1490 (
            .O(N__7177),
            .I(N__7147));
    LocalMux I__1489 (
            .O(N__7174),
            .I(\U712_CHIP_RAM.N_276 ));
    Odrv4 I__1488 (
            .O(N__7171),
            .I(\U712_CHIP_RAM.N_276 ));
    LocalMux I__1487 (
            .O(N__7168),
            .I(\U712_CHIP_RAM.N_276 ));
    LocalMux I__1486 (
            .O(N__7165),
            .I(\U712_CHIP_RAM.N_276 ));
    Odrv4 I__1485 (
            .O(N__7160),
            .I(\U712_CHIP_RAM.N_276 ));
    LocalMux I__1484 (
            .O(N__7155),
            .I(\U712_CHIP_RAM.N_276 ));
    LocalMux I__1483 (
            .O(N__7150),
            .I(\U712_CHIP_RAM.N_276 ));
    LocalMux I__1482 (
            .O(N__7147),
            .I(\U712_CHIP_RAM.N_276 ));
    InMux I__1481 (
            .O(N__7130),
            .I(N__7118));
    InMux I__1480 (
            .O(N__7129),
            .I(N__7118));
    InMux I__1479 (
            .O(N__7128),
            .I(N__7118));
    InMux I__1478 (
            .O(N__7127),
            .I(N__7115));
    CascadeMux I__1477 (
            .O(N__7126),
            .I(N__7109));
    InMux I__1476 (
            .O(N__7125),
            .I(N__7105));
    LocalMux I__1475 (
            .O(N__7118),
            .I(N__7102));
    LocalMux I__1474 (
            .O(N__7115),
            .I(N__7099));
    InMux I__1473 (
            .O(N__7114),
            .I(N__7092));
    InMux I__1472 (
            .O(N__7113),
            .I(N__7092));
    InMux I__1471 (
            .O(N__7112),
            .I(N__7085));
    InMux I__1470 (
            .O(N__7109),
            .I(N__7085));
    InMux I__1469 (
            .O(N__7108),
            .I(N__7085));
    LocalMux I__1468 (
            .O(N__7105),
            .I(N__7078));
    Span4Mux_v I__1467 (
            .O(N__7102),
            .I(N__7078));
    Span4Mux_v I__1466 (
            .O(N__7099),
            .I(N__7078));
    InMux I__1465 (
            .O(N__7098),
            .I(N__7073));
    InMux I__1464 (
            .O(N__7097),
            .I(N__7073));
    LocalMux I__1463 (
            .O(N__7092),
            .I(N__7070));
    LocalMux I__1462 (
            .O(N__7085),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1461 (
            .O(N__7078),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1460 (
            .O(N__7073),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv12 I__1459 (
            .O(N__7070),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__1458 (
            .O(N__7061),
            .I(N__7057));
    InMux I__1457 (
            .O(N__7060),
            .I(N__7054));
    LocalMux I__1456 (
            .O(N__7057),
            .I(N__7051));
    LocalMux I__1455 (
            .O(N__7054),
            .I(N__7048));
    Span4Mux_h I__1454 (
            .O(N__7051),
            .I(N__7045));
    Span4Mux_h I__1453 (
            .O(N__7048),
            .I(N__7038));
    Span4Mux_v I__1452 (
            .O(N__7045),
            .I(N__7038));
    InMux I__1451 (
            .O(N__7044),
            .I(N__7035));
    InMux I__1450 (
            .O(N__7043),
            .I(N__7032));
    Odrv4 I__1449 (
            .O(N__7038),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1448 (
            .O(N__7035),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1447 (
            .O(N__7032),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1446 (
            .O(N__7025),
            .I(N__7022));
    LocalMux I__1445 (
            .O(N__7022),
            .I(N__7019));
    Span4Mux_s3_v I__1444 (
            .O(N__7019),
            .I(N__7016));
    Span4Mux_v I__1443 (
            .O(N__7016),
            .I(N__7013));
    Span4Mux_v I__1442 (
            .O(N__7013),
            .I(N__7010));
    Sp12to4 I__1441 (
            .O(N__7010),
            .I(N__7007));
    Odrv12 I__1440 (
            .O(N__7007),
            .I(CRCSn_c));
    InMux I__1439 (
            .O(N__7004),
            .I(N__7001));
    LocalMux I__1438 (
            .O(N__7001),
            .I(N__6997));
    InMux I__1437 (
            .O(N__7000),
            .I(N__6994));
    Odrv4 I__1436 (
            .O(N__6997),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_a2_0 ));
    LocalMux I__1435 (
            .O(N__6994),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_a2_0 ));
    CascadeMux I__1434 (
            .O(N__6989),
            .I(N__6986));
    InMux I__1433 (
            .O(N__6986),
            .I(N__6983));
    LocalMux I__1432 (
            .O(N__6983),
            .I(N__6980));
    Odrv4 I__1431 (
            .O(N__6980),
            .I(\U712_CHIP_RAM.N_314 ));
    InMux I__1430 (
            .O(N__6977),
            .I(N__6972));
    InMux I__1429 (
            .O(N__6976),
            .I(N__6969));
    InMux I__1428 (
            .O(N__6975),
            .I(N__6966));
    LocalMux I__1427 (
            .O(N__6972),
            .I(N__6959));
    LocalMux I__1426 (
            .O(N__6969),
            .I(N__6956));
    LocalMux I__1425 (
            .O(N__6966),
            .I(N__6951));
    InMux I__1424 (
            .O(N__6965),
            .I(N__6946));
    InMux I__1423 (
            .O(N__6964),
            .I(N__6946));
    InMux I__1422 (
            .O(N__6963),
            .I(N__6943));
    InMux I__1421 (
            .O(N__6962),
            .I(N__6940));
    Span4Mux_v I__1420 (
            .O(N__6959),
            .I(N__6935));
    Span4Mux_v I__1419 (
            .O(N__6956),
            .I(N__6935));
    InMux I__1418 (
            .O(N__6955),
            .I(N__6930));
    InMux I__1417 (
            .O(N__6954),
            .I(N__6930));
    Span4Mux_h I__1416 (
            .O(N__6951),
            .I(N__6925));
    LocalMux I__1415 (
            .O(N__6946),
            .I(N__6925));
    LocalMux I__1414 (
            .O(N__6943),
            .I(\U712_CHIP_RAM.N_293 ));
    LocalMux I__1413 (
            .O(N__6940),
            .I(\U712_CHIP_RAM.N_293 ));
    Odrv4 I__1412 (
            .O(N__6935),
            .I(\U712_CHIP_RAM.N_293 ));
    LocalMux I__1411 (
            .O(N__6930),
            .I(\U712_CHIP_RAM.N_293 ));
    Odrv4 I__1410 (
            .O(N__6925),
            .I(\U712_CHIP_RAM.N_293 ));
    InMux I__1409 (
            .O(N__6914),
            .I(N__6909));
    InMux I__1408 (
            .O(N__6913),
            .I(N__6906));
    InMux I__1407 (
            .O(N__6912),
            .I(N__6903));
    LocalMux I__1406 (
            .O(N__6909),
            .I(N__6898));
    LocalMux I__1405 (
            .O(N__6906),
            .I(N__6898));
    LocalMux I__1404 (
            .O(N__6903),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__1403 (
            .O(N__6898),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    InMux I__1402 (
            .O(N__6893),
            .I(N__6890));
    LocalMux I__1401 (
            .O(N__6890),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i ));
    CascadeMux I__1400 (
            .O(N__6887),
            .I(\U712_CHIP_RAM.REFRESH_RNO_0Z0Z_0_cascade_ ));
    InMux I__1399 (
            .O(N__6884),
            .I(N__6881));
    LocalMux I__1398 (
            .O(N__6881),
            .I(\U712_CHIP_RAM.REFRESHZ0Z_0 ));
    CascadeMux I__1397 (
            .O(N__6878),
            .I(\U712_CHIP_RAM.REFRESH9lt7_cascade_ ));
    InMux I__1396 (
            .O(N__6875),
            .I(N__6872));
    LocalMux I__1395 (
            .O(N__6872),
            .I(N__6869));
    Odrv4 I__1394 (
            .O(N__6869),
            .I(\U712_CHIP_RAM.REFRESHZ0Z_1 ));
    InMux I__1393 (
            .O(N__6866),
            .I(N__6860));
    InMux I__1392 (
            .O(N__6865),
            .I(N__6860));
    LocalMux I__1391 (
            .O(N__6860),
            .I(\U712_CHIP_RAM.REFRESH9lto7_0 ));
    InMux I__1390 (
            .O(N__6857),
            .I(N__6854));
    LocalMux I__1389 (
            .O(N__6854),
            .I(N__6851));
    Span4Mux_v I__1388 (
            .O(N__6851),
            .I(N__6848));
    Sp12to4 I__1387 (
            .O(N__6848),
            .I(N__6845));
    Span12Mux_h I__1386 (
            .O(N__6845),
            .I(N__6842));
    Odrv12 I__1385 (
            .O(N__6842),
            .I(A_c_14));
    CascadeMux I__1384 (
            .O(N__6839),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5_cascade_ ));
    InMux I__1383 (
            .O(N__6836),
            .I(N__6833));
    LocalMux I__1382 (
            .O(N__6833),
            .I(N__6830));
    Sp12to4 I__1381 (
            .O(N__6830),
            .I(N__6827));
    Span12Mux_v I__1380 (
            .O(N__6827),
            .I(N__6824));
    Span12Mux_h I__1379 (
            .O(N__6824),
            .I(N__6821));
    Odrv12 I__1378 (
            .O(N__6821),
            .I(A_c_7));
    InMux I__1377 (
            .O(N__6818),
            .I(N__6815));
    LocalMux I__1376 (
            .O(N__6815),
            .I(N__6812));
    Odrv12 I__1375 (
            .O(N__6812),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__1374 (
            .O(N__6809),
            .I(N__6806));
    LocalMux I__1373 (
            .O(N__6806),
            .I(N__6803));
    Span4Mux_v I__1372 (
            .O(N__6803),
            .I(N__6800));
    Span4Mux_h I__1371 (
            .O(N__6800),
            .I(N__6797));
    Sp12to4 I__1370 (
            .O(N__6797),
            .I(N__6794));
    Odrv12 I__1369 (
            .O(N__6794),
            .I(A_c_15));
    CascadeMux I__1368 (
            .O(N__6791),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6_cascade_ ));
    InMux I__1367 (
            .O(N__6788),
            .I(N__6785));
    LocalMux I__1366 (
            .O(N__6785),
            .I(N__6782));
    Span4Mux_v I__1365 (
            .O(N__6782),
            .I(N__6779));
    Span4Mux_v I__1364 (
            .O(N__6779),
            .I(N__6776));
    Sp12to4 I__1363 (
            .O(N__6776),
            .I(N__6773));
    Span12Mux_h I__1362 (
            .O(N__6773),
            .I(N__6770));
    Odrv12 I__1361 (
            .O(N__6770),
            .I(A_c_8));
    InMux I__1360 (
            .O(N__6767),
            .I(N__6764));
    LocalMux I__1359 (
            .O(N__6764),
            .I(N__6761));
    Span4Mux_v I__1358 (
            .O(N__6761),
            .I(N__6758));
    Span4Mux_v I__1357 (
            .O(N__6758),
            .I(N__6755));
    Sp12to4 I__1356 (
            .O(N__6755),
            .I(N__6752));
    Span12Mux_h I__1355 (
            .O(N__6752),
            .I(N__6749));
    Odrv12 I__1354 (
            .O(N__6749),
            .I(A_c_9));
    InMux I__1353 (
            .O(N__6746),
            .I(N__6743));
    LocalMux I__1352 (
            .O(N__6743),
            .I(N__6740));
    Span4Mux_v I__1351 (
            .O(N__6740),
            .I(N__6737));
    Sp12to4 I__1350 (
            .O(N__6737),
            .I(N__6734));
    Span12Mux_v I__1349 (
            .O(N__6734),
            .I(N__6731));
    Span12Mux_h I__1348 (
            .O(N__6731),
            .I(N__6728));
    Odrv12 I__1347 (
            .O(N__6728),
            .I(A_c_2));
    CascadeMux I__1346 (
            .O(N__6725),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0_cascade_ ));
    CascadeMux I__1345 (
            .O(N__6722),
            .I(\U712_CHIP_RAM.N_315_cascade_ ));
    IoInMux I__1344 (
            .O(N__6719),
            .I(N__6716));
    LocalMux I__1343 (
            .O(N__6716),
            .I(N__6713));
    Span4Mux_s0_v I__1342 (
            .O(N__6713),
            .I(N__6710));
    Sp12to4 I__1341 (
            .O(N__6710),
            .I(N__6707));
    Span12Mux_h I__1340 (
            .O(N__6707),
            .I(N__6704));
    Odrv12 I__1339 (
            .O(N__6704),
            .I(CMA_c_0));
    InMux I__1338 (
            .O(N__6701),
            .I(N__6698));
    LocalMux I__1337 (
            .O(N__6698),
            .I(N__6695));
    Span4Mux_v I__1336 (
            .O(N__6695),
            .I(N__6692));
    Sp12to4 I__1335 (
            .O(N__6692),
            .I(N__6689));
    Span12Mux_h I__1334 (
            .O(N__6689),
            .I(N__6686));
    Span12Mux_v I__1333 (
            .O(N__6686),
            .I(N__6683));
    Odrv12 I__1332 (
            .O(N__6683),
            .I(A_c_3));
    InMux I__1331 (
            .O(N__6680),
            .I(N__6677));
    LocalMux I__1330 (
            .O(N__6677),
            .I(N__6674));
    Span4Mux_v I__1329 (
            .O(N__6674),
            .I(N__6671));
    Span4Mux_h I__1328 (
            .O(N__6671),
            .I(N__6668));
    Sp12to4 I__1327 (
            .O(N__6668),
            .I(N__6665));
    Odrv12 I__1326 (
            .O(N__6665),
            .I(A_c_10));
    CascadeMux I__1325 (
            .O(N__6662),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_ ));
    CascadeMux I__1324 (
            .O(N__6659),
            .I(N__6656));
    InMux I__1323 (
            .O(N__6656),
            .I(N__6653));
    LocalMux I__1322 (
            .O(N__6653),
            .I(N__6650));
    Odrv4 I__1321 (
            .O(N__6650),
            .I(\U712_CHIP_RAM.N_316 ));
    CascadeMux I__1320 (
            .O(N__6647),
            .I(N__6641));
    InMux I__1319 (
            .O(N__6646),
            .I(N__6635));
    InMux I__1318 (
            .O(N__6645),
            .I(N__6632));
    InMux I__1317 (
            .O(N__6644),
            .I(N__6629));
    InMux I__1316 (
            .O(N__6641),
            .I(N__6626));
    InMux I__1315 (
            .O(N__6640),
            .I(N__6619));
    InMux I__1314 (
            .O(N__6639),
            .I(N__6619));
    InMux I__1313 (
            .O(N__6638),
            .I(N__6619));
    LocalMux I__1312 (
            .O(N__6635),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__1311 (
            .O(N__6632),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__1310 (
            .O(N__6629),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__1309 (
            .O(N__6626),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__1308 (
            .O(N__6619),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__1307 (
            .O(N__6608),
            .I(N__6600));
    InMux I__1306 (
            .O(N__6607),
            .I(N__6597));
    InMux I__1305 (
            .O(N__6606),
            .I(N__6590));
    InMux I__1304 (
            .O(N__6605),
            .I(N__6590));
    InMux I__1303 (
            .O(N__6604),
            .I(N__6590));
    InMux I__1302 (
            .O(N__6603),
            .I(N__6587));
    LocalMux I__1301 (
            .O(N__6600),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1300 (
            .O(N__6597),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1299 (
            .O(N__6590),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1298 (
            .O(N__6587),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    InMux I__1297 (
            .O(N__6578),
            .I(N__6571));
    InMux I__1296 (
            .O(N__6577),
            .I(N__6568));
    InMux I__1295 (
            .O(N__6576),
            .I(N__6561));
    InMux I__1294 (
            .O(N__6575),
            .I(N__6561));
    InMux I__1293 (
            .O(N__6574),
            .I(N__6561));
    LocalMux I__1292 (
            .O(N__6571),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__1291 (
            .O(N__6568),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__1290 (
            .O(N__6561),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    InMux I__1289 (
            .O(N__6554),
            .I(N__6548));
    InMux I__1288 (
            .O(N__6553),
            .I(N__6543));
    InMux I__1287 (
            .O(N__6552),
            .I(N__6543));
    InMux I__1286 (
            .O(N__6551),
            .I(N__6540));
    LocalMux I__1285 (
            .O(N__6548),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__1284 (
            .O(N__6543),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__1283 (
            .O(N__6540),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__1282 (
            .O(N__6533),
            .I(N__6527));
    InMux I__1281 (
            .O(N__6532),
            .I(N__6524));
    CascadeMux I__1280 (
            .O(N__6531),
            .I(N__6520));
    InMux I__1279 (
            .O(N__6530),
            .I(N__6516));
    LocalMux I__1278 (
            .O(N__6527),
            .I(N__6511));
    LocalMux I__1277 (
            .O(N__6524),
            .I(N__6511));
    InMux I__1276 (
            .O(N__6523),
            .I(N__6504));
    InMux I__1275 (
            .O(N__6520),
            .I(N__6504));
    InMux I__1274 (
            .O(N__6519),
            .I(N__6504));
    LocalMux I__1273 (
            .O(N__6516),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1272 (
            .O(N__6511),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1271 (
            .O(N__6504),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    IoInMux I__1270 (
            .O(N__6497),
            .I(N__6494));
    LocalMux I__1269 (
            .O(N__6494),
            .I(N__6491));
    Odrv12 I__1268 (
            .O(N__6491),
            .I(CMA_c_2));
    IoInMux I__1267 (
            .O(N__6488),
            .I(N__6485));
    LocalMux I__1266 (
            .O(N__6485),
            .I(N__6482));
    Span4Mux_s3_v I__1265 (
            .O(N__6482),
            .I(N__6479));
    Odrv4 I__1264 (
            .O(N__6479),
            .I(CMA_c_1));
    IoInMux I__1263 (
            .O(N__6476),
            .I(N__6473));
    LocalMux I__1262 (
            .O(N__6473),
            .I(N__6470));
    Span4Mux_s3_v I__1261 (
            .O(N__6470),
            .I(N__6467));
    Span4Mux_h I__1260 (
            .O(N__6467),
            .I(N__6464));
    Span4Mux_h I__1259 (
            .O(N__6464),
            .I(N__6461));
    Odrv4 I__1258 (
            .O(N__6461),
            .I(CMA_c_10));
    InMux I__1257 (
            .O(N__6458),
            .I(N__6455));
    LocalMux I__1256 (
            .O(N__6455),
            .I(N__6452));
    Span4Mux_v I__1255 (
            .O(N__6452),
            .I(N__6449));
    Span4Mux_h I__1254 (
            .O(N__6449),
            .I(N__6446));
    Sp12to4 I__1253 (
            .O(N__6446),
            .I(N__6443));
    Odrv12 I__1252 (
            .O(N__6443),
            .I(A_c_11));
    CascadeMux I__1251 (
            .O(N__6440),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_ ));
    InMux I__1250 (
            .O(N__6437),
            .I(N__6434));
    LocalMux I__1249 (
            .O(N__6434),
            .I(N__6431));
    Span4Mux_v I__1248 (
            .O(N__6431),
            .I(N__6428));
    Sp12to4 I__1247 (
            .O(N__6428),
            .I(N__6425));
    Span12Mux_h I__1246 (
            .O(N__6425),
            .I(N__6422));
    Span12Mux_v I__1245 (
            .O(N__6422),
            .I(N__6419));
    Odrv12 I__1244 (
            .O(N__6419),
            .I(A_c_4));
    InMux I__1243 (
            .O(N__6416),
            .I(N__6413));
    LocalMux I__1242 (
            .O(N__6413),
            .I(\U712_CHIP_RAM.N_317 ));
    CascadeMux I__1241 (
            .O(N__6410),
            .I(N__6407));
    InMux I__1240 (
            .O(N__6407),
            .I(N__6402));
    InMux I__1239 (
            .O(N__6406),
            .I(N__6399));
    InMux I__1238 (
            .O(N__6405),
            .I(N__6396));
    LocalMux I__1237 (
            .O(N__6402),
            .I(\U712_REG_SM.N_292 ));
    LocalMux I__1236 (
            .O(N__6399),
            .I(\U712_REG_SM.N_292 ));
    LocalMux I__1235 (
            .O(N__6396),
            .I(\U712_REG_SM.N_292 ));
    InMux I__1234 (
            .O(N__6389),
            .I(N__6384));
    InMux I__1233 (
            .O(N__6388),
            .I(N__6379));
    InMux I__1232 (
            .O(N__6387),
            .I(N__6379));
    LocalMux I__1231 (
            .O(N__6384),
            .I(\U712_REG_SM.N_298 ));
    LocalMux I__1230 (
            .O(N__6379),
            .I(\U712_REG_SM.N_298 ));
    CascadeMux I__1229 (
            .O(N__6374),
            .I(N__6368));
    InMux I__1228 (
            .O(N__6373),
            .I(N__6365));
    InMux I__1227 (
            .O(N__6372),
            .I(N__6362));
    InMux I__1226 (
            .O(N__6371),
            .I(N__6357));
    InMux I__1225 (
            .O(N__6368),
            .I(N__6357));
    LocalMux I__1224 (
            .O(N__6365),
            .I(\U712_REG_SM.N_294 ));
    LocalMux I__1223 (
            .O(N__6362),
            .I(\U712_REG_SM.N_294 ));
    LocalMux I__1222 (
            .O(N__6357),
            .I(\U712_REG_SM.N_294 ));
    InMux I__1221 (
            .O(N__6350),
            .I(N__6344));
    InMux I__1220 (
            .O(N__6349),
            .I(N__6344));
    LocalMux I__1219 (
            .O(N__6344),
            .I(\U712_REG_SM.N_309 ));
    CascadeMux I__1218 (
            .O(N__6341),
            .I(N__6338));
    InMux I__1217 (
            .O(N__6338),
            .I(N__6334));
    InMux I__1216 (
            .O(N__6337),
            .I(N__6331));
    LocalMux I__1215 (
            .O(N__6334),
            .I(\U712_REG_SM.N_282 ));
    LocalMux I__1214 (
            .O(N__6331),
            .I(\U712_REG_SM.N_282 ));
    CascadeMux I__1213 (
            .O(N__6326),
            .I(\U712_REG_SM.N_282_cascade_ ));
    CascadeMux I__1212 (
            .O(N__6323),
            .I(N__6319));
    InMux I__1211 (
            .O(N__6322),
            .I(N__6316));
    InMux I__1210 (
            .O(N__6319),
            .I(N__6313));
    LocalMux I__1209 (
            .O(N__6316),
            .I(N__6310));
    LocalMux I__1208 (
            .O(N__6313),
            .I(\U712_REG_SM.N_306 ));
    Odrv4 I__1207 (
            .O(N__6310),
            .I(\U712_REG_SM.N_306 ));
    CascadeMux I__1206 (
            .O(N__6305),
            .I(N__6301));
    InMux I__1205 (
            .O(N__6304),
            .I(N__6295));
    InMux I__1204 (
            .O(N__6301),
            .I(N__6295));
    InMux I__1203 (
            .O(N__6300),
            .I(N__6292));
    LocalMux I__1202 (
            .O(N__6295),
            .I(N__6287));
    LocalMux I__1201 (
            .O(N__6292),
            .I(N__6287));
    Span12Mux_v I__1200 (
            .O(N__6287),
            .I(N__6284));
    Span12Mux_h I__1199 (
            .O(N__6284),
            .I(N__6281));
    Span12Mux_v I__1198 (
            .O(N__6281),
            .I(N__6278));
    Odrv12 I__1197 (
            .O(N__6278),
            .I(SIZ_c_1));
    InMux I__1196 (
            .O(N__6275),
            .I(N__6272));
    LocalMux I__1195 (
            .O(N__6272),
            .I(N__6269));
    Odrv4 I__1194 (
            .O(N__6269),
            .I(\U712_BYTE_ENABLE.N_407 ));
    InMux I__1193 (
            .O(N__6266),
            .I(N__6258));
    InMux I__1192 (
            .O(N__6265),
            .I(N__6258));
    InMux I__1191 (
            .O(N__6264),
            .I(N__6253));
    InMux I__1190 (
            .O(N__6263),
            .I(N__6253));
    LocalMux I__1189 (
            .O(N__6258),
            .I(N__6248));
    LocalMux I__1188 (
            .O(N__6253),
            .I(N__6248));
    Span4Mux_v I__1187 (
            .O(N__6248),
            .I(N__6245));
    Sp12to4 I__1186 (
            .O(N__6245),
            .I(N__6242));
    Span12Mux_h I__1185 (
            .O(N__6242),
            .I(N__6239));
    Span12Mux_v I__1184 (
            .O(N__6239),
            .I(N__6236));
    Odrv12 I__1183 (
            .O(N__6236),
            .I(A_c_1));
    InMux I__1182 (
            .O(N__6233),
            .I(N__6225));
    InMux I__1181 (
            .O(N__6232),
            .I(N__6225));
    InMux I__1180 (
            .O(N__6231),
            .I(N__6222));
    InMux I__1179 (
            .O(N__6230),
            .I(N__6219));
    LocalMux I__1178 (
            .O(N__6225),
            .I(N__6214));
    LocalMux I__1177 (
            .O(N__6222),
            .I(N__6214));
    LocalMux I__1176 (
            .O(N__6219),
            .I(N__6211));
    Span4Mux_v I__1175 (
            .O(N__6214),
            .I(N__6208));
    Span4Mux_v I__1174 (
            .O(N__6211),
            .I(N__6205));
    Span4Mux_v I__1173 (
            .O(N__6208),
            .I(N__6198));
    Span4Mux_v I__1172 (
            .O(N__6205),
            .I(N__6198));
    InMux I__1171 (
            .O(N__6204),
            .I(N__6193));
    InMux I__1170 (
            .O(N__6203),
            .I(N__6193));
    Span4Mux_h I__1169 (
            .O(N__6198),
            .I(N__6190));
    LocalMux I__1168 (
            .O(N__6193),
            .I(N__6187));
    Sp12to4 I__1167 (
            .O(N__6190),
            .I(N__6182));
    Span12Mux_v I__1166 (
            .O(N__6187),
            .I(N__6182));
    Odrv12 I__1165 (
            .O(N__6182),
            .I(A_c_0));
    InMux I__1164 (
            .O(N__6179),
            .I(N__6176));
    LocalMux I__1163 (
            .O(N__6176),
            .I(\U712_BYTE_ENABLE.N_409 ));
    InMux I__1162 (
            .O(N__6173),
            .I(N__6170));
    LocalMux I__1161 (
            .O(N__6170),
            .I(N__6166));
    IoInMux I__1160 (
            .O(N__6169),
            .I(N__6163));
    Span4Mux_v I__1159 (
            .O(N__6166),
            .I(N__6160));
    LocalMux I__1158 (
            .O(N__6163),
            .I(N__6157));
    Sp12to4 I__1157 (
            .O(N__6160),
            .I(N__6154));
    Span4Mux_s3_h I__1156 (
            .O(N__6157),
            .I(N__6151));
    Span12Mux_h I__1155 (
            .O(N__6154),
            .I(N__6146));
    Sp12to4 I__1154 (
            .O(N__6151),
            .I(N__6146));
    Span12Mux_v I__1153 (
            .O(N__6146),
            .I(N__6143));
    Odrv12 I__1152 (
            .O(N__6143),
            .I(C1_c));
    InMux I__1151 (
            .O(N__6140),
            .I(N__6137));
    LocalMux I__1150 (
            .O(N__6137),
            .I(N__6134));
    Span12Mux_h I__1149 (
            .O(N__6134),
            .I(N__6131));
    Span12Mux_v I__1148 (
            .O(N__6131),
            .I(N__6128));
    Odrv12 I__1147 (
            .O(N__6128),
            .I(C3_c));
    InMux I__1146 (
            .O(N__6125),
            .I(N__6121));
    InMux I__1145 (
            .O(N__6124),
            .I(N__6118));
    LocalMux I__1144 (
            .O(N__6121),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    LocalMux I__1143 (
            .O(N__6118),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    CascadeMux I__1142 (
            .O(N__6113),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0_cascade_ ));
    IoInMux I__1141 (
            .O(N__6110),
            .I(N__6107));
    LocalMux I__1140 (
            .O(N__6107),
            .I(N__6104));
    Span4Mux_s3_h I__1139 (
            .O(N__6104),
            .I(N__6101));
    Span4Mux_v I__1138 (
            .O(N__6101),
            .I(N__6098));
    Sp12to4 I__1137 (
            .O(N__6098),
            .I(N__6095));
    Span12Mux_h I__1136 (
            .O(N__6095),
            .I(N__6092));
    Odrv12 I__1135 (
            .O(N__6092),
            .I(N_192_i));
    InMux I__1134 (
            .O(N__6089),
            .I(N__6086));
    LocalMux I__1133 (
            .O(N__6086),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0 ));
    IoInMux I__1132 (
            .O(N__6083),
            .I(N__6080));
    LocalMux I__1131 (
            .O(N__6080),
            .I(N__6077));
    Span12Mux_s6_h I__1130 (
            .O(N__6077),
            .I(N__6074));
    Span12Mux_h I__1129 (
            .O(N__6074),
            .I(N__6071));
    Span12Mux_v I__1128 (
            .O(N__6071),
            .I(N__6068));
    Odrv12 I__1127 (
            .O(N__6068),
            .I(N_194_i));
    InMux I__1126 (
            .O(N__6065),
            .I(N__6062));
    LocalMux I__1125 (
            .O(N__6062),
            .I(N__6059));
    Span4Mux_v I__1124 (
            .O(N__6059),
            .I(N__6055));
    InMux I__1123 (
            .O(N__6058),
            .I(N__6052));
    Sp12to4 I__1122 (
            .O(N__6055),
            .I(N__6047));
    LocalMux I__1121 (
            .O(N__6052),
            .I(N__6047));
    Span12Mux_h I__1120 (
            .O(N__6047),
            .I(N__6044));
    Span12Mux_v I__1119 (
            .O(N__6044),
            .I(N__6041));
    Odrv12 I__1118 (
            .O(N__6041),
            .I(SIZ_c_0));
    IoInMux I__1117 (
            .O(N__6038),
            .I(N__6035));
    LocalMux I__1116 (
            .O(N__6035),
            .I(N__6032));
    Span4Mux_s3_v I__1115 (
            .O(N__6032),
            .I(N__6029));
    Span4Mux_v I__1114 (
            .O(N__6029),
            .I(N__6026));
    Span4Mux_v I__1113 (
            .O(N__6026),
            .I(N__6021));
    InMux I__1112 (
            .O(N__6025),
            .I(N__6018));
    InMux I__1111 (
            .O(N__6024),
            .I(N__6015));
    Span4Mux_h I__1110 (
            .O(N__6021),
            .I(N__6011));
    LocalMux I__1109 (
            .O(N__6018),
            .I(N__6006));
    LocalMux I__1108 (
            .O(N__6015),
            .I(N__6006));
    InMux I__1107 (
            .O(N__6014),
            .I(N__6003));
    Odrv4 I__1106 (
            .O(N__6011),
            .I(DBENn_c));
    Odrv4 I__1105 (
            .O(N__6006),
            .I(DBENn_c));
    LocalMux I__1104 (
            .O(N__6003),
            .I(DBENn_c));
    IoInMux I__1103 (
            .O(N__5996),
            .I(N__5993));
    LocalMux I__1102 (
            .O(N__5993),
            .I(N__5990));
    Span4Mux_s2_v I__1101 (
            .O(N__5990),
            .I(N__5987));
    Span4Mux_h I__1100 (
            .O(N__5987),
            .I(N__5984));
    Span4Mux_h I__1099 (
            .O(N__5984),
            .I(N__5979));
    InMux I__1098 (
            .O(N__5983),
            .I(N__5974));
    InMux I__1097 (
            .O(N__5982),
            .I(N__5974));
    Sp12to4 I__1096 (
            .O(N__5979),
            .I(N__5969));
    LocalMux I__1095 (
            .O(N__5974),
            .I(N__5966));
    InMux I__1094 (
            .O(N__5973),
            .I(N__5963));
    InMux I__1093 (
            .O(N__5972),
            .I(N__5960));
    Span12Mux_s9_v I__1092 (
            .O(N__5969),
            .I(N__5948));
    Sp12to4 I__1091 (
            .O(N__5966),
            .I(N__5948));
    LocalMux I__1090 (
            .O(N__5963),
            .I(N__5948));
    LocalMux I__1089 (
            .O(N__5960),
            .I(N__5948));
    InMux I__1088 (
            .O(N__5959),
            .I(N__5941));
    InMux I__1087 (
            .O(N__5958),
            .I(N__5941));
    InMux I__1086 (
            .O(N__5957),
            .I(N__5941));
    Odrv12 I__1085 (
            .O(N__5948),
            .I(RAMENn_c));
    LocalMux I__1084 (
            .O(N__5941),
            .I(RAMENn_c));
    CascadeMux I__1083 (
            .O(N__5936),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_cascade_ ));
    IoInMux I__1082 (
            .O(N__5933),
            .I(N__5930));
    LocalMux I__1081 (
            .O(N__5930),
            .I(N__5927));
    Span12Mux_s6_h I__1080 (
            .O(N__5927),
            .I(N__5924));
    Span12Mux_h I__1079 (
            .O(N__5924),
            .I(N__5921));
    Span12Mux_v I__1078 (
            .O(N__5921),
            .I(N__5918));
    Odrv12 I__1077 (
            .O(N__5918),
            .I(N_196_i));
    InMux I__1076 (
            .O(N__5915),
            .I(N__5907));
    InMux I__1075 (
            .O(N__5914),
            .I(N__5907));
    InMux I__1074 (
            .O(N__5913),
            .I(N__5902));
    InMux I__1073 (
            .O(N__5912),
            .I(N__5902));
    LocalMux I__1072 (
            .O(N__5907),
            .I(\U712_BYTE_ENABLE.N_404 ));
    LocalMux I__1071 (
            .O(N__5902),
            .I(\U712_BYTE_ENABLE.N_404 ));
    InMux I__1070 (
            .O(N__5897),
            .I(N__5894));
    LocalMux I__1069 (
            .O(N__5894),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0 ));
    CascadeMux I__1068 (
            .O(N__5891),
            .I(\U712_BYTE_ENABLE.N_411_cascade_ ));
    IoInMux I__1067 (
            .O(N__5888),
            .I(N__5885));
    LocalMux I__1066 (
            .O(N__5885),
            .I(N__5882));
    IoSpan4Mux I__1065 (
            .O(N__5882),
            .I(N__5879));
    Sp12to4 I__1064 (
            .O(N__5879),
            .I(N__5876));
    Span12Mux_s7_v I__1063 (
            .O(N__5876),
            .I(N__5873));
    Odrv12 I__1062 (
            .O(N__5873),
            .I(N_198_i));
    InMux I__1061 (
            .O(N__5870),
            .I(N__5867));
    LocalMux I__1060 (
            .O(N__5867),
            .I(\U712_BYTE_ENABLE.N_405 ));
    CascadeMux I__1059 (
            .O(N__5864),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_cascade_ ));
    InMux I__1058 (
            .O(N__5861),
            .I(N__5858));
    LocalMux I__1057 (
            .O(N__5858),
            .I(\U712_CHIP_RAM.DBENn_7_0_a2_0 ));
    CascadeMux I__1056 (
            .O(N__5855),
            .I(N__5852));
    InMux I__1055 (
            .O(N__5852),
            .I(N__5847));
    InMux I__1054 (
            .O(N__5851),
            .I(N__5844));
    InMux I__1053 (
            .O(N__5850),
            .I(N__5841));
    LocalMux I__1052 (
            .O(N__5847),
            .I(N__5838));
    LocalMux I__1051 (
            .O(N__5844),
            .I(N__5835));
    LocalMux I__1050 (
            .O(N__5841),
            .I(\U712_CHIP_RAM.N_347 ));
    Odrv4 I__1049 (
            .O(N__5838),
            .I(\U712_CHIP_RAM.N_347 ));
    Odrv4 I__1048 (
            .O(N__5835),
            .I(\U712_CHIP_RAM.N_347 ));
    InMux I__1047 (
            .O(N__5828),
            .I(N__5825));
    LocalMux I__1046 (
            .O(N__5825),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_3_1 ));
    CascadeMux I__1045 (
            .O(N__5822),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_2_1_cascade_ ));
    InMux I__1044 (
            .O(N__5819),
            .I(N__5814));
    InMux I__1043 (
            .O(N__5818),
            .I(N__5811));
    InMux I__1042 (
            .O(N__5817),
            .I(N__5808));
    LocalMux I__1041 (
            .O(N__5814),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER50 ));
    LocalMux I__1040 (
            .O(N__5811),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER50 ));
    LocalMux I__1039 (
            .O(N__5808),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER50 ));
    InMux I__1038 (
            .O(N__5801),
            .I(N__5795));
    InMux I__1037 (
            .O(N__5800),
            .I(N__5784));
    CascadeMux I__1036 (
            .O(N__5799),
            .I(N__5778));
    InMux I__1035 (
            .O(N__5798),
            .I(N__5775));
    LocalMux I__1034 (
            .O(N__5795),
            .I(N__5772));
    InMux I__1033 (
            .O(N__5794),
            .I(N__5765));
    InMux I__1032 (
            .O(N__5793),
            .I(N__5765));
    InMux I__1031 (
            .O(N__5792),
            .I(N__5765));
    InMux I__1030 (
            .O(N__5791),
            .I(N__5758));
    InMux I__1029 (
            .O(N__5790),
            .I(N__5758));
    InMux I__1028 (
            .O(N__5789),
            .I(N__5758));
    InMux I__1027 (
            .O(N__5788),
            .I(N__5753));
    InMux I__1026 (
            .O(N__5787),
            .I(N__5753));
    LocalMux I__1025 (
            .O(N__5784),
            .I(N__5750));
    CascadeMux I__1024 (
            .O(N__5783),
            .I(N__5747));
    CascadeMux I__1023 (
            .O(N__5782),
            .I(N__5743));
    CascadeMux I__1022 (
            .O(N__5781),
            .I(N__5738));
    InMux I__1021 (
            .O(N__5778),
            .I(N__5728));
    LocalMux I__1020 (
            .O(N__5775),
            .I(N__5723));
    Span4Mux_v I__1019 (
            .O(N__5772),
            .I(N__5723));
    LocalMux I__1018 (
            .O(N__5765),
            .I(N__5720));
    LocalMux I__1017 (
            .O(N__5758),
            .I(N__5713));
    LocalMux I__1016 (
            .O(N__5753),
            .I(N__5713));
    Span4Mux_h I__1015 (
            .O(N__5750),
            .I(N__5713));
    InMux I__1014 (
            .O(N__5747),
            .I(N__5706));
    InMux I__1013 (
            .O(N__5746),
            .I(N__5706));
    InMux I__1012 (
            .O(N__5743),
            .I(N__5706));
    InMux I__1011 (
            .O(N__5742),
            .I(N__5701));
    InMux I__1010 (
            .O(N__5741),
            .I(N__5701));
    InMux I__1009 (
            .O(N__5738),
            .I(N__5696));
    InMux I__1008 (
            .O(N__5737),
            .I(N__5696));
    InMux I__1007 (
            .O(N__5736),
            .I(N__5693));
    InMux I__1006 (
            .O(N__5735),
            .I(N__5686));
    InMux I__1005 (
            .O(N__5734),
            .I(N__5686));
    InMux I__1004 (
            .O(N__5733),
            .I(N__5686));
    InMux I__1003 (
            .O(N__5732),
            .I(N__5681));
    InMux I__1002 (
            .O(N__5731),
            .I(N__5681));
    LocalMux I__1001 (
            .O(N__5728),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1000 (
            .O(N__5723),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv12 I__999 (
            .O(N__5720),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__998 (
            .O(N__5713),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__997 (
            .O(N__5706),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__996 (
            .O(N__5701),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__995 (
            .O(N__5696),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__994 (
            .O(N__5693),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__993 (
            .O(N__5686),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__992 (
            .O(N__5681),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__991 (
            .O(N__5660),
            .I(N__5653));
    CascadeMux I__990 (
            .O(N__5659),
            .I(N__5650));
    CascadeMux I__989 (
            .O(N__5658),
            .I(N__5647));
    CascadeMux I__988 (
            .O(N__5657),
            .I(N__5643));
    InMux I__987 (
            .O(N__5656),
            .I(N__5639));
    LocalMux I__986 (
            .O(N__5653),
            .I(N__5634));
    InMux I__985 (
            .O(N__5650),
            .I(N__5629));
    InMux I__984 (
            .O(N__5647),
            .I(N__5629));
    InMux I__983 (
            .O(N__5646),
            .I(N__5626));
    InMux I__982 (
            .O(N__5643),
            .I(N__5623));
    InMux I__981 (
            .O(N__5642),
            .I(N__5620));
    LocalMux I__980 (
            .O(N__5639),
            .I(N__5617));
    CascadeMux I__979 (
            .O(N__5638),
            .I(N__5608));
    InMux I__978 (
            .O(N__5637),
            .I(N__5602));
    Span4Mux_v I__977 (
            .O(N__5634),
            .I(N__5597));
    LocalMux I__976 (
            .O(N__5629),
            .I(N__5597));
    LocalMux I__975 (
            .O(N__5626),
            .I(N__5592));
    LocalMux I__974 (
            .O(N__5623),
            .I(N__5592));
    LocalMux I__973 (
            .O(N__5620),
            .I(N__5587));
    Span4Mux_v I__972 (
            .O(N__5617),
            .I(N__5587));
    InMux I__971 (
            .O(N__5616),
            .I(N__5582));
    InMux I__970 (
            .O(N__5615),
            .I(N__5582));
    InMux I__969 (
            .O(N__5614),
            .I(N__5579));
    InMux I__968 (
            .O(N__5613),
            .I(N__5572));
    InMux I__967 (
            .O(N__5612),
            .I(N__5572));
    InMux I__966 (
            .O(N__5611),
            .I(N__5572));
    InMux I__965 (
            .O(N__5608),
            .I(N__5567));
    InMux I__964 (
            .O(N__5607),
            .I(N__5567));
    InMux I__963 (
            .O(N__5606),
            .I(N__5562));
    InMux I__962 (
            .O(N__5605),
            .I(N__5562));
    LocalMux I__961 (
            .O(N__5602),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__960 (
            .O(N__5597),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__959 (
            .O(N__5592),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__958 (
            .O(N__5587),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__957 (
            .O(N__5582),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__956 (
            .O(N__5579),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__955 (
            .O(N__5572),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__954 (
            .O(N__5567),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__953 (
            .O(N__5562),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__952 (
            .O(N__5543),
            .I(N__5536));
    InMux I__951 (
            .O(N__5542),
            .I(N__5536));
    CascadeMux I__950 (
            .O(N__5541),
            .I(N__5532));
    LocalMux I__949 (
            .O(N__5536),
            .I(N__5528));
    InMux I__948 (
            .O(N__5535),
            .I(N__5525));
    InMux I__947 (
            .O(N__5532),
            .I(N__5520));
    InMux I__946 (
            .O(N__5531),
            .I(N__5520));
    Odrv4 I__945 (
            .O(N__5528),
            .I(\U712_CHIP_RAM.N_273 ));
    LocalMux I__944 (
            .O(N__5525),
            .I(\U712_CHIP_RAM.N_273 ));
    LocalMux I__943 (
            .O(N__5520),
            .I(\U712_CHIP_RAM.N_273 ));
    CascadeMux I__942 (
            .O(N__5513),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_1_0_cascade_ ));
    InMux I__941 (
            .O(N__5510),
            .I(N__5506));
    InMux I__940 (
            .O(N__5509),
            .I(N__5503));
    LocalMux I__939 (
            .O(N__5506),
            .I(\U712_CHIP_RAM.N_305 ));
    LocalMux I__938 (
            .O(N__5503),
            .I(\U712_CHIP_RAM.N_305 ));
    CascadeMux I__937 (
            .O(N__5498),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_0_cascade_ ));
    InMux I__936 (
            .O(N__5495),
            .I(N__5487));
    InMux I__935 (
            .O(N__5494),
            .I(N__5487));
    InMux I__934 (
            .O(N__5493),
            .I(N__5482));
    InMux I__933 (
            .O(N__5492),
            .I(N__5482));
    LocalMux I__932 (
            .O(N__5487),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ));
    LocalMux I__931 (
            .O(N__5482),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ));
    CascadeMux I__930 (
            .O(N__5477),
            .I(\U712_CHIP_RAM.REFRESH_RST_cascade_ ));
    InMux I__929 (
            .O(N__5474),
            .I(N__5471));
    LocalMux I__928 (
            .O(N__5471),
            .I(\U712_CHIP_RAM.N_289 ));
    CascadeMux I__927 (
            .O(N__5468),
            .I(\U712_CHIP_RAM.N_425_cascade_ ));
    InMux I__926 (
            .O(N__5465),
            .I(N__5461));
    InMux I__925 (
            .O(N__5464),
            .I(N__5458));
    LocalMux I__924 (
            .O(N__5461),
            .I(\U712_CHIP_RAM.N_424 ));
    LocalMux I__923 (
            .O(N__5458),
            .I(\U712_CHIP_RAM.N_424 ));
    InMux I__922 (
            .O(N__5453),
            .I(N__5450));
    LocalMux I__921 (
            .O(N__5450),
            .I(\U712_CHIP_RAM.N_302 ));
    InMux I__920 (
            .O(N__5447),
            .I(N__5443));
    CascadeMux I__919 (
            .O(N__5446),
            .I(N__5439));
    LocalMux I__918 (
            .O(N__5443),
            .I(N__5435));
    InMux I__917 (
            .O(N__5442),
            .I(N__5428));
    InMux I__916 (
            .O(N__5439),
            .I(N__5428));
    InMux I__915 (
            .O(N__5438),
            .I(N__5428));
    Odrv4 I__914 (
            .O(N__5435),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__913 (
            .O(N__5428),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__912 (
            .O(N__5423),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_START_2_0_a2_1_cascade_ ));
    InMux I__911 (
            .O(N__5420),
            .I(N__5416));
    InMux I__910 (
            .O(N__5419),
            .I(N__5413));
    LocalMux I__909 (
            .O(N__5416),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ));
    LocalMux I__908 (
            .O(N__5413),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ));
    InMux I__907 (
            .O(N__5408),
            .I(N__5403));
    CascadeMux I__906 (
            .O(N__5407),
            .I(N__5398));
    InMux I__905 (
            .O(N__5406),
            .I(N__5392));
    LocalMux I__904 (
            .O(N__5403),
            .I(N__5388));
    InMux I__903 (
            .O(N__5402),
            .I(N__5385));
    InMux I__902 (
            .O(N__5401),
            .I(N__5376));
    InMux I__901 (
            .O(N__5398),
            .I(N__5376));
    InMux I__900 (
            .O(N__5397),
            .I(N__5376));
    InMux I__899 (
            .O(N__5396),
            .I(N__5376));
    InMux I__898 (
            .O(N__5395),
            .I(N__5373));
    LocalMux I__897 (
            .O(N__5392),
            .I(N__5370));
    InMux I__896 (
            .O(N__5391),
            .I(N__5367));
    Odrv4 I__895 (
            .O(N__5388),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__894 (
            .O(N__5385),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__893 (
            .O(N__5376),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__892 (
            .O(N__5373),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv12 I__891 (
            .O(N__5370),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__890 (
            .O(N__5367),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    CascadeMux I__889 (
            .O(N__5354),
            .I(N__5350));
    CascadeMux I__888 (
            .O(N__5353),
            .I(N__5346));
    InMux I__887 (
            .O(N__5350),
            .I(N__5343));
    InMux I__886 (
            .O(N__5349),
            .I(N__5340));
    InMux I__885 (
            .O(N__5346),
            .I(N__5335));
    LocalMux I__884 (
            .O(N__5343),
            .I(N__5331));
    LocalMux I__883 (
            .O(N__5340),
            .I(N__5328));
    InMux I__882 (
            .O(N__5339),
            .I(N__5320));
    InMux I__881 (
            .O(N__5338),
            .I(N__5317));
    LocalMux I__880 (
            .O(N__5335),
            .I(N__5314));
    InMux I__879 (
            .O(N__5334),
            .I(N__5311));
    Span4Mux_v I__878 (
            .O(N__5331),
            .I(N__5306));
    Span4Mux_v I__877 (
            .O(N__5328),
            .I(N__5306));
    InMux I__876 (
            .O(N__5327),
            .I(N__5303));
    InMux I__875 (
            .O(N__5326),
            .I(N__5300));
    InMux I__874 (
            .O(N__5325),
            .I(N__5297));
    InMux I__873 (
            .O(N__5324),
            .I(N__5292));
    InMux I__872 (
            .O(N__5323),
            .I(N__5292));
    LocalMux I__871 (
            .O(N__5320),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__870 (
            .O(N__5317),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv12 I__869 (
            .O(N__5314),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__868 (
            .O(N__5311),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__867 (
            .O(N__5306),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__866 (
            .O(N__5303),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__865 (
            .O(N__5300),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__864 (
            .O(N__5297),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__863 (
            .O(N__5292),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__862 (
            .O(N__5273),
            .I(N__5270));
    LocalMux I__861 (
            .O(N__5270),
            .I(\U712_CHIP_RAM.N_438 ));
    InMux I__860 (
            .O(N__5267),
            .I(N__5264));
    LocalMux I__859 (
            .O(N__5264),
            .I(N__5254));
    InMux I__858 (
            .O(N__5263),
            .I(N__5251));
    InMux I__857 (
            .O(N__5262),
            .I(N__5248));
    InMux I__856 (
            .O(N__5261),
            .I(N__5243));
    InMux I__855 (
            .O(N__5260),
            .I(N__5240));
    InMux I__854 (
            .O(N__5259),
            .I(N__5233));
    InMux I__853 (
            .O(N__5258),
            .I(N__5233));
    InMux I__852 (
            .O(N__5257),
            .I(N__5233));
    Span4Mux_h I__851 (
            .O(N__5254),
            .I(N__5228));
    LocalMux I__850 (
            .O(N__5251),
            .I(N__5228));
    LocalMux I__849 (
            .O(N__5248),
            .I(N__5225));
    InMux I__848 (
            .O(N__5247),
            .I(N__5220));
    InMux I__847 (
            .O(N__5246),
            .I(N__5220));
    LocalMux I__846 (
            .O(N__5243),
            .I(\U712_CHIP_RAM.N_284 ));
    LocalMux I__845 (
            .O(N__5240),
            .I(\U712_CHIP_RAM.N_284 ));
    LocalMux I__844 (
            .O(N__5233),
            .I(\U712_CHIP_RAM.N_284 ));
    Odrv4 I__843 (
            .O(N__5228),
            .I(\U712_CHIP_RAM.N_284 ));
    Odrv4 I__842 (
            .O(N__5225),
            .I(\U712_CHIP_RAM.N_284 ));
    LocalMux I__841 (
            .O(N__5220),
            .I(\U712_CHIP_RAM.N_284 ));
    CascadeMux I__840 (
            .O(N__5207),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_1_cascade_ ));
    InMux I__839 (
            .O(N__5204),
            .I(N__5197));
    InMux I__838 (
            .O(N__5203),
            .I(N__5197));
    InMux I__837 (
            .O(N__5202),
            .I(N__5193));
    LocalMux I__836 (
            .O(N__5197),
            .I(N__5190));
    InMux I__835 (
            .O(N__5196),
            .I(N__5187));
    LocalMux I__834 (
            .O(N__5193),
            .I(N__5182));
    Span4Mux_v I__833 (
            .O(N__5190),
            .I(N__5182));
    LocalMux I__832 (
            .O(N__5187),
            .I(\U712_CHIP_RAM.N_272 ));
    Odrv4 I__831 (
            .O(N__5182),
            .I(\U712_CHIP_RAM.N_272 ));
    InMux I__830 (
            .O(N__5177),
            .I(N__5174));
    LocalMux I__829 (
            .O(N__5174),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0 ));
    InMux I__828 (
            .O(N__5171),
            .I(N__5168));
    LocalMux I__827 (
            .O(N__5168),
            .I(\U712_CHIP_RAM.N_310 ));
    CascadeMux I__826 (
            .O(N__5165),
            .I(\U712_CHIP_RAM.N_310_cascade_ ));
    InMux I__825 (
            .O(N__5162),
            .I(N__5155));
    InMux I__824 (
            .O(N__5161),
            .I(N__5155));
    InMux I__823 (
            .O(N__5160),
            .I(N__5152));
    LocalMux I__822 (
            .O(N__5155),
            .I(\U712_CHIP_RAM.N_46 ));
    LocalMux I__821 (
            .O(N__5152),
            .I(\U712_CHIP_RAM.N_46 ));
    CascadeMux I__820 (
            .O(N__5147),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_3_0_a2_i_0_cascade_ ));
    CascadeMux I__819 (
            .O(N__5144),
            .I(\U712_CHIP_RAM.N_179_cascade_ ));
    IoInMux I__818 (
            .O(N__5141),
            .I(N__5138));
    LocalMux I__817 (
            .O(N__5138),
            .I(N__5135));
    IoSpan4Mux I__816 (
            .O(N__5135),
            .I(N__5132));
    Span4Mux_s3_h I__815 (
            .O(N__5132),
            .I(N__5129));
    Span4Mux_h I__814 (
            .O(N__5129),
            .I(N__5126));
    Sp12to4 I__813 (
            .O(N__5126),
            .I(N__5123));
    Span12Mux_h I__812 (
            .O(N__5123),
            .I(N__5119));
    InMux I__811 (
            .O(N__5122),
            .I(N__5116));
    Odrv12 I__810 (
            .O(N__5119),
            .I(CLK_EN_c));
    LocalMux I__809 (
            .O(N__5116),
            .I(CLK_EN_c));
    InMux I__808 (
            .O(N__5111),
            .I(N__5106));
    InMux I__807 (
            .O(N__5110),
            .I(N__5101));
    InMux I__806 (
            .O(N__5109),
            .I(N__5101));
    LocalMux I__805 (
            .O(N__5106),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    LocalMux I__804 (
            .O(N__5101),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    InMux I__803 (
            .O(N__5096),
            .I(N__5092));
    CascadeMux I__802 (
            .O(N__5095),
            .I(N__5086));
    LocalMux I__801 (
            .O(N__5092),
            .I(N__5082));
    CascadeMux I__800 (
            .O(N__5091),
            .I(N__5078));
    InMux I__799 (
            .O(N__5090),
            .I(N__5071));
    InMux I__798 (
            .O(N__5089),
            .I(N__5068));
    InMux I__797 (
            .O(N__5086),
            .I(N__5065));
    InMux I__796 (
            .O(N__5085),
            .I(N__5062));
    Span4Mux_h I__795 (
            .O(N__5082),
            .I(N__5059));
    InMux I__794 (
            .O(N__5081),
            .I(N__5056));
    InMux I__793 (
            .O(N__5078),
            .I(N__5053));
    InMux I__792 (
            .O(N__5077),
            .I(N__5048));
    InMux I__791 (
            .O(N__5076),
            .I(N__5048));
    InMux I__790 (
            .O(N__5075),
            .I(N__5043));
    InMux I__789 (
            .O(N__5074),
            .I(N__5043));
    LocalMux I__788 (
            .O(N__5071),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__787 (
            .O(N__5068),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__786 (
            .O(N__5065),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__785 (
            .O(N__5062),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__784 (
            .O(N__5059),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__783 (
            .O(N__5056),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__782 (
            .O(N__5053),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__781 (
            .O(N__5048),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__780 (
            .O(N__5043),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__779 (
            .O(N__5024),
            .I(\U712_CHIP_RAM.N_438_cascade_ ));
    CascadeMux I__778 (
            .O(N__5021),
            .I(\U712_REG_SM.N_292_cascade_ ));
    CascadeMux I__777 (
            .O(N__5018),
            .I(N__5015));
    InMux I__776 (
            .O(N__5015),
            .I(N__5011));
    InMux I__775 (
            .O(N__5014),
            .I(N__5008));
    LocalMux I__774 (
            .O(N__5011),
            .I(\U712_REG_SM.N_507 ));
    LocalMux I__773 (
            .O(N__5008),
            .I(\U712_REG_SM.N_507 ));
    InMux I__772 (
            .O(N__5003),
            .I(N__5000));
    LocalMux I__771 (
            .O(N__5000),
            .I(N__4994));
    InMux I__770 (
            .O(N__4999),
            .I(N__4991));
    InMux I__769 (
            .O(N__4998),
            .I(N__4988));
    InMux I__768 (
            .O(N__4997),
            .I(N__4985));
    Span4Mux_v I__767 (
            .O(N__4994),
            .I(N__4978));
    LocalMux I__766 (
            .O(N__4991),
            .I(N__4978));
    LocalMux I__765 (
            .O(N__4988),
            .I(N__4978));
    LocalMux I__764 (
            .O(N__4985),
            .I(N__4975));
    Span4Mux_v I__763 (
            .O(N__4978),
            .I(N__4972));
    Span4Mux_v I__762 (
            .O(N__4975),
            .I(N__4969));
    Sp12to4 I__761 (
            .O(N__4972),
            .I(N__4964));
    Sp12to4 I__760 (
            .O(N__4969),
            .I(N__4964));
    Span12Mux_h I__759 (
            .O(N__4964),
            .I(N__4961));
    Span12Mux_v I__758 (
            .O(N__4961),
            .I(N__4958));
    Odrv12 I__757 (
            .O(N__4958),
            .I(RnW_c));
    CascadeMux I__756 (
            .O(N__4955),
            .I(N__4952));
    InMux I__755 (
            .O(N__4952),
            .I(N__4949));
    LocalMux I__754 (
            .O(N__4949),
            .I(\U712_REG_SM.N_104 ));
    InMux I__753 (
            .O(N__4946),
            .I(N__4941));
    InMux I__752 (
            .O(N__4945),
            .I(N__4938));
    InMux I__751 (
            .O(N__4944),
            .I(N__4935));
    LocalMux I__750 (
            .O(N__4941),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__749 (
            .O(N__4938),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__748 (
            .O(N__4935),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    InMux I__747 (
            .O(N__4928),
            .I(N__4925));
    LocalMux I__746 (
            .O(N__4925),
            .I(\U712_REG_SM.N_372 ));
    CascadeMux I__745 (
            .O(N__4922),
            .I(N__4917));
    InMux I__744 (
            .O(N__4921),
            .I(N__4914));
    InMux I__743 (
            .O(N__4920),
            .I(N__4911));
    InMux I__742 (
            .O(N__4917),
            .I(N__4908));
    LocalMux I__741 (
            .O(N__4914),
            .I(N__4903));
    LocalMux I__740 (
            .O(N__4911),
            .I(N__4903));
    LocalMux I__739 (
            .O(N__4908),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    Odrv4 I__738 (
            .O(N__4903),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    IoInMux I__737 (
            .O(N__4898),
            .I(N__4895));
    LocalMux I__736 (
            .O(N__4895),
            .I(N__4891));
    IoInMux I__735 (
            .O(N__4894),
            .I(N__4888));
    IoSpan4Mux I__734 (
            .O(N__4891),
            .I(N__4885));
    LocalMux I__733 (
            .O(N__4888),
            .I(N__4882));
    Span4Mux_s2_v I__732 (
            .O(N__4885),
            .I(N__4879));
    IoSpan4Mux I__731 (
            .O(N__4882),
            .I(N__4876));
    Sp12to4 I__730 (
            .O(N__4879),
            .I(N__4873));
    Span4Mux_s2_v I__729 (
            .O(N__4876),
            .I(N__4870));
    Span12Mux_v I__728 (
            .O(N__4873),
            .I(N__4867));
    Sp12to4 I__727 (
            .O(N__4870),
            .I(N__4864));
    Span12Mux_h I__726 (
            .O(N__4867),
            .I(N__4859));
    Span12Mux_v I__725 (
            .O(N__4864),
            .I(N__4859));
    Odrv12 I__724 (
            .O(N__4859),
            .I(ASn_c));
    CEMux I__723 (
            .O(N__4856),
            .I(N__4853));
    LocalMux I__722 (
            .O(N__4853),
            .I(\U712_REG_SM.N_186_0 ));
    CascadeMux I__721 (
            .O(N__4850),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_cascade_ ));
    CascadeMux I__720 (
            .O(N__4847),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_0_a2_2_cascade_ ));
    CascadeMux I__719 (
            .O(N__4844),
            .I(N__4841));
    InMux I__718 (
            .O(N__4841),
            .I(N__4838));
    LocalMux I__717 (
            .O(N__4838),
            .I(\U712_CHIP_RAM.N_393 ));
    InMux I__716 (
            .O(N__4835),
            .I(N__4829));
    InMux I__715 (
            .O(N__4834),
            .I(N__4824));
    InMux I__714 (
            .O(N__4833),
            .I(N__4824));
    InMux I__713 (
            .O(N__4832),
            .I(N__4821));
    LocalMux I__712 (
            .O(N__4829),
            .I(N__4818));
    LocalMux I__711 (
            .O(N__4824),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    LocalMux I__710 (
            .O(N__4821),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    Odrv4 I__709 (
            .O(N__4818),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    CascadeMux I__708 (
            .O(N__4811),
            .I(\U712_REG_SM.N_301_cascade_ ));
    CascadeMux I__707 (
            .O(N__4808),
            .I(N__4804));
    CascadeMux I__706 (
            .O(N__4807),
            .I(N__4801));
    InMux I__705 (
            .O(N__4804),
            .I(N__4797));
    InMux I__704 (
            .O(N__4801),
            .I(N__4794));
    InMux I__703 (
            .O(N__4800),
            .I(N__4791));
    LocalMux I__702 (
            .O(N__4797),
            .I(\U712_REG_SM.N_288 ));
    LocalMux I__701 (
            .O(N__4794),
            .I(\U712_REG_SM.N_288 ));
    LocalMux I__700 (
            .O(N__4791),
            .I(\U712_REG_SM.N_288 ));
    InMux I__699 (
            .O(N__4784),
            .I(N__4779));
    InMux I__698 (
            .O(N__4783),
            .I(N__4776));
    InMux I__697 (
            .O(N__4782),
            .I(N__4773));
    LocalMux I__696 (
            .O(N__4779),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__695 (
            .O(N__4776),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__694 (
            .O(N__4773),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    InMux I__693 (
            .O(N__4766),
            .I(N__4760));
    InMux I__692 (
            .O(N__4765),
            .I(N__4760));
    LocalMux I__691 (
            .O(N__4760),
            .I(\U712_REG_SM.N_301 ));
    InMux I__690 (
            .O(N__4757),
            .I(N__4748));
    InMux I__689 (
            .O(N__4756),
            .I(N__4748));
    InMux I__688 (
            .O(N__4755),
            .I(N__4748));
    LocalMux I__687 (
            .O(N__4748),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    InMux I__686 (
            .O(N__4745),
            .I(N__4742));
    LocalMux I__685 (
            .O(N__4742),
            .I(N__4739));
    Span4Mux_v I__684 (
            .O(N__4739),
            .I(N__4733));
    InMux I__683 (
            .O(N__4738),
            .I(N__4726));
    InMux I__682 (
            .O(N__4737),
            .I(N__4726));
    InMux I__681 (
            .O(N__4736),
            .I(N__4726));
    Odrv4 I__680 (
            .O(N__4733),
            .I(REG_CYCLEm));
    LocalMux I__679 (
            .O(N__4726),
            .I(REG_CYCLEm));
    IoInMux I__678 (
            .O(N__4721),
            .I(N__4718));
    LocalMux I__677 (
            .O(N__4718),
            .I(N__4715));
    IoSpan4Mux I__676 (
            .O(N__4715),
            .I(N__4712));
    IoSpan4Mux I__675 (
            .O(N__4712),
            .I(N__4709));
    IoSpan4Mux I__674 (
            .O(N__4709),
            .I(N__4706));
    Span4Mux_s3_v I__673 (
            .O(N__4706),
            .I(N__4703));
    Sp12to4 I__672 (
            .O(N__4703),
            .I(N__4700));
    Span12Mux_v I__671 (
            .O(N__4700),
            .I(N__4697));
    Odrv12 I__670 (
            .O(N__4697),
            .I(DRDENn_c));
    CascadeMux I__669 (
            .O(N__4694),
            .I(N__4691));
    InMux I__668 (
            .O(N__4691),
            .I(N__4687));
    InMux I__667 (
            .O(N__4690),
            .I(N__4684));
    LocalMux I__666 (
            .O(N__4687),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__665 (
            .O(N__4684),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    InMux I__664 (
            .O(N__4679),
            .I(N__4673));
    InMux I__663 (
            .O(N__4678),
            .I(N__4673));
    LocalMux I__662 (
            .O(N__4673),
            .I(\U712_REG_SM.N_341 ));
    CascadeMux I__661 (
            .O(N__4670),
            .I(\U712_REG_SM.N_294_cascade_ ));
    InMux I__660 (
            .O(N__4667),
            .I(N__4664));
    LocalMux I__659 (
            .O(N__4664),
            .I(N__4661));
    Odrv4 I__658 (
            .O(N__4661),
            .I(\U712_REG_SM.N_373 ));
    InMux I__657 (
            .O(N__4658),
            .I(N__4652));
    InMux I__656 (
            .O(N__4657),
            .I(N__4652));
    LocalMux I__655 (
            .O(N__4652),
            .I(N__4649));
    Odrv4 I__654 (
            .O(N__4649),
            .I(\U712_CHIP_RAM.N_296_i ));
    CascadeMux I__653 (
            .O(N__4646),
            .I(\U712_CHIP_RAM.SDRAM_CMD_e_1_2_cascade_ ));
    CascadeMux I__652 (
            .O(N__4643),
            .I(N__4640));
    InMux I__651 (
            .O(N__4640),
            .I(N__4637));
    LocalMux I__650 (
            .O(N__4637),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_0_3 ));
    CEMux I__649 (
            .O(N__4634),
            .I(N__4631));
    LocalMux I__648 (
            .O(N__4631),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0 ));
    IoInMux I__647 (
            .O(N__4628),
            .I(N__4625));
    LocalMux I__646 (
            .O(N__4625),
            .I(N__4622));
    Span4Mux_s2_v I__645 (
            .O(N__4622),
            .I(N__4618));
    CascadeMux I__644 (
            .O(N__4621),
            .I(N__4615));
    Sp12to4 I__643 (
            .O(N__4618),
            .I(N__4611));
    InMux I__642 (
            .O(N__4615),
            .I(N__4608));
    CascadeMux I__641 (
            .O(N__4614),
            .I(N__4605));
    Span12Mux_h I__640 (
            .O(N__4611),
            .I(N__4602));
    LocalMux I__639 (
            .O(N__4608),
            .I(N__4599));
    InMux I__638 (
            .O(N__4605),
            .I(N__4596));
    Odrv12 I__637 (
            .O(N__4602),
            .I(DBDIR_c));
    Odrv4 I__636 (
            .O(N__4599),
            .I(DBDIR_c));
    LocalMux I__635 (
            .O(N__4596),
            .I(DBDIR_c));
    IoInMux I__634 (
            .O(N__4589),
            .I(N__4586));
    LocalMux I__633 (
            .O(N__4586),
            .I(N__4583));
    IoSpan4Mux I__632 (
            .O(N__4583),
            .I(N__4580));
    Span4Mux_s2_h I__631 (
            .O(N__4580),
            .I(N__4577));
    Sp12to4 I__630 (
            .O(N__4577),
            .I(N__4574));
    Span12Mux_s11_h I__629 (
            .O(N__4574),
            .I(N__4571));
    Span12Mux_v I__628 (
            .O(N__4571),
            .I(N__4568));
    Odrv12 I__627 (
            .O(N__4568),
            .I(N_188));
    InMux I__626 (
            .O(N__4565),
            .I(N__4562));
    LocalMux I__625 (
            .O(N__4562),
            .I(N__4559));
    Span4Mux_v I__624 (
            .O(N__4559),
            .I(N__4554));
    InMux I__623 (
            .O(N__4558),
            .I(N__4549));
    InMux I__622 (
            .O(N__4557),
            .I(N__4549));
    Odrv4 I__621 (
            .O(N__4554),
            .I(U712_REG_SM_DBR_SYNC_1));
    LocalMux I__620 (
            .O(N__4549),
            .I(U712_REG_SM_DBR_SYNC_1));
    CascadeMux I__619 (
            .O(N__4544),
            .I(\U712_REG_SM.N_288_cascade_ ));
    InMux I__618 (
            .O(N__4541),
            .I(N__4538));
    LocalMux I__617 (
            .O(N__4538),
            .I(N__4534));
    InMux I__616 (
            .O(N__4537),
            .I(N__4529));
    Span4Mux_v I__615 (
            .O(N__4534),
            .I(N__4526));
    InMux I__614 (
            .O(N__4533),
            .I(N__4521));
    InMux I__613 (
            .O(N__4532),
            .I(N__4521));
    LocalMux I__612 (
            .O(N__4529),
            .I(U712_REG_SM_DBR_SYNC_0));
    Odrv4 I__611 (
            .O(N__4526),
            .I(U712_REG_SM_DBR_SYNC_0));
    LocalMux I__610 (
            .O(N__4521),
            .I(U712_REG_SM_DBR_SYNC_0));
    CascadeMux I__609 (
            .O(N__4514),
            .I(\U712_CHIP_RAM.N_347_cascade_ ));
    CascadeMux I__608 (
            .O(N__4511),
            .I(\U712_CHIP_RAM.N_378_cascade_ ));
    InMux I__607 (
            .O(N__4508),
            .I(N__4505));
    LocalMux I__606 (
            .O(N__4505),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_tz ));
    InMux I__605 (
            .O(N__4502),
            .I(N__4499));
    LocalMux I__604 (
            .O(N__4499),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_0_a2_0_a2_0 ));
    CascadeMux I__603 (
            .O(N__4496),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_0_cascade_ ));
    CascadeMux I__602 (
            .O(N__4493),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER50_cascade_ ));
    InMux I__601 (
            .O(N__4490),
            .I(N__4486));
    InMux I__600 (
            .O(N__4489),
            .I(N__4483));
    LocalMux I__599 (
            .O(N__4486),
            .I(N__4478));
    LocalMux I__598 (
            .O(N__4483),
            .I(N__4478));
    Span12Mux_h I__597 (
            .O(N__4478),
            .I(N__4475));
    Span12Mux_v I__596 (
            .O(N__4475),
            .I(N__4472));
    Odrv12 I__595 (
            .O(N__4472),
            .I(AWEn_c));
    InMux I__594 (
            .O(N__4469),
            .I(N__4466));
    LocalMux I__593 (
            .O(N__4466),
            .I(\U712_CHIP_RAM.N_287 ));
    CascadeMux I__592 (
            .O(N__4463),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_1_0_cascade_ ));
    CascadeMux I__591 (
            .O(N__4460),
            .I(\U712_CHIP_RAM.N_273_cascade_ ));
    InMux I__590 (
            .O(N__4457),
            .I(N__4452));
    InMux I__589 (
            .O(N__4456),
            .I(N__4449));
    InMux I__588 (
            .O(N__4455),
            .I(N__4446));
    LocalMux I__587 (
            .O(N__4452),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3 ));
    LocalMux I__586 (
            .O(N__4449),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3 ));
    LocalMux I__585 (
            .O(N__4446),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3 ));
    InMux I__584 (
            .O(N__4439),
            .I(N__4436));
    LocalMux I__583 (
            .O(N__4436),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_0 ));
    InMux I__582 (
            .O(N__4433),
            .I(N__4429));
    CascadeMux I__581 (
            .O(N__4432),
            .I(N__4425));
    LocalMux I__580 (
            .O(N__4429),
            .I(N__4421));
    InMux I__579 (
            .O(N__4428),
            .I(N__4414));
    InMux I__578 (
            .O(N__4425),
            .I(N__4414));
    InMux I__577 (
            .O(N__4424),
            .I(N__4414));
    Span4Mux_v I__576 (
            .O(N__4421),
            .I(N__4411));
    LocalMux I__575 (
            .O(N__4414),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    Odrv4 I__574 (
            .O(N__4411),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__573 (
            .O(N__4406),
            .I(N__4403));
    LocalMux I__572 (
            .O(N__4403),
            .I(N__4398));
    InMux I__571 (
            .O(N__4402),
            .I(N__4393));
    InMux I__570 (
            .O(N__4401),
            .I(N__4393));
    Odrv4 I__569 (
            .O(N__4398),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__568 (
            .O(N__4393),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    CascadeMux I__567 (
            .O(N__4388),
            .I(N__4384));
    CascadeMux I__566 (
            .O(N__4387),
            .I(N__4381));
    InMux I__565 (
            .O(N__4384),
            .I(N__4376));
    InMux I__564 (
            .O(N__4381),
            .I(N__4376));
    LocalMux I__563 (
            .O(N__4376),
            .I(\U712_REG_SM.LDS_OUT_2_0_a2Z0Z_0 ));
    CascadeMux I__562 (
            .O(N__4373),
            .I(N__4370));
    InMux I__561 (
            .O(N__4370),
            .I(N__4367));
    LocalMux I__560 (
            .O(N__4367),
            .I(N__4360));
    InMux I__559 (
            .O(N__4366),
            .I(N__4357));
    InMux I__558 (
            .O(N__4365),
            .I(N__4350));
    InMux I__557 (
            .O(N__4364),
            .I(N__4350));
    InMux I__556 (
            .O(N__4363),
            .I(N__4350));
    Odrv4 I__555 (
            .O(N__4360),
            .I(\U712_REG_SM.N_342 ));
    LocalMux I__554 (
            .O(N__4357),
            .I(\U712_REG_SM.N_342 ));
    LocalMux I__553 (
            .O(N__4350),
            .I(\U712_REG_SM.N_342 ));
    InMux I__552 (
            .O(N__4343),
            .I(N__4339));
    InMux I__551 (
            .O(N__4342),
            .I(N__4336));
    LocalMux I__550 (
            .O(N__4339),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    LocalMux I__549 (
            .O(N__4336),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    IoInMux I__548 (
            .O(N__4331),
            .I(N__4328));
    LocalMux I__547 (
            .O(N__4328),
            .I(N__4325));
    IoSpan4Mux I__546 (
            .O(N__4325),
            .I(N__4322));
    Span4Mux_s3_v I__545 (
            .O(N__4322),
            .I(N__4319));
    Span4Mux_h I__544 (
            .O(N__4319),
            .I(N__4316));
    Sp12to4 I__543 (
            .O(N__4316),
            .I(N__4313));
    Span12Mux_v I__542 (
            .O(N__4313),
            .I(N__4310));
    Odrv12 I__541 (
            .O(N__4310),
            .I(U712_REG_SM_un1_LDSn_i));
    InMux I__540 (
            .O(N__4307),
            .I(N__4304));
    LocalMux I__539 (
            .O(N__4304),
            .I(N__4300));
    InMux I__538 (
            .O(N__4303),
            .I(N__4297));
    Odrv4 I__537 (
            .O(N__4300),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    LocalMux I__536 (
            .O(N__4297),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    InMux I__535 (
            .O(N__4292),
            .I(N__4288));
    InMux I__534 (
            .O(N__4291),
            .I(N__4285));
    LocalMux I__533 (
            .O(N__4288),
            .I(N__4281));
    LocalMux I__532 (
            .O(N__4285),
            .I(N__4278));
    InMux I__531 (
            .O(N__4284),
            .I(N__4275));
    Odrv12 I__530 (
            .O(N__4281),
            .I(\U712_REG_SM.DS_ENZ0 ));
    Odrv4 I__529 (
            .O(N__4278),
            .I(\U712_REG_SM.DS_ENZ0 ));
    LocalMux I__528 (
            .O(N__4275),
            .I(\U712_REG_SM.DS_ENZ0 ));
    IoInMux I__527 (
            .O(N__4268),
            .I(N__4265));
    LocalMux I__526 (
            .O(N__4265),
            .I(N__4262));
    IoSpan4Mux I__525 (
            .O(N__4262),
            .I(N__4259));
    IoSpan4Mux I__524 (
            .O(N__4259),
            .I(N__4256));
    Sp12to4 I__523 (
            .O(N__4256),
            .I(N__4253));
    Span12Mux_v I__522 (
            .O(N__4253),
            .I(N__4250));
    Odrv12 I__521 (
            .O(N__4250),
            .I(U712_REG_SM_un1_UDSn_i));
    CascadeMux I__520 (
            .O(N__4247),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_ ));
    CascadeMux I__519 (
            .O(N__4244),
            .I(N__4241));
    InMux I__518 (
            .O(N__4241),
            .I(N__4238));
    LocalMux I__517 (
            .O(N__4238),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6 ));
    InMux I__516 (
            .O(N__4235),
            .I(N__4231));
    InMux I__515 (
            .O(N__4234),
            .I(N__4228));
    LocalMux I__514 (
            .O(N__4231),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__513 (
            .O(N__4228),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__512 (
            .O(N__4223),
            .I(N__4218));
    InMux I__511 (
            .O(N__4222),
            .I(N__4215));
    InMux I__510 (
            .O(N__4221),
            .I(N__4212));
    LocalMux I__509 (
            .O(N__4218),
            .I(N__4209));
    LocalMux I__508 (
            .O(N__4215),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__507 (
            .O(N__4212),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    Odrv4 I__506 (
            .O(N__4209),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__505 (
            .O(N__4202),
            .I(N__4197));
    InMux I__504 (
            .O(N__4201),
            .I(N__4192));
    InMux I__503 (
            .O(N__4200),
            .I(N__4192));
    InMux I__502 (
            .O(N__4197),
            .I(N__4189));
    LocalMux I__501 (
            .O(N__4192),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__500 (
            .O(N__4189),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    CascadeMux I__499 (
            .O(N__4184),
            .I(N__4181));
    InMux I__498 (
            .O(N__4181),
            .I(N__4175));
    InMux I__497 (
            .O(N__4180),
            .I(N__4172));
    InMux I__496 (
            .O(N__4179),
            .I(N__4169));
    InMux I__495 (
            .O(N__4178),
            .I(N__4166));
    LocalMux I__494 (
            .O(N__4175),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__493 (
            .O(N__4172),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__492 (
            .O(N__4169),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__491 (
            .O(N__4166),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__490 (
            .O(N__4157),
            .I(N__4154));
    InMux I__489 (
            .O(N__4154),
            .I(N__4150));
    InMux I__488 (
            .O(N__4153),
            .I(N__4147));
    LocalMux I__487 (
            .O(N__4150),
            .I(REG_TACK));
    LocalMux I__486 (
            .O(N__4147),
            .I(REG_TACK));
    InMux I__485 (
            .O(N__4142),
            .I(N__4139));
    LocalMux I__484 (
            .O(N__4139),
            .I(N__4135));
    InMux I__483 (
            .O(N__4138),
            .I(N__4132));
    Span4Mux_v I__482 (
            .O(N__4135),
            .I(N__4127));
    LocalMux I__481 (
            .O(N__4132),
            .I(N__4127));
    Span4Mux_v I__480 (
            .O(N__4127),
            .I(N__4124));
    Span4Mux_v I__479 (
            .O(N__4124),
            .I(N__4121));
    Sp12to4 I__478 (
            .O(N__4121),
            .I(N__4118));
    Span12Mux_h I__477 (
            .O(N__4118),
            .I(N__4115));
    Odrv12 I__476 (
            .O(N__4115),
            .I(TSn_c));
    InMux I__475 (
            .O(N__4112),
            .I(N__4109));
    LocalMux I__474 (
            .O(N__4109),
            .I(N__4106));
    Span4Mux_v I__473 (
            .O(N__4106),
            .I(N__4103));
    Sp12to4 I__472 (
            .O(N__4103),
            .I(N__4100));
    Span12Mux_h I__471 (
            .O(N__4100),
            .I(N__4097));
    Span12Mux_v I__470 (
            .O(N__4097),
            .I(N__4094));
    Odrv12 I__469 (
            .O(N__4094),
            .I(REGSPACEn_c));
    InMux I__468 (
            .O(N__4091),
            .I(N__4085));
    InMux I__467 (
            .O(N__4090),
            .I(N__4085));
    LocalMux I__466 (
            .O(N__4085),
            .I(\U712_REG_SM.REG_CYCLE_GOZ0 ));
    InMux I__465 (
            .O(N__4082),
            .I(N__4079));
    LocalMux I__464 (
            .O(N__4079),
            .I(\U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1 ));
    CascadeMux I__463 (
            .O(N__4076),
            .I(\U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_ ));
    CascadeMux I__462 (
            .O(N__4073),
            .I(N__4070));
    InMux I__461 (
            .O(N__4070),
            .I(N__4067));
    LocalMux I__460 (
            .O(N__4067),
            .I(N__4064));
    Span4Mux_v I__459 (
            .O(N__4064),
            .I(N__4061));
    Sp12to4 I__458 (
            .O(N__4061),
            .I(N__4058));
    Span12Mux_h I__457 (
            .O(N__4058),
            .I(N__4055));
    Span12Mux_v I__456 (
            .O(N__4055),
            .I(N__4052));
    Odrv12 I__455 (
            .O(N__4052),
            .I(RAMSPACEn_c));
    InMux I__454 (
            .O(N__4049),
            .I(N__4046));
    LocalMux I__453 (
            .O(N__4046),
            .I(N__4043));
    Span4Mux_v I__452 (
            .O(N__4043),
            .I(N__4040));
    Sp12to4 I__451 (
            .O(N__4040),
            .I(N__4037));
    Span12Mux_h I__450 (
            .O(N__4037),
            .I(N__4034));
    Span12Mux_v I__449 (
            .O(N__4034),
            .I(N__4031));
    Odrv12 I__448 (
            .O(N__4031),
            .I(DBRn_c));
    CascadeMux I__447 (
            .O(N__4028),
            .I(\U712_CHIP_RAM.N_287_cascade_ ));
    InMux I__446 (
            .O(N__4025),
            .I(N__4022));
    LocalMux I__445 (
            .O(N__4022),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_1_0 ));
    CascadeMux I__444 (
            .O(N__4019),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_cascade_ ));
    CascadeMux I__443 (
            .O(N__4016),
            .I(N__4013));
    InMux I__442 (
            .O(N__4013),
            .I(N__4006));
    InMux I__441 (
            .O(N__4012),
            .I(N__4006));
    InMux I__440 (
            .O(N__4011),
            .I(N__4003));
    LocalMux I__439 (
            .O(N__4006),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__438 (
            .O(N__4003),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__437 (
            .O(N__3998),
            .I(N__3994));
    InMux I__436 (
            .O(N__3997),
            .I(N__3991));
    LocalMux I__435 (
            .O(N__3994),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    LocalMux I__434 (
            .O(N__3991),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__433 (
            .O(N__3986),
            .I(N__3983));
    LocalMux I__432 (
            .O(N__3983),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ));
    CascadeMux I__431 (
            .O(N__3980),
            .I(\U712_CYCLE_TERM.N_307_i_0_en_cascade_ ));
    InMux I__430 (
            .O(N__3977),
            .I(N__3972));
    InMux I__429 (
            .O(N__3976),
            .I(N__3967));
    InMux I__428 (
            .O(N__3975),
            .I(N__3967));
    LocalMux I__427 (
            .O(N__3972),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__426 (
            .O(N__3967),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CascadeMux I__425 (
            .O(N__3962),
            .I(N__3958));
    InMux I__424 (
            .O(N__3961),
            .I(N__3955));
    InMux I__423 (
            .O(N__3958),
            .I(N__3951));
    LocalMux I__422 (
            .O(N__3955),
            .I(N__3948));
    InMux I__421 (
            .O(N__3954),
            .I(N__3945));
    LocalMux I__420 (
            .O(N__3951),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    Odrv4 I__419 (
            .O(N__3948),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__418 (
            .O(N__3945),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__417 (
            .O(N__3938),
            .I(N__3935));
    LocalMux I__416 (
            .O(N__3935),
            .I(N__3932));
    Sp12to4 I__415 (
            .O(N__3932),
            .I(N__3929));
    Odrv12 I__414 (
            .O(N__3929),
            .I(TACK_EN_i_ess));
    CEMux I__413 (
            .O(N__3926),
            .I(N__3923));
    LocalMux I__412 (
            .O(N__3923),
            .I(N__3920));
    Odrv12 I__411 (
            .O(N__3920),
            .I(\U712_CYCLE_TERM.N_307_i_0_en_0 ));
    IoInMux I__410 (
            .O(N__3917),
            .I(N__3914));
    LocalMux I__409 (
            .O(N__3914),
            .I(N__3911));
    Span12Mux_s2_v I__408 (
            .O(N__3911),
            .I(N__3908));
    Odrv12 I__407 (
            .O(N__3908),
            .I(VBENn_c));
    CascadeMux I__406 (
            .O(N__3905),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3_cascade_ ));
    CascadeMux I__405 (
            .O(N__3902),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_ ));
    InMux I__404 (
            .O(N__3899),
            .I(N__3896));
    LocalMux I__403 (
            .O(N__3896),
            .I(\U712_CHIP_RAM.N_181 ));
    InMux I__402 (
            .O(N__3893),
            .I(N__3883));
    InMux I__401 (
            .O(N__3892),
            .I(N__3883));
    InMux I__400 (
            .O(N__3891),
            .I(N__3883));
    InMux I__399 (
            .O(N__3890),
            .I(N__3880));
    LocalMux I__398 (
            .O(N__3883),
            .I(N__3877));
    LocalMux I__397 (
            .O(N__3880),
            .I(N__3872));
    Span4Mux_v I__396 (
            .O(N__3877),
            .I(N__3872));
    Span4Mux_v I__395 (
            .O(N__3872),
            .I(N__3869));
    Sp12to4 I__394 (
            .O(N__3869),
            .I(N__3866));
    Span12Mux_h I__393 (
            .O(N__3866),
            .I(N__3863));
    Odrv12 I__392 (
            .O(N__3863),
            .I(CLK40_OUT_i));
    IoInMux I__391 (
            .O(N__3860),
            .I(N__3857));
    LocalMux I__390 (
            .O(N__3857),
            .I(N__3854));
    Span12Mux_s8_h I__389 (
            .O(N__3854),
            .I(N__3851));
    Span12Mux_v I__388 (
            .O(N__3851),
            .I(N__3847));
    InMux I__387 (
            .O(N__3850),
            .I(N__3844));
    Odrv12 I__386 (
            .O(N__3847),
            .I(TACK_OUTn));
    LocalMux I__385 (
            .O(N__3844),
            .I(TACK_OUTn));
    InMux I__384 (
            .O(N__3839),
            .I(N__3827));
    InMux I__383 (
            .O(N__3838),
            .I(N__3827));
    InMux I__382 (
            .O(N__3837),
            .I(N__3827));
    InMux I__381 (
            .O(N__3836),
            .I(N__3827));
    LocalMux I__380 (
            .O(N__3827),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__379 (
            .O(N__3824),
            .I(N__3820));
    InMux I__378 (
            .O(N__3823),
            .I(N__3817));
    LocalMux I__377 (
            .O(N__3820),
            .I(CPU_TACKm));
    LocalMux I__376 (
            .O(N__3817),
            .I(CPU_TACKm));
    CascadeMux I__375 (
            .O(N__3812),
            .I(N__3809));
    InMux I__374 (
            .O(N__3809),
            .I(N__3805));
    InMux I__373 (
            .O(N__3808),
            .I(N__3802));
    LocalMux I__372 (
            .O(N__3805),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__371 (
            .O(N__3802),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__370 (
            .O(N__3797),
            .I(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ));
    InMux I__369 (
            .O(N__3794),
            .I(N__3791));
    LocalMux I__368 (
            .O(N__3791),
            .I(N__3788));
    Span4Mux_v I__367 (
            .O(N__3788),
            .I(N__3785));
    Sp12to4 I__366 (
            .O(N__3785),
            .I(N__3782));
    Odrv12 I__365 (
            .O(N__3782),
            .I(A_c_13));
    CascadeMux I__364 (
            .O(N__3779),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4_cascade_ ));
    InMux I__363 (
            .O(N__3776),
            .I(N__3773));
    LocalMux I__362 (
            .O(N__3773),
            .I(N__3770));
    Span4Mux_h I__361 (
            .O(N__3770),
            .I(N__3767));
    Sp12to4 I__360 (
            .O(N__3767),
            .I(N__3764));
    Span12Mux_v I__359 (
            .O(N__3764),
            .I(N__3761));
    Odrv12 I__358 (
            .O(N__3761),
            .I(A_c_6));
    IoInMux I__357 (
            .O(N__3758),
            .I(N__3755));
    LocalMux I__356 (
            .O(N__3755),
            .I(N__3752));
    Span12Mux_s9_h I__355 (
            .O(N__3752),
            .I(N__3749));
    Span12Mux_h I__354 (
            .O(N__3749),
            .I(N__3746));
    Odrv12 I__353 (
            .O(N__3746),
            .I(CMA_c_3));
    InMux I__352 (
            .O(N__3743),
            .I(N__3740));
    LocalMux I__351 (
            .O(N__3740),
            .I(\U712_CHIP_RAM.N_319 ));
    IoInMux I__350 (
            .O(N__3737),
            .I(N__3734));
    LocalMux I__349 (
            .O(N__3734),
            .I(N__3731));
    Span4Mux_s2_h I__348 (
            .O(N__3731),
            .I(N__3728));
    Span4Mux_v I__347 (
            .O(N__3728),
            .I(N__3725));
    Span4Mux_v I__346 (
            .O(N__3725),
            .I(N__3722));
    Sp12to4 I__345 (
            .O(N__3722),
            .I(N__3719));
    Span12Mux_s11_h I__344 (
            .O(N__3719),
            .I(N__3716));
    Odrv12 I__343 (
            .O(N__3716),
            .I(CMA_c_4));
    InMux I__342 (
            .O(N__3713),
            .I(N__3710));
    LocalMux I__341 (
            .O(N__3710),
            .I(N__3707));
    Span4Mux_v I__340 (
            .O(N__3707),
            .I(N__3704));
    Sp12to4 I__339 (
            .O(N__3704),
            .I(N__3701));
    Odrv12 I__338 (
            .O(N__3701),
            .I(A_c_12));
    CascadeMux I__337 (
            .O(N__3698),
            .I(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_ ));
    InMux I__336 (
            .O(N__3695),
            .I(N__3692));
    LocalMux I__335 (
            .O(N__3692),
            .I(N__3689));
    Sp12to4 I__334 (
            .O(N__3689),
            .I(N__3686));
    Span12Mux_v I__333 (
            .O(N__3686),
            .I(N__3683));
    Odrv12 I__332 (
            .O(N__3683),
            .I(A_c_5));
    InMux I__331 (
            .O(N__3680),
            .I(N__3677));
    LocalMux I__330 (
            .O(N__3677),
            .I(\U712_CHIP_RAM.N_318 ));
    IoInMux I__329 (
            .O(N__3674),
            .I(N__3671));
    LocalMux I__328 (
            .O(N__3671),
            .I(N__3668));
    Span4Mux_s3_h I__327 (
            .O(N__3668),
            .I(N__3665));
    Span4Mux_h I__326 (
            .O(N__3665),
            .I(N__3662));
    Span4Mux_v I__325 (
            .O(N__3662),
            .I(N__3659));
    Odrv4 I__324 (
            .O(N__3659),
            .I(CLK40_OUT_i_i));
    CascadeMux I__323 (
            .O(N__3656),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_0_a2_i_0_cascade_ ));
    IoInMux I__322 (
            .O(N__3653),
            .I(N__3650));
    LocalMux I__321 (
            .O(N__3650),
            .I(N__3647));
    IoSpan4Mux I__320 (
            .O(N__3647),
            .I(N__3644));
    Span4Mux_s2_v I__319 (
            .O(N__3644),
            .I(N__3641));
    Span4Mux_v I__318 (
            .O(N__3641),
            .I(N__3638));
    Odrv4 I__317 (
            .O(N__3638),
            .I(CLK80_OUT_i_i));
    IoInMux I__316 (
            .O(N__3635),
            .I(N__3632));
    LocalMux I__315 (
            .O(N__3632),
            .I(N__3629));
    IoSpan4Mux I__314 (
            .O(N__3629),
            .I(N__3626));
    Span4Mux_s3_h I__313 (
            .O(N__3626),
            .I(N__3623));
    Span4Mux_h I__312 (
            .O(N__3623),
            .I(N__3620));
    Odrv4 I__311 (
            .O(N__3620),
            .I(N_839_i));
    IoInMux I__310 (
            .O(N__3617),
            .I(N__3614));
    LocalMux I__309 (
            .O(N__3614),
            .I(N__3611));
    IoSpan4Mux I__308 (
            .O(N__3611),
            .I(N__3608));
    Span4Mux_s2_v I__307 (
            .O(N__3608),
            .I(N__3605));
    Sp12to4 I__306 (
            .O(N__3605),
            .I(N__3602));
    Span12Mux_v I__305 (
            .O(N__3602),
            .I(N__3599));
    Odrv12 I__304 (
            .O(N__3599),
            .I(CLK40_IN_c));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_8_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7634),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__6169),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_5_1_5.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_5_1_5.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_5_1_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_5_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9248),
            .lcout(CLK80_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_obuft_RNO_LC_6_18_0.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_6_18_0.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_6_18_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_obuft_RNO_LC_6_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3938),
            .lcout(N_839_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_7_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_7_4_6 .LUT_INIT=16'b0000111101010011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_7_4_6  (
            .in0(N__7583),
            .in1(N__6818),
            .in2(N__8521),
            .in3(N__8134),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_7_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_7_4_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_7_4_7  (
            .in0(N__8135),
            .in1(N__3794),
            .in2(N__3779),
            .in3(N__3776),
            .lcout(\U712_CHIP_RAM.N_319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_7_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_7_5_3 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_7_5_3  (
            .in0(N__3680),
            .in1(_gnd_net_),
            .in2(N__8641),
            .in3(N__8756),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9231),
            .ce(N__7967),
            .sr(N__9046));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_7_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_7_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_7_5_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_7_5_6  (
            .in0(N__8755),
            .in1(N__8631),
            .in2(_gnd_net_),
            .in3(N__3743),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9231),
            .ce(N__7967),
            .sr(N__9046));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_7_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_7_6_0 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_7_6_0  (
            .in0(N__8507),
            .in1(N__7880),
            .in2(N__8169),
            .in3(N__7466),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_7_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_7_6_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_7_6_1  (
            .in0(N__8158),
            .in1(N__3713),
            .in2(N__3698),
            .in3(N__3695),
            .lcout(\U712_CHIP_RAM.N_318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLK40C_obuf_RNO_LC_7_6_5.C_ON=1'b0;
    defparam CLK40C_obuf_RNO_LC_7_6_5.SEQ_MODE=4'b0000;
    defparam CLK40C_obuf_RNO_LC_7_6_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLK40C_obuf_RNO_LC_7_6_5 (
            .in0(N__3890),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_8_6 .LUT_INIT=16'b1001100110111011;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_8_6  (
            .in0(N__5800),
            .in1(N__5656),
            .in2(_gnd_net_),
            .in3(N__5349),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_0_a2_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_8_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_8_7  (
            .in0(N__5267),
            .in1(N__7203),
            .in2(N__3656),
            .in3(N__5096),
            .lcout(\U712_CHIP_RAM.N_181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_7_9_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_7_9_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_7_9_0  (
            .in0(N__3837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3893),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9239),
            .ce(),
            .sr(N__9019));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_7_9_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_7_9_1 .LUT_INIT=16'b1111101000110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_7_9_1  (
            .in0(N__3891),
            .in1(N__3976),
            .in2(N__3962),
            .in3(N__3839),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9239),
            .ce(),
            .sr(N__9019));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_7_9_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_7_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3998),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9239),
            .ce(),
            .sr(N__9019));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_7_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_7_9_3 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_7_9_3  (
            .in0(N__3824),
            .in1(N__5801),
            .in2(N__8174),
            .in3(N__3899),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9239),
            .ce(),
            .sr(N__9019));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_7_9_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_7_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4012),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9239),
            .ce(),
            .sr(N__9019));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_7_9_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_7_9_6 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_7_9_6 .LUT_INIT=16'b1111110011110100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_7_9_6  (
            .in0(N__3838),
            .in1(N__3850),
            .in2(N__4016),
            .in3(N__3892),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9239),
            .ce(),
            .sr(N__9019));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_7_9_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_7_9_7 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_7_9_7 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_7_9_7  (
            .in0(N__3986),
            .in1(N__3975),
            .in2(N__3812),
            .in3(N__3836),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9239),
            .ce(),
            .sr(N__9019));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_7_10_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_7_10_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(N__4153),
            .in2(_gnd_net_),
            .in3(N__3823),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_7_10_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_7_10_5 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_7_10_5  (
            .in0(N__7701),
            .in1(N__3808),
            .in2(N__3797),
            .in3(N__3954),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_307_i_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_7_10_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_7_10_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_7_10_6  (
            .in0(N__9083),
            .in1(_gnd_net_),
            .in2(N__3980),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.N_307_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_11_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_11_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_11_0 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_11_0  (
            .in0(N__7691),
            .in1(N__3977),
            .in2(_gnd_net_),
            .in3(N__3961),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9243),
            .ce(N__3926),
            .sr(N__9004));
    defparam \U712_REG_SM.LDS_OUT_2_0_a2_0_LC_7_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_2_0_a2_0_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_2_0_a2_0_LC_7_12_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_REG_SM.LDS_OUT_2_0_a2_0_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__6058),
            .in2(_gnd_net_),
            .in3(N__4997),
            .lcout(\U712_REG_SM.LDS_OUT_2_0_a2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_4_3 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_4_3  (
            .in0(N__4457),
            .in1(N__9089),
            .in2(N__4184),
            .in3(N__5090),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9222),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_5  (
            .in0(N__4745),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8137),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_8_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_8_5_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_8_5_0  (
            .in0(N__5731),
            .in1(N__5325),
            .in2(_gnd_net_),
            .in3(N__5605),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_8_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_8_5_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_8_5_5  (
            .in0(N__5606),
            .in1(N__5334),
            .in2(_gnd_net_),
            .in3(N__5732),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_8_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_8_5_6 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_8_5_6  (
            .in0(N__4222),
            .in1(N__4180),
            .in2(N__3905),
            .in3(N__5089),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_5_7 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3902),
            .in3(N__9086),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9227),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_8_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_8_6_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_8_6_0  (
            .in0(N__4533),
            .in1(N__4558),
            .in2(N__5446),
            .in3(N__5406),
            .lcout(\U712_CHIP_RAM.N_272 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_6_2 .LUT_INIT=16'b0000001110101011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_6_2  (
            .in0(N__5442),
            .in1(N__4142),
            .in2(N__4073),
            .in3(N__8162),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9232),
            .ce(),
            .sr(N__9030));
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_8_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_8_6_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_8_6_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DBR_SYNC_0_LC_8_6_3  (
            .in0(N__4049),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(U712_REG_SM_DBR_SYNC_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9232),
            .ce(),
            .sr(N__9030));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_8_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_8_6_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_8_6_5  (
            .in0(N__4557),
            .in1(N__4532),
            .in2(_gnd_net_),
            .in3(N__5438),
            .lcout(\U712_CHIP_RAM.N_287 ),
            .ltout(\U712_CHIP_RAM.N_287_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRB433_1_LC_8_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRB433_1_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRB433_1_LC_8_6_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRB433_1_LC_8_6_6  (
            .in0(N__5614),
            .in1(N__4439),
            .in2(N__4028),
            .in3(N__5736),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVNIQ6_3_LC_8_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVNIQ6_3_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVNIQ6_3_LC_8_6_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVNIQ6_3_LC_8_6_7  (
            .in0(N__4025),
            .in1(N__7177),
            .in2(N__4019),
            .in3(N__5081),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DBR_SYNC_1_LC_8_7_1 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_8_7_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_8_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_1_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4537),
            .lcout(U712_REG_SM_DBR_SYNC_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9234),
            .ce(),
            .sr(N__9024));
    defparam \U712_CHIP_RAM.DBDIR_LC_8_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_8_7_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_8_7_2 .LUT_INIT=16'b1111000001110100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_8_7_2  (
            .in0(N__4489),
            .in1(N__7000),
            .in2(N__4614),
            .in3(N__6976),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9234),
            .ce(),
            .sr(N__9024));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_9_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__4011),
            .in2(_gnd_net_),
            .in3(N__3997),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_LC_8_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_8_10_1 .LUT_INIT=16'b1111101101010000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_8_10_1  (
            .in0(N__4832),
            .in1(N__4800),
            .in2(N__4157),
            .in3(N__4782),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9240),
            .ce(),
            .sr(N__9005));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_10_2 .LUT_INIT=16'b0101000001110011;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_8_10_2  (
            .in0(N__4091),
            .in1(N__4138),
            .in2(N__4432),
            .in3(N__4112),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9240),
            .ce(),
            .sr(N__9005));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_8_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_8_10_3 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_8_10_3  (
            .in0(N__4945),
            .in1(N__4366),
            .in2(_gnd_net_),
            .in3(N__6322),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9240),
            .ce(),
            .sr(N__9005));
    defparam \U712_REG_SM.DS_EN_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_8_10_5 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \U712_REG_SM.DS_EN_LC_8_10_5  (
            .in0(N__4284),
            .in1(N__4928),
            .in2(N__4955),
            .in3(N__4082),
            .lcout(\U712_REG_SM.DS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9240),
            .ce(),
            .sr(N__9005));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_10_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_10_6 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_8_10_6  (
            .in0(N__4424),
            .in1(N__4402),
            .in2(N__5018),
            .in3(N__6373),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9240),
            .ce(),
            .sr(N__9005));
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_8_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_8_10_7 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_GO_LC_8_10_7  (
            .in0(N__4401),
            .in1(N__4090),
            .in2(N__4373),
            .in3(N__4428),
            .lcout(\U712_REG_SM.REG_CYCLE_GOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9240),
            .ce(),
            .sr(N__9005));
    defparam \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_8_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_8_11_2 .LUT_INIT=16'b0000111100000001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_8_11_2  (
            .in0(N__6387),
            .in1(N__4678),
            .in2(N__6374),
            .in3(N__5014),
            .lcout(\U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1 ),
            .ltout(\U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_1_ess_RNO_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_1_ess_RNO_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REGENn_1_ess_RNO_LC_8_11_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_REG_SM.REGENn_1_ess_RNO_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4076),
            .in3(N__9081),
            .lcout(\U712_REG_SM.N_186_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_8_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_8_11_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_8_11_5  (
            .in0(N__4679),
            .in1(N__6371),
            .in2(_gnd_net_),
            .in3(N__6388),
            .lcout(\U712_REG_SM.N_342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDS_OUT_LC_8_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.LDS_OUT_LC_8_12_4 .LUT_INIT=16'b1100110010101111;
    LogicCell40 \U712_REG_SM.LDS_OUT_LC_8_12_4  (
            .in0(N__6203),
            .in1(N__4342),
            .in2(N__4387),
            .in3(N__4364),
            .lcout(\U712_REG_SM.LDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9244),
            .ce(),
            .sr(N__8994));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_8_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_8_12_5 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_8_12_5  (
            .in0(N__4363),
            .in1(N__4433),
            .in2(N__4694),
            .in3(N__4406),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9244),
            .ce(),
            .sr(N__8994));
    defparam \U712_REG_SM.UDS_OUT_LC_8_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.UDS_OUT_LC_8_12_6 .LUT_INIT=16'b1100110001011111;
    LogicCell40 \U712_REG_SM.UDS_OUT_LC_8_12_6  (
            .in0(N__6204),
            .in1(N__4303),
            .in2(N__4388),
            .in3(N__4365),
            .lcout(\U712_REG_SM.UDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9244),
            .ce(),
            .sr(N__8994));
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_13_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__4291),
            .in2(_gnd_net_),
            .in3(N__4343),
            .lcout(U712_REG_SM_un1_LDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_8_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_8_14_7 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_REG_SM.UDS_OUT_RNIUP9B_LC_8_14_7  (
            .in0(N__4307),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4292),
            .lcout(U712_REG_SM_un1_UDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_4_1 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_4_1  (
            .in0(N__5637),
            .in1(N__5339),
            .in2(N__5799),
            .in3(N__5160),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9214),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_9_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_9_4_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_9_4_3  (
            .in0(N__4221),
            .in1(N__4179),
            .in2(N__5095),
            .in3(N__4455),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_4_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_4_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_4_4  (
            .in0(N__9087),
            .in1(_gnd_net_),
            .in2(N__4247),
            .in3(N__4201),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9214),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_4_7 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_4_7  (
            .in0(N__4200),
            .in1(N__9088),
            .in2(N__4244),
            .in3(N__4235),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9214),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_5_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_5_0  (
            .in0(N__4234),
            .in1(N__4223),
            .in2(N__4202),
            .in3(N__4178),
            .lcout(\U712_CHIP_RAM.N_276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_5_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_5_1  (
            .in0(N__5798),
            .in1(N__5642),
            .in2(_gnd_net_),
            .in3(N__5161),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9223),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_5_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_5_2  (
            .in0(N__5261),
            .in1(N__5402),
            .in2(_gnd_net_),
            .in3(N__4469),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_5_3 .LUT_INIT=16'b0000000001100111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_5_3  (
            .in0(N__6962),
            .in1(N__5742),
            .in2(N__4463),
            .in3(N__5171),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9223),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_9_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_9_5_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__5323),
            .in2(_gnd_net_),
            .in3(N__5074),
            .lcout(\U712_CHIP_RAM.N_273 ),
            .ltout(\U712_CHIP_RAM.N_273_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINN5O1_LC_9_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINN5O1_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINN5O1_LC_9_5_5 .LUT_INIT=16'b0000111111000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINN5O1_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__5741),
            .in2(N__4460),
            .in3(N__7127),
            .lcout(\U712_CHIP_RAM.N_296_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_5_6  (
            .in0(N__5162),
            .in1(N__4456),
            .in2(_gnd_net_),
            .in3(N__5075),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9223),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICGJU_LC_9_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICGJU_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICGJU_LC_9_5_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICGJU_LC_9_5_7  (
            .in0(N__5324),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5391),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a2_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_9_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_9_6_0 .LUT_INIT=16'b0000000010000100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_9_6_0  (
            .in0(N__5616),
            .in1(N__7114),
            .in2(N__5781),
            .in3(N__5817),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_0_a2_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_9_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_9_6_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__7178),
            .in2(_gnd_net_),
            .in3(N__7708),
            .lcout(\U712_CHIP_RAM.N_347 ),
            .ltout(\U712_CHIP_RAM.N_347_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHBQU6_0_LC_9_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHBQU6_0_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHBQU6_0_LC_9_6_2 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIHBQU6_0_LC_9_6_2  (
            .in0(N__5737),
            .in1(N__7216),
            .in2(N__4514),
            .in3(N__5465),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_378_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8KLPE_0_LC_9_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8KLPE_0_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8KLPE_0_LC_9_6_3 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI8KLPE_0_LC_9_6_3  (
            .in0(N__5262),
            .in1(N__7709),
            .in2(N__4511),
            .in3(N__4508),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_9_6_4 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_9_6_4  (
            .in0(N__7179),
            .in1(_gnd_net_),
            .in2(N__5541),
            .in3(N__4502),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_9_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_9_6_5 .LUT_INIT=16'b0000101011111010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_LC_9_6_5  (
            .in0(N__5110),
            .in1(_gnd_net_),
            .in2(N__4496),
            .in3(N__6975),
            .lcout(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9228),
            .ce(),
            .sr(N__9025));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_9_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_9_6_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__5419),
            .in2(_gnd_net_),
            .in3(N__5109),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER50 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER50_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_9_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_9_6_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_9_6_7  (
            .in0(N__7113),
            .in1(N__5615),
            .in2(N__4493),
            .in3(N__5531),
            .lcout(\U712_CHIP_RAM.N_424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_3_LC_9_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_3_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_3_LC_9_7_0 .LUT_INIT=16'b0000100011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_3_LC_9_7_0  (
            .in0(N__5792),
            .in1(N__7129),
            .in2(N__5658),
            .in3(N__4657),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_7_1 .LUT_INIT=16'b1111100000101101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_7_1  (
            .in0(N__7128),
            .in1(N__5819),
            .in2(N__5657),
            .in3(N__5793),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_7_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_7_2  (
            .in0(N__5003),
            .in1(N__4490),
            .in2(_gnd_net_),
            .in3(N__5395),
            .lcout(\U712_CHIP_RAM.N_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_3_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_3_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_3_LC_9_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_sbtinv_3_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5492),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_9_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_9_7_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_9_7_4  (
            .in0(N__5263),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5196),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_7_6 .LUT_INIT=16'b0110100011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_7_6  (
            .in0(N__5794),
            .in1(N__7130),
            .in2(N__5659),
            .in3(N__4658),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_e_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_7_7 .LUT_INIT=16'b1111111000110010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_7_7  (
            .in0(N__5850),
            .in1(N__5493),
            .in2(N__4646),
            .in3(N__8717),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9233),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_3_LC_9_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_3_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_3_LC_9_8_0 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_3_LC_9_8_0  (
            .in0(N__5851),
            .in1(N__5660),
            .in2(N__4643),
            .in3(N__5510),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9235),
            .ce(N__4634),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_9_9_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_9_9_0 .LUT_INIT=16'b1100110000001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_9_9_0  (
            .in0(N__4783),
            .in1(N__6350),
            .in2(N__4807),
            .in3(N__4834),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9236),
            .ce(),
            .sr(N__9006));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_9_9_4 .LUT_INIT=16'b0001000101010000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_9_9_4  (
            .in0(N__4667),
            .in1(N__6349),
            .in2(N__4922),
            .in3(N__4833),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9236),
            .ce(),
            .sr(N__9006));
    defparam \U712_BUFFERS.DRDDIR_i_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_LC_9_10_0 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_LC_9_10_0  (
            .in0(N__4737),
            .in1(N__5982),
            .in2(N__4621),
            .in3(N__4999),
            .lcout(N_188),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_9_10_1 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_9_10_1  (
            .in0(N__6337),
            .in1(N__6577),
            .in2(_gnd_net_),
            .in3(N__6532),
            .lcout(\U712_REG_SM.N_288 ),
            .ltout(\U712_REG_SM.N_288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_10_2 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__4565),
            .in2(N__4544),
            .in3(N__4541),
            .lcout(\U712_REG_SM.N_301 ),
            .ltout(\U712_REG_SM.N_301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_9_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_10_3 .LUT_INIT=16'b1101110110001100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_9_10_3  (
            .in0(N__4835),
            .in1(N__4756),
            .in2(N__4811),
            .in3(N__4736),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9237),
            .ce(),
            .sr(N__8998));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_10_5 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_9_10_5  (
            .in0(N__4766),
            .in1(N__4784),
            .in2(N__4808),
            .in3(N__4757),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9237),
            .ce(),
            .sr(N__8998));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_10_6 .LUT_INIT=16'b0010111000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_9_10_6  (
            .in0(N__4755),
            .in1(N__4946),
            .in2(N__6323),
            .in3(N__4765),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9237),
            .ce(),
            .sr(N__8998));
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_9_10_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a2_LC_9_10_7  (
            .in0(N__5983),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4738),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_9_11_0 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_9_11_0  (
            .in0(N__6575),
            .in1(_gnd_net_),
            .in2(N__6531),
            .in3(N__4690),
            .lcout(\U712_REG_SM.N_341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_9_11_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_9_11_1  (
            .in0(N__6552),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6125),
            .lcout(\U712_REG_SM.N_294 ),
            .ltout(\U712_REG_SM.N_294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_9_11_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_9_11_2  (
            .in0(N__6405),
            .in1(N__6606),
            .in2(N__4670),
            .in3(N__6640),
            .lcout(\U712_REG_SM.N_373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_9_11_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__6574),
            .in2(_gnd_net_),
            .in3(N__6519),
            .lcout(\U712_REG_SM.N_292 ),
            .ltout(\U712_REG_SM.N_292_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_9_11_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_9_11_4  (
            .in0(N__4920),
            .in1(N__6605),
            .in2(N__5021),
            .in3(N__6639),
            .lcout(\U712_REG_SM.N_507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_9_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_9_11_5 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_9_11_5  (
            .in0(N__6553),
            .in1(N__6644),
            .in2(_gnd_net_),
            .in3(N__4998),
            .lcout(\U712_REG_SM.N_104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_9_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_9_11_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__6604),
            .in2(_gnd_net_),
            .in3(N__6638),
            .lcout(\U712_REG_SM.N_298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_9_11_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_1_LC_9_11_7  (
            .in0(N__4944),
            .in1(N__6576),
            .in2(N__6341),
            .in3(N__6523),
            .lcout(\U712_REG_SM.N_372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_1_ess_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_1_ess_LC_9_12_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_1_ess_LC_9_12_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_REG_SM.REGENn_1_ess_LC_9_12_2  (
            .in0(N__4921),
            .in1(N__6645),
            .in2(N__6410),
            .in3(N__6607),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9242),
            .ce(N__4856),
            .sr(N__8992));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_10_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_10_4_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_10_4_0 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_10_4_0  (
            .in0(N__5259),
            .in1(N__6955),
            .in2(N__4844),
            .in3(N__5204),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_10_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_10_4_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_10_4_1 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_10_4_1  (
            .in0(N__8063),
            .in1(N__6963),
            .in2(N__4850),
            .in3(N__5408),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9210),
            .ce(),
            .sr(N__9031));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_2_LC_10_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_2_LC_10_4_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_2_LC_10_4_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNO_2_LC_10_4_2  (
            .in0(N__5613),
            .in1(N__5746),
            .in2(N__5353),
            .in3(N__8062),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_1_LC_10_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_1_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_1_LC_10_4_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNO_1_LC_10_4_3  (
            .in0(N__5085),
            .in1(N__5257),
            .in2(N__4847),
            .in3(N__7189),
            .lcout(\U712_CHIP_RAM.N_393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJV8G1_2_LC_10_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJV8G1_2_LC_10_4_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJV8G1_2_LC_10_4_4 .LUT_INIT=16'b0001100000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIJV8G1_2_LC_10_4_4  (
            .in0(N__5611),
            .in1(N__5327),
            .in2(N__5091),
            .in3(N__8061),
            .lcout(\U712_CHIP_RAM.N_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6IFV8_0_LC_10_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6IFV8_0_LC_10_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6IFV8_0_LC_10_4_5 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6IFV8_0_LC_10_4_5  (
            .in0(N__7181),
            .in1(N__9084),
            .in2(N__5783),
            .in3(N__5453),
            .lcout(\U712_CHIP_RAM.N_310 ),
            .ltout(\U712_CHIP_RAM.N_310_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDCLTE_0_LC_10_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDCLTE_0_LC_10_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDCLTE_0_LC_10_4_6 .LUT_INIT=16'b1111000011111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIDCLTE_0_LC_10_4_6  (
            .in0(N__5258),
            .in1(N__5203),
            .in2(N__5165),
            .in3(N__6954),
            .lcout(\U712_CHIP_RAM.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_10_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_10_4_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_10_4_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_10_4_7  (
            .in0(N__7180),
            .in1(N__5612),
            .in2(N__5782),
            .in3(N__5535),
            .lcout(\U712_CHIP_RAM.N_293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_0 .LUT_INIT=16'b1111101111111110;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_5_0  (
            .in0(N__5247),
            .in1(N__5734),
            .in2(N__5638),
            .in3(N__5338),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_3_0_a2_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_5_1 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_5_1  (
            .in0(_gnd_net_),
            .in1(N__7193),
            .in2(N__5147),
            .in3(N__5077),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_179_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_10_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_10_5_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_10_5_2 .LUT_INIT=16'b1010110010101111;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_10_5_2  (
            .in0(N__5122),
            .in1(N__6914),
            .in2(N__5144),
            .in3(N__5735),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9215),
            .ce(),
            .sr(N__9026));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_10_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_10_5_3 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_10_5_3  (
            .in0(N__7097),
            .in1(N__5420),
            .in2(_gnd_net_),
            .in3(N__5111),
            .lcout(\U712_CHIP_RAM.N_284 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_5_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_5_5  (
            .in0(_gnd_net_),
            .in1(N__5607),
            .in2(_gnd_net_),
            .in3(N__5076),
            .lcout(\U712_CHIP_RAM.N_438 ),
            .ltout(\U712_CHIP_RAM.N_438_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILE372_2_LC_10_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILE372_2_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILE372_2_LC_10_5_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNILE372_2_LC_10_5_6  (
            .in0(N__5326),
            .in1(N__7098),
            .in2(N__5024),
            .in3(N__5733),
            .lcout(\U712_CHIP_RAM.N_425 ),
            .ltout(\U712_CHIP_RAM.N_425_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI94U46_2_LC_10_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI94U46_2_LC_10_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI94U46_2_LC_10_5_7 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI94U46_2_LC_10_5_7  (
            .in0(N__5474),
            .in1(N__5246),
            .in2(N__5468),
            .in3(N__5464),
            .lcout(\U712_CHIP_RAM.N_302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_6_0 .LUT_INIT=16'b0101110100001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_6_0  (
            .in0(N__5958),
            .in1(N__8786),
            .in2(N__8813),
            .in3(N__5401),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9224),
            .ce(),
            .sr(N__9020));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNO_0_LC_10_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNO_0_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNO_0_LC_10_6_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNO_0_LC_10_6_1  (
            .in0(N__5397),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5447),
            .lcout(),
            .ltout(\U712_CHIP_RAM.REFRESH_CYCLE_START_2_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_10_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_10_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_10_6_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_10_6_2  (
            .in0(N__5959),
            .in1(N__6875),
            .in2(N__5423),
            .in3(N__8132),
            .lcout(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9224),
            .ce(),
            .sr(N__9020));
    defparam \U712_CHIP_RAM.DMA_CYCLE_1_LC_10_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_1_LC_10_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_1_LC_10_6_3 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_1_LC_10_6_3  (
            .in0(N__6965),
            .in1(N__5957),
            .in2(N__5407),
            .in3(N__5177),
            .lcout(RAMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9224),
            .ce(),
            .sr(N__9020));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_10_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_10_6_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_10_6_4  (
            .in0(_gnd_net_),
            .in1(N__7916),
            .in2(_gnd_net_),
            .in3(N__5396),
            .lcout(\U712_CHIP_RAM.DBENn_7_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_10_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_10_6_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_10_6_5  (
            .in0(N__5787),
            .in1(N__7188),
            .in2(N__5354),
            .in3(N__5273),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIB6KL9_2_LC_10_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIB6KL9_2_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIB6KL9_2_LC_10_6_6 .LUT_INIT=16'b0101000101010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIB6KL9_2_LC_10_6_6  (
            .in0(N__5260),
            .in1(N__6964),
            .in2(N__5207),
            .in3(N__5202),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_10_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_10_6_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_10_6_7 .LUT_INIT=16'b1010110011111100;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_10_6_7  (
            .in0(N__5788),
            .in1(N__6014),
            .in2(N__5864),
            .in3(N__5861),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9224),
            .ce(),
            .sr(N__9020));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_7_0 .LUT_INIT=16'b1111111011110110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_7_0  (
            .in0(N__5790),
            .in1(N__5542),
            .in2(N__5855),
            .in3(N__7112),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_i_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_7_1 .LUT_INIT=16'b1010101011111100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_7_1  (
            .in0(N__8480),
            .in1(N__5828),
            .in2(N__5822),
            .in3(N__5494),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9229),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVS9V_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVS9V_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVS9V_LC_10_7_2 .LUT_INIT=16'b0010001001100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVS9V_LC_10_7_2  (
            .in0(N__5789),
            .in1(N__7108),
            .in2(_gnd_net_),
            .in3(N__5818),
            .lcout(\U712_CHIP_RAM.N_305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_7_3 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_7_3  (
            .in0(N__6913),
            .in1(N__5791),
            .in2(N__7126),
            .in3(N__5646),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_7_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_7_4  (
            .in0(N__7205),
            .in1(N__5543),
            .in2(N__5513),
            .in3(N__7702),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_i_0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_7_5 .LUT_INIT=16'b1010101011111100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_7_5  (
            .in0(N__8569),
            .in1(N__5509),
            .in2(N__5498),
            .in3(N__5495),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9229),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNITDMK_3_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNITDMK_3_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNITDMK_3_LC_10_7_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNITDMK_3_LC_10_7_6  (
            .in0(N__8718),
            .in1(N__8568),
            .in2(N__8470),
            .in3(N__7043),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(\U712_CHIP_RAM.REFRESH_RST_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI9T531_3_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI9T531_3_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI9T531_3_LC_10_7_7 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI9T531_3_LC_10_7_7  (
            .in0(N__8696),
            .in1(N__8471),
            .in2(N__5477),
            .in3(N__7044),
            .lcout(\U712_CHIP_RAM.un1_CMA31_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_8_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_10_8_1  (
            .in0(N__5972),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6024),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0 ),
            .ltout(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_192_i_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_192_i_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_192_i_LC_10_8_2 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \U712_BYTE_ENABLE.N_192_i_LC_10_8_2  (
            .in0(N__8858),
            .in1(N__5914),
            .in2(N__6113),
            .in3(N__5870),
            .lcout(N_192_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_194_i_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_194_i_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_194_i_LC_10_8_3 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \U712_BYTE_ENABLE.N_194_i_LC_10_8_3  (
            .in0(N__5915),
            .in1(N__6089),
            .in2(N__8900),
            .in3(N__6275),
            .lcout(N_194_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_10_9_1 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_10_9_1  (
            .in0(N__6065),
            .in1(N__6304),
            .in2(_gnd_net_),
            .in3(N__8150),
            .lcout(\U712_BYTE_ENABLE.N_404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_0_LC_10_9_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_0_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_0_LC_10_9_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_0_LC_10_9_2  (
            .in0(N__6025),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5973),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0 ),
            .ltout(\U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_196_i_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_196_i_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_196_i_LC_10_9_3 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_196_i_LC_10_9_3  (
            .in0(N__5912),
            .in1(N__6179),
            .in2(N__5936),
            .in3(N__8853),
            .lcout(N_196_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_LC_10_9_4 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_LC_10_9_4  (
            .in0(N__8148),
            .in1(N__6265),
            .in2(N__6305),
            .in3(N__6232),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_411_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_198_i_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_198_i_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_198_i_LC_10_9_5 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_198_i_LC_10_9_5  (
            .in0(N__5913),
            .in1(N__5897),
            .in2(N__5891),
            .in3(N__8893),
            .lcout(N_198_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_0_LC_10_9_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_0_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_0_LC_10_9_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_0_LC_10_9_6  (
            .in0(N__8149),
            .in1(N__6233),
            .in2(_gnd_net_),
            .in3(N__6266),
            .lcout(\U712_BYTE_ENABLE.N_405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_10_10_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_10_10_0  (
            .in0(N__6406),
            .in1(N__6389),
            .in2(_gnd_net_),
            .in3(N__6372),
            .lcout(\U712_REG_SM.N_309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_10_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_10_1  (
            .in0(N__6124),
            .in1(N__6603),
            .in2(N__6647),
            .in3(N__6551),
            .lcout(\U712_REG_SM.N_282 ),
            .ltout(\U712_REG_SM.N_282_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_10_2 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__6578),
            .in2(N__6326),
            .in3(N__6533),
            .lcout(\U712_REG_SM.N_306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_10_10_6 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_10_10_6  (
            .in0(N__6300),
            .in1(N__6264),
            .in2(N__8168),
            .in3(N__6231),
            .lcout(\U712_BYTE_ENABLE.N_407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_10_10_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_10_10_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_10_10_7  (
            .in0(N__6263),
            .in1(N__6230),
            .in2(_gnd_net_),
            .in3(N__8151),
            .lcout(\U712_BYTE_ENABLE.N_409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_0_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_10_11_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_10_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6173),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9238),
            .ce(),
            .sr(N__8993));
    defparam \U712_REG_SM.C3_SYNC_0_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_10_11_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_10_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6140),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9238),
            .ce(),
            .sr(N__8993));
    defparam \U712_REG_SM.C1_SYNC_2_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_2_LC_10_11_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_2_LC_10_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_2_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6608),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9238),
            .ce(),
            .sr(N__8993));
    defparam \U712_REG_SM.C1_SYNC_1_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_10_11_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_10_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6646),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9238),
            .ce(),
            .sr(N__8993));
    defparam \U712_REG_SM.C3_SYNC_2_LC_10_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_2_LC_10_11_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_2_LC_10_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_2_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6530),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9238),
            .ce(),
            .sr(N__8993));
    defparam \U712_REG_SM.C3_SYNC_1_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_10_12_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_10_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6554),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9241),
            .ce(),
            .sr(N__8991));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_2_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_2_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_2_1 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_11_2_1  (
            .in0(N__6416),
            .in1(_gnd_net_),
            .in2(N__8639),
            .in3(N__8759),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9203),
            .ce(N__7964),
            .sr(N__9036));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_11_2_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_11_2_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_11_2_2 .LUT_INIT=16'b1111000011010001;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_11_2_2  (
            .in0(N__8518),
            .in1(N__8620),
            .in2(N__6659),
            .in3(N__8758),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9203),
            .ce(N__7964),
            .sr(N__9036));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_11_2_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_11_2_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_11_2_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_11_2_3  (
            .in0(N__8757),
            .in1(N__8519),
            .in2(N__8638),
            .in3(N__7061),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9203),
            .ce(N__7964),
            .sr(N__9036));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_3_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_3_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_3_2  (
            .in0(N__7325),
            .in1(N__8092),
            .in2(N__7421),
            .in3(N__8520),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_3_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_3_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_3_3  (
            .in0(N__8093),
            .in1(N__6458),
            .in2(N__6440),
            .in3(N__6437),
            .lcout(\U712_CHIP_RAM.N_317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_4_1 .LUT_INIT=16'b0000001111110101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_4_1  (
            .in0(N__7235),
            .in1(N__7592),
            .in2(N__8146),
            .in3(N__8503),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_4_2 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_4_2  (
            .in0(N__8106),
            .in1(N__6857),
            .in2(N__6839),
            .in3(N__6836),
            .lcout(\U712_CHIP_RAM.N_320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_11_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_11_4_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_11_4_4  (
            .in0(N__7622),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9207),
            .ce(N__7837),
            .sr(N__9027));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_4_5 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_4_5  (
            .in0(N__7241),
            .in1(N__8502),
            .in2(N__8147),
            .in3(N__7538),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_4_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_11_4_6  (
            .in0(N__8107),
            .in1(N__6809),
            .in2(N__6791),
            .in3(N__6788),
            .lcout(\U712_CHIP_RAM.N_321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_5_0 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_5_0  (
            .in0(N__8496),
            .in1(N__7229),
            .in2(N__8133),
            .in3(N__9257),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_5_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_5_1  (
            .in0(N__6767),
            .in1(N__6746),
            .in2(N__6725),
            .in3(N__8080),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_315_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_11_5_2 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_11_5_2  (
            .in0(N__8753),
            .in1(_gnd_net_),
            .in2(N__6722),
            .in3(N__8619),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9211),
            .ce(N__7951),
            .sr(N__9021));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_5_3 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_5_3  (
            .in0(N__7223),
            .in1(N__8076),
            .in2(N__8514),
            .in3(N__7499),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_5_4 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_5_4  (
            .in0(N__6701),
            .in1(N__6680),
            .in2(N__6662),
            .in3(N__8099),
            .lcout(\U712_CHIP_RAM.N_316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_11_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_11_6_0 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_11_6_0  (
            .in0(N__7125),
            .in1(N__7217),
            .in2(_gnd_net_),
            .in3(N__7204),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9216),
            .ce(),
            .sr(N__9013));
    defparam \U712_CHIP_RAM.CRCSn_LC_11_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_11_6_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_11_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7060),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9216),
            .ce(),
            .sr(N__9013));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_11_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_11_7_1 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_11_7_1  (
            .in0(N__6912),
            .in1(N__7004),
            .in2(N__6989),
            .in3(N__6977),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9225),
            .ce(),
            .sr(N__9007));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIV62J1_3_LC_11_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIV62J1_3_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIV62J1_3_LC_11_7_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIV62J1_3_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__9082),
            .in2(_gnd_net_),
            .in3(N__6893),
            .lcout(\U712_CHIP_RAM.un1_CMA31_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_0_LC_11_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_0_LC_11_8_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_0_LC_11_8_0  (
            .in0(N__7363),
            .in1(N__7743),
            .in2(N__7346),
            .in3(N__7795),
            .lcout(),
            .ltout(\U712_CHIP_RAM.REFRESH_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_0_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_0_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_0_LC_11_8_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_0_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__7393),
            .in2(N__6887),
            .in3(N__6865),
            .lcout(\U712_CHIP_RAM.REFRESHZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9230),
            .ce(),
            .sr(N__8999));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_1_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_1_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_1_LC_11_8_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_1_LC_11_8_3  (
            .in0(N__7794),
            .in1(N__7341),
            .in2(_gnd_net_),
            .in3(N__7362),
            .lcout(),
            .ltout(\U712_CHIP_RAM.REFRESH9lt7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_1_LC_11_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_1_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_1_LC_11_8_4 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_1_LC_11_8_4  (
            .in0(N__6866),
            .in1(N__6884),
            .in2(N__6878),
            .in3(N__7744),
            .lcout(\U712_CHIP_RAM.REFRESHZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9230),
            .ce(),
            .sr(N__8999));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_RNILI9L_5_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_RNILI9L_5_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_RNILI9L_5_LC_11_9_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_RNILI9L_5_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__7762),
            .in2(_gnd_net_),
            .in3(N__7777),
            .lcout(\U712_CHIP_RAM.REFRESH9lto7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_3_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7489),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9202),
            .ce(N__7833),
            .sr(N__9023));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_4_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_4_4 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_12_4_4  (
            .in0(N__8627),
            .in1(_gnd_net_),
            .in2(N__8767),
            .in3(N__7319),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9205),
            .ce(N__7965),
            .sr(N__9018));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_4_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_4_6 .LUT_INIT=16'b1111101100000001;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_12_4_6  (
            .in0(N__8760),
            .in1(N__8506),
            .in2(N__8640),
            .in3(N__7292),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9205),
            .ce(N__7965),
            .sr(N__9018));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_4_7 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_12_4_7  (
            .in0(N__7271),
            .in1(N__8204),
            .in2(N__7574),
            .in3(N__8136),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9205),
            .ce(N__7965),
            .sr(N__9018));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_12_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_12_5_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_12_5_2  (
            .in0(N__8309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9206),
            .ce(N__7832),
            .sr(N__9012));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_12_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_12_5_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_12_5_4  (
            .in0(N__7564),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9206),
            .ce(N__7832),
            .sr(N__9012));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_5_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_5_5  (
            .in0(N__7529),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9206),
            .ce(N__7832),
            .sr(N__9012));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7453),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9206),
            .ce(N__7832),
            .sr(N__9012));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_6_0  (
            .in0(N__7525),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9209),
            .ce(N__9116),
            .sr(N__9003));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_6_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_12_6_3  (
            .in0(N__7493),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9209),
            .ce(N__9116),
            .sr(N__9003));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7457),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9209),
            .ce(N__9116),
            .sr(N__9003));
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_12_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_12_7_0 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_12_7_0  (
            .in0(N__9080),
            .in1(N__8779),
            .in2(_gnd_net_),
            .in3(N__8802),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_7_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_7_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_7_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_8_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_8_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(N__7382),
            .in2(_gnd_net_),
            .in3(N__7376),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(bfn_12_8_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__7730),
            .ce(),
            .sr(N__7721));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_8_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_8_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__7373),
            .in2(_gnd_net_),
            .in3(N__7367),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__7730),
            .ce(),
            .sr(N__7721));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_8_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_8_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(N__7364),
            .in2(_gnd_net_),
            .in3(N__7349),
            .lcout(\U712_CHIP_RAM.REFRESH9lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__7730),
            .ce(),
            .sr(N__7721));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_8_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_8_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(N__7345),
            .in2(_gnd_net_),
            .in3(N__7328),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__7730),
            .ce(),
            .sr(N__7721));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_8_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_8_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(N__7796),
            .in2(_gnd_net_),
            .in3(N__7781),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__7730),
            .ce(),
            .sr(N__7721));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_8_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_8_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(N__7778),
            .in2(_gnd_net_),
            .in3(N__7766),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__7730),
            .ce(),
            .sr(N__7721));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_8_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_8_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_8_6  (
            .in0(_gnd_net_),
            .in1(N__7763),
            .in2(_gnd_net_),
            .in3(N__7751),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__7730),
            .ce(),
            .sr(N__7721));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_8_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_8_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__7745),
            .in2(_gnd_net_),
            .in3(N__7748),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7730),
            .ce(),
            .sr(N__7721));
    defparam RESETn_ibuf_RNIM9SF_LC_12_14_5.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_14_5.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_14_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7685),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_4_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7618),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9208),
            .ce(N__9108),
            .sr(N__9028));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_4_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7907),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9208),
            .ce(N__9108),
            .sr(N__9028));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_4_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7871),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9208),
            .ce(N__9108),
            .sr(N__9028));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_4_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7565),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9208),
            .ce(N__9108),
            .sr(N__9028));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_5_0 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_5_0  (
            .in0(N__7844),
            .in1(N__8505),
            .in2(N__8173),
            .in3(N__8273),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_5_1 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_5_1  (
            .in0(N__8166),
            .in1(N__8267),
            .in2(N__8249),
            .in3(N__8246),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_322_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_5_2 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_13_5_2  (
            .in0(N__8615),
            .in1(_gnd_net_),
            .in2(N__8228),
            .in3(N__8754),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9212),
            .ce(N__7966),
            .sr(N__9022));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_5_5 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_5_5  (
            .in0(N__8504),
            .in1(N__8749),
            .in2(_gnd_net_),
            .in3(N__8614),
            .lcout(\U712_CHIP_RAM.CMA_5_i_0_8 ),
            .ltout(\U712_CHIP_RAM.CMA_5_i_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_5_6 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_13_5_6  (
            .in0(N__8198),
            .in1(N__8377),
            .in2(N__8177),
            .in3(N__8167),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9212),
            .ce(N__7966),
            .sr(N__9022));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_13_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_13_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_13_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9295),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9217),
            .ce(N__7838),
            .sr(N__9014));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_13_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_13_6_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_13_6_4  (
            .in0(N__7906),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9217),
            .ce(N__7838),
            .sr(N__9014));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_13_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_13_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7867),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9217),
            .ce(N__7838),
            .sr(N__9014));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_13_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_13_7_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_13_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__8892),
            .in2(_gnd_net_),
            .in3(N__8857),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9226),
            .ce(),
            .sr(N__9008));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_7_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8806),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9226),
            .ce(),
            .sr(N__9008));
    defparam \U712_CHIP_RAM.RASn_LC_14_1_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_14_1_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_14_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_14_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8768),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9204),
            .ce(),
            .sr(N__9050));
    defparam \U712_CHIP_RAM.WEn_LC_14_1_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_14_1_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_14_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_14_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8642),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9204),
            .ce(),
            .sr(N__9050));
    defparam \U712_CHIP_RAM.CASn_LC_14_1_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_14_1_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_14_1_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_14_1_7  (
            .in0(N__8522),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9204),
            .ce(),
            .sr(N__9050));
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_14_3_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_14_3_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_14_3_3 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_14_3_3  (
            .in0(N__9085),
            .in1(N__8326),
            .in2(_gnd_net_),
            .in3(N__8315),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_14_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_14_4_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_14_4_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_14_4_0  (
            .in0(N__8378),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8342),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9213),
            .ce(),
            .sr(N__9032));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_14_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_14_4_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_14_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_14_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8327),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9213),
            .ce(),
            .sr(N__9032));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_5_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_5_0  (
            .in0(N__8308),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9218),
            .ce(N__9112),
            .sr(N__9029));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9296),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9218),
            .ce(N__9112),
            .sr(N__9029));
endmodule // U712_TOP

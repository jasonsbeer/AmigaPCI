// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 12 2025 17:26:36

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U400_TOP" view "INTERFACE"

module U400_TOP (
    SIZ,
    MA,
    A,
    LBENn,
    CS0n,
    UUBEn,
    TAn,
    CLK40,
    RnW,
    BANK1,
    UMBEn,
    WEn,
    LLBEn,
    TSn,
    LMBEn,
    RASn,
    CS1n,
    RESETn,
    CLK_EN,
    CASn,
    BANK0);

    input [1:0] SIZ;
    output [12:0] MA;
    input [31:0] A;
    output LBENn;
    output CS0n;
    output UUBEn;
    output TAn;
    input CLK40;
    input RnW;
    output BANK1;
    output UMBEn;
    output WEn;
    output LLBEn;
    input TSn;
    output LMBEn;
    output RASn;
    output CS1n;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;

    wire N__7469;
    wire N__7468;
    wire N__7467;
    wire N__7460;
    wire N__7459;
    wire N__7458;
    wire N__7451;
    wire N__7450;
    wire N__7449;
    wire N__7442;
    wire N__7441;
    wire N__7440;
    wire N__7433;
    wire N__7432;
    wire N__7431;
    wire N__7424;
    wire N__7423;
    wire N__7422;
    wire N__7415;
    wire N__7414;
    wire N__7413;
    wire N__7406;
    wire N__7405;
    wire N__7404;
    wire N__7397;
    wire N__7396;
    wire N__7395;
    wire N__7388;
    wire N__7387;
    wire N__7386;
    wire N__7379;
    wire N__7378;
    wire N__7377;
    wire N__7370;
    wire N__7369;
    wire N__7368;
    wire N__7361;
    wire N__7360;
    wire N__7359;
    wire N__7352;
    wire N__7351;
    wire N__7350;
    wire N__7343;
    wire N__7342;
    wire N__7341;
    wire N__7334;
    wire N__7333;
    wire N__7332;
    wire N__7325;
    wire N__7324;
    wire N__7323;
    wire N__7316;
    wire N__7315;
    wire N__7314;
    wire N__7307;
    wire N__7306;
    wire N__7305;
    wire N__7298;
    wire N__7297;
    wire N__7296;
    wire N__7289;
    wire N__7288;
    wire N__7287;
    wire N__7280;
    wire N__7279;
    wire N__7278;
    wire N__7271;
    wire N__7270;
    wire N__7269;
    wire N__7262;
    wire N__7261;
    wire N__7260;
    wire N__7253;
    wire N__7252;
    wire N__7251;
    wire N__7244;
    wire N__7243;
    wire N__7242;
    wire N__7235;
    wire N__7234;
    wire N__7233;
    wire N__7226;
    wire N__7225;
    wire N__7224;
    wire N__7217;
    wire N__7216;
    wire N__7215;
    wire N__7208;
    wire N__7207;
    wire N__7206;
    wire N__7199;
    wire N__7198;
    wire N__7197;
    wire N__7190;
    wire N__7189;
    wire N__7188;
    wire N__7181;
    wire N__7180;
    wire N__7179;
    wire N__7172;
    wire N__7171;
    wire N__7170;
    wire N__7163;
    wire N__7162;
    wire N__7161;
    wire N__7154;
    wire N__7153;
    wire N__7152;
    wire N__7145;
    wire N__7144;
    wire N__7143;
    wire N__7136;
    wire N__7135;
    wire N__7134;
    wire N__7127;
    wire N__7126;
    wire N__7125;
    wire N__7118;
    wire N__7117;
    wire N__7116;
    wire N__7109;
    wire N__7108;
    wire N__7107;
    wire N__7100;
    wire N__7099;
    wire N__7098;
    wire N__7091;
    wire N__7090;
    wire N__7089;
    wire N__7082;
    wire N__7081;
    wire N__7080;
    wire N__7073;
    wire N__7072;
    wire N__7071;
    wire N__7064;
    wire N__7063;
    wire N__7062;
    wire N__7055;
    wire N__7054;
    wire N__7053;
    wire N__7046;
    wire N__7045;
    wire N__7044;
    wire N__7037;
    wire N__7036;
    wire N__7035;
    wire N__7028;
    wire N__7027;
    wire N__7026;
    wire N__7019;
    wire N__7018;
    wire N__7017;
    wire N__7010;
    wire N__7009;
    wire N__7008;
    wire N__7001;
    wire N__7000;
    wire N__6999;
    wire N__6992;
    wire N__6991;
    wire N__6990;
    wire N__6983;
    wire N__6982;
    wire N__6981;
    wire N__6974;
    wire N__6973;
    wire N__6972;
    wire N__6965;
    wire N__6964;
    wire N__6963;
    wire N__6956;
    wire N__6955;
    wire N__6954;
    wire N__6947;
    wire N__6946;
    wire N__6945;
    wire N__6938;
    wire N__6937;
    wire N__6936;
    wire N__6929;
    wire N__6928;
    wire N__6927;
    wire N__6920;
    wire N__6919;
    wire N__6918;
    wire N__6911;
    wire N__6910;
    wire N__6909;
    wire N__6902;
    wire N__6901;
    wire N__6900;
    wire N__6893;
    wire N__6892;
    wire N__6891;
    wire N__6874;
    wire N__6871;
    wire N__6868;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6858;
    wire N__6853;
    wire N__6852;
    wire N__6851;
    wire N__6850;
    wire N__6849;
    wire N__6846;
    wire N__6843;
    wire N__6836;
    wire N__6835;
    wire N__6834;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6817;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6801;
    wire N__6800;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6790;
    wire N__6787;
    wire N__6784;
    wire N__6781;
    wire N__6778;
    wire N__6777;
    wire N__6776;
    wire N__6767;
    wire N__6764;
    wire N__6761;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6747;
    wire N__6746;
    wire N__6743;
    wire N__6742;
    wire N__6741;
    wire N__6740;
    wire N__6739;
    wire N__6738;
    wire N__6737;
    wire N__6736;
    wire N__6735;
    wire N__6734;
    wire N__6733;
    wire N__6732;
    wire N__6731;
    wire N__6730;
    wire N__6697;
    wire N__6694;
    wire N__6691;
    wire N__6688;
    wire N__6687;
    wire N__6686;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6676;
    wire N__6673;
    wire N__6670;
    wire N__6667;
    wire N__6664;
    wire N__6661;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6640;
    wire N__6639;
    wire N__6636;
    wire N__6635;
    wire N__6632;
    wire N__6627;
    wire N__6626;
    wire N__6625;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6613;
    wire N__6612;
    wire N__6611;
    wire N__6610;
    wire N__6609;
    wire N__6608;
    wire N__6607;
    wire N__6606;
    wire N__6605;
    wire N__6604;
    wire N__6603;
    wire N__6602;
    wire N__6599;
    wire N__6598;
    wire N__6591;
    wire N__6588;
    wire N__6585;
    wire N__6582;
    wire N__6581;
    wire N__6580;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6562;
    wire N__6557;
    wire N__6556;
    wire N__6555;
    wire N__6552;
    wire N__6547;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6530;
    wire N__6523;
    wire N__6520;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6505;
    wire N__6500;
    wire N__6493;
    wire N__6490;
    wire N__6485;
    wire N__6480;
    wire N__6477;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6461;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6438;
    wire N__6435;
    wire N__6432;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6408;
    wire N__6407;
    wire N__6404;
    wire N__6403;
    wire N__6402;
    wire N__6401;
    wire N__6396;
    wire N__6391;
    wire N__6390;
    wire N__6389;
    wire N__6388;
    wire N__6383;
    wire N__6380;
    wire N__6377;
    wire N__6372;
    wire N__6371;
    wire N__6368;
    wire N__6367;
    wire N__6358;
    wire N__6357;
    wire N__6354;
    wire N__6351;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6334;
    wire N__6331;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6306;
    wire N__6305;
    wire N__6304;
    wire N__6299;
    wire N__6298;
    wire N__6297;
    wire N__6292;
    wire N__6291;
    wire N__6290;
    wire N__6289;
    wire N__6288;
    wire N__6285;
    wire N__6280;
    wire N__6277;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6257;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6249;
    wire N__6246;
    wire N__6243;
    wire N__6238;
    wire N__6235;
    wire N__6232;
    wire N__6223;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6193;
    wire N__6190;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6175;
    wire N__6172;
    wire N__6169;
    wire N__6166;
    wire N__6163;
    wire N__6160;
    wire N__6157;
    wire N__6154;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6124;
    wire N__6121;
    wire N__6118;
    wire N__6115;
    wire N__6112;
    wire N__6109;
    wire N__6106;
    wire N__6103;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6037;
    wire N__6036;
    wire N__6035;
    wire N__6034;
    wire N__6033;
    wire N__6032;
    wire N__6031;
    wire N__6028;
    wire N__6027;
    wire N__6026;
    wire N__6025;
    wire N__6024;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6012;
    wire N__6007;
    wire N__6006;
    wire N__6001;
    wire N__5996;
    wire N__5995;
    wire N__5994;
    wire N__5989;
    wire N__5980;
    wire N__5979;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5947;
    wire N__5942;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5928;
    wire N__5925;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5907;
    wire N__5902;
    wire N__5893;
    wire N__5892;
    wire N__5889;
    wire N__5888;
    wire N__5887;
    wire N__5886;
    wire N__5883;
    wire N__5880;
    wire N__5875;
    wire N__5872;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5856;
    wire N__5853;
    wire N__5852;
    wire N__5851;
    wire N__5848;
    wire N__5847;
    wire N__5846;
    wire N__5843;
    wire N__5838;
    wire N__5835;
    wire N__5830;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5809;
    wire N__5808;
    wire N__5807;
    wire N__5806;
    wire N__5805;
    wire N__5804;
    wire N__5803;
    wire N__5802;
    wire N__5801;
    wire N__5800;
    wire N__5797;
    wire N__5792;
    wire N__5789;
    wire N__5788;
    wire N__5787;
    wire N__5786;
    wire N__5785;
    wire N__5784;
    wire N__5783;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5768;
    wire N__5765;
    wire N__5758;
    wire N__5755;
    wire N__5752;
    wire N__5747;
    wire N__5742;
    wire N__5739;
    wire N__5736;
    wire N__5733;
    wire N__5728;
    wire N__5727;
    wire N__5726;
    wire N__5725;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5704;
    wire N__5699;
    wire N__5696;
    wire N__5691;
    wire N__5688;
    wire N__5677;
    wire N__5668;
    wire N__5665;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5649;
    wire N__5648;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5634;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5622;
    wire N__5617;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5604;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5596;
    wire N__5593;
    wire N__5586;
    wire N__5581;
    wire N__5578;
    wire N__5577;
    wire N__5576;
    wire N__5573;
    wire N__5568;
    wire N__5565;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5547;
    wire N__5542;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5505;
    wire N__5502;
    wire N__5497;
    wire N__5496;
    wire N__5493;
    wire N__5490;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5473;
    wire N__5470;
    wire N__5469;
    wire N__5466;
    wire N__5463;
    wire N__5462;
    wire N__5461;
    wire N__5456;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5434;
    wire N__5433;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5407;
    wire N__5404;
    wire N__5401;
    wire N__5400;
    wire N__5397;
    wire N__5394;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5292;
    wire N__5289;
    wire N__5286;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5265;
    wire N__5262;
    wire N__5259;
    wire N__5256;
    wire N__5253;
    wire N__5248;
    wire N__5247;
    wire N__5246;
    wire N__5245;
    wire N__5244;
    wire N__5243;
    wire N__5242;
    wire N__5241;
    wire N__5240;
    wire N__5239;
    wire N__5238;
    wire N__5237;
    wire N__5236;
    wire N__5235;
    wire N__5234;
    wire N__5233;
    wire N__5232;
    wire N__5231;
    wire N__5230;
    wire N__5229;
    wire N__5228;
    wire N__5227;
    wire N__5226;
    wire N__5225;
    wire N__5224;
    wire N__5223;
    wire N__5222;
    wire N__5167;
    wire N__5164;
    wire N__5161;
    wire N__5160;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5148;
    wire N__5145;
    wire N__5144;
    wire N__5137;
    wire N__5134;
    wire N__5133;
    wire N__5130;
    wire N__5127;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5101;
    wire N__5098;
    wire N__5095;
    wire N__5092;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5062;
    wire N__5061;
    wire N__5056;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5040;
    wire N__5037;
    wire N__5034;
    wire N__5029;
    wire N__5026;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5014;
    wire N__5013;
    wire N__5012;
    wire N__5011;
    wire N__5010;
    wire N__5007;
    wire N__5004;
    wire N__5003;
    wire N__5002;
    wire N__5001;
    wire N__5000;
    wire N__4997;
    wire N__4996;
    wire N__4993;
    wire N__4990;
    wire N__4989;
    wire N__4988;
    wire N__4987;
    wire N__4986;
    wire N__4985;
    wire N__4984;
    wire N__4983;
    wire N__4978;
    wire N__4975;
    wire N__4972;
    wire N__4967;
    wire N__4962;
    wire N__4959;
    wire N__4954;
    wire N__4953;
    wire N__4950;
    wire N__4949;
    wire N__4948;
    wire N__4947;
    wire N__4944;
    wire N__4939;
    wire N__4936;
    wire N__4933;
    wire N__4924;
    wire N__4923;
    wire N__4922;
    wire N__4919;
    wire N__4914;
    wire N__4909;
    wire N__4904;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4888;
    wire N__4885;
    wire N__4882;
    wire N__4871;
    wire N__4858;
    wire N__4857;
    wire N__4856;
    wire N__4855;
    wire N__4854;
    wire N__4853;
    wire N__4850;
    wire N__4849;
    wire N__4848;
    wire N__4847;
    wire N__4844;
    wire N__4837;
    wire N__4834;
    wire N__4833;
    wire N__4832;
    wire N__4831;
    wire N__4828;
    wire N__4821;
    wire N__4820;
    wire N__4819;
    wire N__4818;
    wire N__4815;
    wire N__4810;
    wire N__4807;
    wire N__4802;
    wire N__4801;
    wire N__4800;
    wire N__4799;
    wire N__4798;
    wire N__4797;
    wire N__4796;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4781;
    wire N__4772;
    wire N__4767;
    wire N__4762;
    wire N__4755;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4731;
    wire N__4728;
    wire N__4725;
    wire N__4724;
    wire N__4723;
    wire N__4722;
    wire N__4721;
    wire N__4720;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4708;
    wire N__4699;
    wire N__4696;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4668;
    wire N__4665;
    wire N__4660;
    wire N__4659;
    wire N__4658;
    wire N__4657;
    wire N__4656;
    wire N__4655;
    wire N__4654;
    wire N__4653;
    wire N__4652;
    wire N__4649;
    wire N__4648;
    wire N__4647;
    wire N__4646;
    wire N__4645;
    wire N__4644;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4631;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4619;
    wire N__4612;
    wire N__4609;
    wire N__4608;
    wire N__4607;
    wire N__4604;
    wire N__4603;
    wire N__4602;
    wire N__4601;
    wire N__4600;
    wire N__4599;
    wire N__4598;
    wire N__4593;
    wire N__4588;
    wire N__4581;
    wire N__4576;
    wire N__4571;
    wire N__4568;
    wire N__4563;
    wire N__4560;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4539;
    wire N__4534;
    wire N__4531;
    wire N__4522;
    wire N__4507;
    wire N__4504;
    wire N__4503;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4477;
    wire N__4476;
    wire N__4475;
    wire N__4472;
    wire N__4467;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4453;
    wire N__4452;
    wire N__4449;
    wire N__4448;
    wire N__4441;
    wire N__4438;
    wire N__4437;
    wire N__4436;
    wire N__4433;
    wire N__4428;
    wire N__4423;
    wire N__4420;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4412;
    wire N__4405;
    wire N__4402;
    wire N__4401;
    wire N__4400;
    wire N__4399;
    wire N__4398;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4369;
    wire N__4366;
    wire N__4365;
    wire N__4364;
    wire N__4363;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4348;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4330;
    wire N__4329;
    wire N__4326;
    wire N__4325;
    wire N__4322;
    wire N__4317;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4299;
    wire N__4296;
    wire N__4293;
    wire N__4282;
    wire N__4279;
    wire N__4276;
    wire N__4273;
    wire N__4270;
    wire N__4267;
    wire N__4266;
    wire N__4263;
    wire N__4260;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4245;
    wire N__4242;
    wire N__4239;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4222;
    wire N__4219;
    wire N__4218;
    wire N__4215;
    wire N__4212;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4200;
    wire N__4197;
    wire N__4194;
    wire N__4189;
    wire N__4188;
    wire N__4185;
    wire N__4182;
    wire N__4177;
    wire N__4174;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4149;
    wire N__4148;
    wire N__4147;
    wire N__4146;
    wire N__4145;
    wire N__4144;
    wire N__4141;
    wire N__4136;
    wire N__4131;
    wire N__4126;
    wire N__4117;
    wire N__4116;
    wire N__4115;
    wire N__4112;
    wire N__4107;
    wire N__4102;
    wire N__4101;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4078;
    wire N__4077;
    wire N__4076;
    wire N__4075;
    wire N__4072;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4061;
    wire N__4056;
    wire N__4055;
    wire N__4050;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4038;
    wire N__4035;
    wire N__4026;
    wire N__4021;
    wire N__4018;
    wire N__4017;
    wire N__4016;
    wire N__4015;
    wire N__4014;
    wire N__4011;
    wire N__4010;
    wire N__4009;
    wire N__4008;
    wire N__4007;
    wire N__4006;
    wire N__4005;
    wire N__4004;
    wire N__4003;
    wire N__4002;
    wire N__4001;
    wire N__4000;
    wire N__3999;
    wire N__3992;
    wire N__3991;
    wire N__3990;
    wire N__3983;
    wire N__3978;
    wire N__3977;
    wire N__3972;
    wire N__3971;
    wire N__3970;
    wire N__3963;
    wire N__3956;
    wire N__3953;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3941;
    wire N__3938;
    wire N__3935;
    wire N__3934;
    wire N__3931;
    wire N__3926;
    wire N__3921;
    wire N__3916;
    wire N__3913;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3893;
    wire N__3880;
    wire N__3879;
    wire N__3876;
    wire N__3875;
    wire N__3872;
    wire N__3867;
    wire N__3862;
    wire N__3859;
    wire N__3856;
    wire N__3855;
    wire N__3852;
    wire N__3851;
    wire N__3850;
    wire N__3849;
    wire N__3848;
    wire N__3847;
    wire N__3846;
    wire N__3843;
    wire N__3840;
    wire N__3837;
    wire N__3834;
    wire N__3831;
    wire N__3830;
    wire N__3827;
    wire N__3826;
    wire N__3825;
    wire N__3824;
    wire N__3823;
    wire N__3822;
    wire N__3819;
    wire N__3816;
    wire N__3815;
    wire N__3814;
    wire N__3813;
    wire N__3810;
    wire N__3805;
    wire N__3802;
    wire N__3799;
    wire N__3792;
    wire N__3789;
    wire N__3784;
    wire N__3781;
    wire N__3776;
    wire N__3769;
    wire N__3764;
    wire N__3753;
    wire N__3742;
    wire N__3739;
    wire N__3736;
    wire N__3733;
    wire N__3730;
    wire N__3727;
    wire N__3726;
    wire N__3723;
    wire N__3720;
    wire N__3715;
    wire N__3714;
    wire N__3711;
    wire N__3708;
    wire N__3703;
    wire N__3700;
    wire N__3699;
    wire N__3696;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3678;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3666;
    wire N__3661;
    wire N__3658;
    wire N__3655;
    wire N__3652;
    wire N__3649;
    wire N__3646;
    wire N__3643;
    wire N__3640;
    wire N__3639;
    wire N__3638;
    wire N__3637;
    wire N__3636;
    wire N__3635;
    wire N__3632;
    wire N__3627;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3617;
    wire N__3612;
    wire N__3609;
    wire N__3598;
    wire N__3597;
    wire N__3596;
    wire N__3593;
    wire N__3590;
    wire N__3587;
    wire N__3584;
    wire N__3581;
    wire N__3580;
    wire N__3577;
    wire N__3572;
    wire N__3569;
    wire N__3562;
    wire N__3559;
    wire N__3558;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3548;
    wire N__3541;
    wire N__3538;
    wire N__3535;
    wire N__3532;
    wire N__3529;
    wire N__3526;
    wire N__3523;
    wire N__3522;
    wire N__3519;
    wire N__3516;
    wire N__3513;
    wire N__3510;
    wire N__3505;
    wire N__3502;
    wire N__3499;
    wire N__3496;
    wire N__3493;
    wire N__3490;
    wire N__3487;
    wire N__3484;
    wire N__3481;
    wire N__3478;
    wire N__3475;
    wire N__3472;
    wire N__3469;
    wire N__3466;
    wire N__3463;
    wire N__3460;
    wire N__3457;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3445;
    wire N__3442;
    wire N__3439;
    wire N__3436;
    wire N__3433;
    wire N__3432;
    wire N__3429;
    wire N__3426;
    wire N__3423;
    wire N__3420;
    wire N__3415;
    wire N__3412;
    wire N__3409;
    wire N__3406;
    wire N__3403;
    wire N__3400;
    wire N__3397;
    wire N__3394;
    wire N__3391;
    wire N__3388;
    wire N__3385;
    wire N__3384;
    wire N__3381;
    wire N__3378;
    wire N__3373;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3363;
    wire N__3360;
    wire N__3357;
    wire N__3354;
    wire N__3351;
    wire N__3348;
    wire N__3343;
    wire N__3340;
    wire N__3337;
    wire N__3334;
    wire N__3331;
    wire N__3328;
    wire N__3325;
    wire N__3324;
    wire N__3323;
    wire N__3320;
    wire N__3317;
    wire N__3314;
    wire N__3307;
    wire N__3304;
    wire N__3301;
    wire N__3298;
    wire N__3295;
    wire N__3292;
    wire N__3289;
    wire N__3286;
    wire N__3283;
    wire N__3280;
    wire N__3279;
    wire N__3276;
    wire N__3273;
    wire N__3268;
    wire N__3267;
    wire N__3264;
    wire N__3261;
    wire N__3256;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3241;
    wire N__3240;
    wire N__3237;
    wire N__3234;
    wire N__3229;
    wire N__3226;
    wire N__3223;
    wire N__3222;
    wire N__3221;
    wire N__3216;
    wire N__3213;
    wire N__3208;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3190;
    wire N__3187;
    wire N__3184;
    wire N__3181;
    wire N__3178;
    wire N__3175;
    wire N__3172;
    wire N__3169;
    wire N__3166;
    wire N__3163;
    wire N__3160;
    wire N__3157;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3121;
    wire N__3118;
    wire N__3115;
    wire N__3112;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3097;
    wire N__3094;
    wire N__3091;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3070;
    wire N__3067;
    wire N__3064;
    wire N__3061;
    wire N__3058;
    wire N__3055;
    wire N__3052;
    wire N__3049;
    wire N__3046;
    wire N__3043;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3031;
    wire N__3028;
    wire N__3025;
    wire N__3022;
    wire N__3019;
    wire N__3016;
    wire N__3013;
    wire N__3010;
    wire N__3007;
    wire N__3004;
    wire N__3001;
    wire N__2998;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2986;
    wire N__2983;
    wire N__2980;
    wire N__2977;
    wire N__2974;
    wire N__2971;
    wire N__2968;
    wire N__2965;
    wire N__2962;
    wire N__2959;
    wire N__2956;
    wire N__2953;
    wire N__2950;
    wire N__2947;
    wire N__2944;
    wire N__2941;
    wire N__2938;
    wire N__2935;
    wire N__2932;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2920;
    wire N__2917;
    wire N__2914;
    wire N__2913;
    wire N__2910;
    wire N__2907;
    wire N__2902;
    wire N__2901;
    wire N__2898;
    wire N__2895;
    wire N__2890;
    wire N__2889;
    wire N__2886;
    wire N__2883;
    wire N__2878;
    wire N__2877;
    wire N__2874;
    wire N__2871;
    wire N__2866;
    wire N__2865;
    wire N__2862;
    wire N__2859;
    wire N__2854;
    wire N__2851;
    wire N__2850;
    wire N__2847;
    wire N__2844;
    wire N__2839;
    wire N__2836;
    wire N__2833;
    wire N__2830;
    wire N__2827;
    wire N__2824;
    wire N__2821;
    wire N__2818;
    wire N__2815;
    wire N__2812;
    wire N__2811;
    wire N__2808;
    wire N__2805;
    wire N__2800;
    wire N__2799;
    wire N__2798;
    wire N__2795;
    wire N__2792;
    wire N__2789;
    wire N__2786;
    wire N__2779;
    wire N__2776;
    wire N__2773;
    wire N__2770;
    wire N__2767;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2755;
    wire N__2752;
    wire N__2749;
    wire CLK40_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \INVU400_SDRAM.REFRESH_COUNTER_0C_net ;
    wire A_c_31;
    wire A_c_27;
    wire \INVU400_SDRAM.REFRESH_COUNTER_1C_net ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_0 ;
    wire bfn_2_4_0_;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_1 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_2 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_3 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_4 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_5 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_6 ;
    wire \U400_SDRAM.un3_REFRESH_COUNTER_cry_7 ;
    wire \INVU400_SDRAM.REFRESH_COUNTER_2C_net ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_8 ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U400_SDRAM.un1_REFRESH_COUNTERlt7_0_cascade_ ;
    wire \U400_SDRAM.REFRESH_COUNTERZ0Z_6 ;
    wire CASn_c;
    wire WEn_c;
    wire \INVU400_SDRAM.CASnC_net ;
    wire RASn_c;
    wire \INVU400_SDRAM.RASnC_net ;
    wire A_c_30;
    wire A_c_29;
    wire A_c_28;
    wire \U400_ADDRESS_DECODE.m2Z0Z_1 ;
    wire \INVU400_SDRAM.SDRAM_COUNTER_1C_net ;
    wire \INVU400_SDRAM.RAM_CYCLEC_net ;
    wire \U400_ADDRESS_DECODE.N_185_cascade_ ;
    wire \U400_ADDRESS_DECODE.m84_amZ0_cascade_ ;
    wire \U400_ADDRESS_DECODE.m84_bmZ0 ;
    wire N_85_0;
    wire \U400_ADDRESS_DECODE.N_46_0 ;
    wire \U400_ADDRESS_DECODE.N_47_0_cascade_ ;
    wire \U400_ADDRESS_DECODE.m71_amZ0Z_1 ;
    wire \U400_ADDRESS_DECODE.m71_amZ0_cascade_ ;
    wire \U400_ADDRESS_DECODE.m71_bmZ0 ;
    wire \U400_ADDRESS_DECODE.N_72_0_cascade_ ;
    wire N_73_0_cascade_;
    wire \INVU400_SDRAM.SDRAM_CMD_2C_net ;
    wire \U400_ADDRESS_DECODE.m56_amZ0 ;
    wire N_57_0;
    wire \U400_ADDRESS_DECODE.N_7_0_cascade_ ;
    wire \INVU400_SDRAM.SDRAM_CMD_0C_net ;
    wire RESETn_c_i;
    wire A_c_9;
    wire A_c_17;
    wire MA_c_7;
    wire A_c_18;
    wire A_c_24;
    wire MA_c_8;
    wire \INVU400_SDRAM.MA_nesr_7C_net ;
    wire A_c_8;
    wire A_c_16;
    wire MA_c_6;
    wire \INVU400_SDRAM.MA_nesr_6C_net ;
    wire bfn_5_3_0_;
    wire \U400_SDRAM.SDRAM_COUNTER_s_1 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_0 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_1 ;
    wire \U400_SDRAM.SDRAM_COUNTER_s_3 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_2 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_3 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_4 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_5 ;
    wire \U400_SDRAM.SDRAM_COUNTER_cry_6 ;
    wire \INVU400_SDRAM.SDRAM_COUNTER_2C_net ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U400_SDRAM.SDRAM_COUNTERZ0Z_4 ;
    wire N_60_cascade_;
    wire \U400_ADDRESS_DECODE.N_98_0_cascade_ ;
    wire U400_SDRAM_SDRAM_CMD_5_sqmuxa;
    wire \U400_ADDRESS_DECODE.m41_amZ0_cascade_ ;
    wire \U400_ADDRESS_DECODE.m41_bmZ0 ;
    wire \U400_ADDRESS_DECODE.m54Z0Z_0_cascade_ ;
    wire \U400_ADDRESS_DECODE.m56_bmZ0 ;
    wire \U400_ADDRESS_DECODE.N_185 ;
    wire \U400_ADDRESS_DECODE.N_185_mux_cascade_ ;
    wire \U400_ADDRESS_DECODE.N_42_0 ;
    wire \U400_ADDRESS_DECODE.m43_bmZ0_cascade_ ;
    wire N_44_0;
    wire \U400_ADDRESS_DECODE.N_33_0 ;
    wire \U400_ADDRESS_DECODE.m43_amZ0 ;
    wire \U400_ADDRESS_DECODE.m87_nsZ0Z_1 ;
    wire \U400_ADDRESS_DECODE.N_88_0_cascade_ ;
    wire N_96_0_cascade_;
    wire N_73_0;
    wire \INVU400_SDRAM.SDRAM_CMD_1C_net ;
    wire \U400_ADDRESS_DECODE.m63_nsZ0Z_1 ;
    wire \U400_ADDRESS_DECODE.N_139_0_cascade_ ;
    wire \U400_ADDRESS_DECODE.m133Z0Z_0 ;
    wire \U400_ADDRESS_DECODE.N_47_0 ;
    wire \U400_ADDRESS_DECODE.N_62_0 ;
    wire \U400_ADDRESS_DECODE.N_62_0_cascade_ ;
    wire \U400_ADDRESS_DECODE.m141_bmZ0_cascade_ ;
    wire \U400_ADDRESS_DECODE.m141_amZ0 ;
    wire \U400_SDRAM.CS0_ENZ0 ;
    wire CS0n_c;
    wire \INVU400_SDRAM.CS0_ENC_net ;
    wire A_c_26;
    wire MA_c_12;
    wire A_c_19;
    wire MA_c_9;
    wire \INVU400_SDRAM.MA_nesr_12C_net ;
    wire U400_SDRAM_RAM_CYCLE;
    wire U400_SDRAM_RAM_CYCLE_START_2_0;
    wire \U400_ADDRESS_DECODE.N_8_0_cascade_ ;
    wire \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2 ;
    wire TSn_c;
    wire \U400_ADDRESS_DECODE.m165_nsZ0Z_1 ;
    wire N_13_0_cascade_;
    wire \U400_ADDRESS_DECODE.N_10_0 ;
    wire \U400_ADDRESS_DECODE.N_8_0 ;
    wire \U400_ADDRESS_DECODE.N_179_mux_cascade_ ;
    wire \U400_ADDRESS_DECODE.m94_amZ0Z_1 ;
    wire \U400_ADDRESS_DECODE.m94_amZ0_cascade_ ;
    wire \U400_ADDRESS_DECODE.N_95_0 ;
    wire U400_SDRAM_RAM_CYCLE_START;
    wire \U400_ADDRESS_DECODE.N_15_0 ;
    wire N_13_0;
    wire U400_SDRAM_SDRAM_CMD11;
    wire \U400_ADDRESS_DECODE.m20_amZ0_cascade_ ;
    wire U400_SDRAM_SDRAM_COUNTER_3;
    wire \U400_ADDRESS_DECODE.N_6_0 ;
    wire \U400_ADDRESS_DECODE.m94_bmZ0 ;
    wire U400_SDRAM_SDRAM_COUNTER_1;
    wire \U400_ADDRESS_DECODE.m20_bmZ0 ;
    wire \U400_ADDRESS_DECODE.N_20_0 ;
    wire \U400_ADDRESS_DECODE.N_179_mux ;
    wire RnW_c;
    wire U400_SDRAM_WRITE_CYCLE;
    wire N_48;
    wire N_142_0;
    wire \INVU400_SDRAM.WRITE_CYCLEC_net ;
    wire \U400_ADDRESS_DECODE.N_12_0 ;
    wire \U400_ADDRESS_DECODE.N_21_0 ;
    wire A_c_23;
    wire N_137_0;
    wire N_190_mux;
    wire N_138_0;
    wire N_23_0;
    wire \U400_SDRAM.CS1_ENZ0 ;
    wire CS1n_c;
    wire \INVU400_SDRAM.CS1_ENC_net ;
    wire U400_SDRAM_TA_COUNTER_4;
    wire U400_SDRAM_TA_COUNTER_1;
    wire \U400_ADDRESS_DECODE.N_177_mux_cascade_ ;
    wire U400_SDRAM_TA_COUNTER_0;
    wire U400_SDRAM_TACK;
    wire U400_SDRAM_TA_COUNTER_5;
    wire \U400_SDRAM.N_252_0_0_cascade_ ;
    wire U400_SDRAM_TA_COUNTER_2;
    wire U400_SDRAM_TA_COUNTER_3;
    wire A_c_22;
    wire BANK1_c;
    wire A_c_21;
    wire U400_SDRAM_un1_SDRAM_COUNTER59_2_0;
    wire BANK0_c;
    wire U400_SDRAM_SDRAM_CMD_1_sqmuxa_1;
    wire \INVU400_SDRAM.BANK1C_net ;
    wire U400_SDRAM_SDRAM_COUNTER_2;
    wire N_60;
    wire \U400_ADDRESS_DECODE.m145_nsZ0Z_1 ;
    wire N_100_0_i;
    wire CONSTANT_ONE_NET;
    wire U400_SDRAM_SDRAM_COUNTER_0;
    wire \INVU400_SDRAM.SDRAM_COUNTER_0C_net ;
    wire U400_SDRAM_SDRAM_COUNTERe_0_i;
    wire \U400_ADDRESS_DECODE.N_135_0 ;
    wire \U400_ADDRESS_DECODE.N_146_0 ;
    wire N_14_i;
    wire \U400_ADDRESS_DECODE.N_147_0_cascade_ ;
    wire \U400_ADDRESS_DECODE.N_136_0 ;
    wire N_43;
    wire A_c_20;
    wire MA_c_10;
    wire A_c_25;
    wire MA_c_11;
    wire \INVU400_SDRAM.MA_nesr_10C_net ;
    wire \U400_ADDRESS_DECODE.N_4_0_cascade_ ;
    wire N_124_0;
    wire \U400_SDRAM.N_252_0_0 ;
    wire \U400_SDRAM.N_252_0_0_en ;
    wire N_174;
    wire U400_SDRAM_TA_OUT_5_0;
    wire U400_SDRAM_N_252_0;
    wire TA_OUT;
    wire CLK40_c_g;
    wire U400_SDRAM_BURST;
    wire \U400_ADDRESS_DECODE.N_114_0 ;
    wire N_65_0;
    wire U400_SDRAM_SDRAM_CONFIGURED;
    wire \INVU400_SDRAM.SDRAM_CONFIGUREDC_net ;
    wire N_129_0;
    wire N_127_0;
    wire A_c_1;
    wire N_128_0;
    wire \U400_ADDRESS_DECODE.N_122_0 ;
    wire SIZ_c_0;
    wire A_c_0;
    wire \U400_ADDRESS_DECODE.N_4_0 ;
    wire SIZ_c_1;
    wire \U400_ADDRESS_DECODE.N_186_mux ;
    wire A_c_7;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_1 ;
    wire A_c_3;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_0 ;
    wire A_c_11;
    wire \U400_SDRAM.MA_5_iv_0_1 ;
    wire MA_c_1;
    wire A_c_15;
    wire \U400_SDRAM.MA_5_iv_0_5 ;
    wire MA_c_5;
    wire A_c_5;
    wire A_c_13;
    wire MA_c_3;
    wire \INVU400_SDRAM.MA_nesr_1C_net ;
    wire A_c_4;
    wire A_c_12;
    wire MA_c_2;
    wire A_c_6;
    wire A_c_14;
    wire MA_c_4;
    wire A_c_2;
    wire \U400_SDRAM.SDRAM_CMDZ0Z_2 ;
    wire A_c_10;
    wire \U400_SDRAM.MA19 ;
    wire MA_c_0;
    wire \INVU400_SDRAM.MA_nesr_2C_net ;
    wire \U400_SDRAM.un1_MA20_0_i_0 ;
    wire RESETn_c_i_g;
    wire \U400_ADDRESS_DECODE.N_170_mux ;
    wire RESETn_c;
    wire N_4_0_i;
    wire TA_EN_i;
    wire N_304_i;
    wire _gnd_net_;

    IO_PAD MA_obuf_7_iopad (
            .OE(N__7469),
            .DIN(N__7468),
            .DOUT(N__7467),
            .PACKAGEPIN(MA[7]));
    defparam MA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_7_preio (
            .PADOEN(N__7469),
            .PADOUT(N__7468),
            .PADIN(N__7467),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3037),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__7460),
            .DIN(N__7459),
            .DOUT(N__7458),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__7460),
            .PADOUT(N__7459),
            .PADIN(N__7458),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__7451),
            .DIN(N__7450),
            .DOUT(N__7449),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__7451),
            .PADOUT(N__7450),
            .PADIN(N__7449),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2839),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__7442),
            .DIN(N__7441),
            .DOUT(N__7440),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__7442),
            .PADOUT(N__7441),
            .PADIN(N__7440),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5104),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_8_iopad (
            .OE(N__7433),
            .DIN(N__7432),
            .DOUT(N__7431),
            .PACKAGEPIN(MA[8]));
    defparam MA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_8_preio (
            .PADOEN(N__7433),
            .PADOUT(N__7432),
            .PADIN(N__7431),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3175),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_10_iopad (
            .OE(N__7424),
            .DIN(N__7423),
            .DOUT(N__7422),
            .PACKAGEPIN(MA[10]));
    defparam MA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_10_preio (
            .PADOEN(N__7424),
            .PADOUT(N__7423),
            .PADIN(N__7422),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5356),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__7415),
            .DIN(N__7414),
            .DOUT(N__7413),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__7415),
            .PADOUT(N__7414),
            .PADIN(N__7413),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_2_iopad (
            .OE(N__7406),
            .DIN(N__7405),
            .DOUT(N__7404),
            .PACKAGEPIN(MA[2]));
    defparam MA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_2_preio (
            .PADOEN(N__7406),
            .PADOUT(N__7405),
            .PADIN(N__7404),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6097),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__7397),
            .DIN(N__7396),
            .DOUT(N__7395),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__7397),
            .PADOUT(N__7396),
            .PADIN(N__7395),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__7388),
            .DIN(N__7387),
            .DOUT(N__7386),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__7388),
            .PADOUT(N__7387),
            .PADIN(N__7386),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__7379),
            .DIN(N__7378),
            .DOUT(N__7377),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__7379),
            .PADOUT(N__7378),
            .PADIN(N__7377),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5317),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__7370),
            .DIN(N__7369),
            .DOUT(N__7368),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__7370),
            .PADOUT(N__7369),
            .PADIN(N__7368),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__7361),
            .DIN(N__7360),
            .DOUT(N__7359),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__7361),
            .PADOUT(N__7360),
            .PADIN(N__7359),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__7352),
            .DIN(N__7351),
            .DOUT(N__7350),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__7352),
            .PADOUT(N__7351),
            .PADIN(N__7350),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_12_iopad (
            .OE(N__7343),
            .DIN(N__7342),
            .DOUT(N__7341),
            .PACKAGEPIN(MA[12]));
    defparam MA_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_12_preio (
            .PADOEN(N__7343),
            .PADOUT(N__7342),
            .PADIN(N__7341),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3469),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_1_iopad (
            .OE(N__7334),
            .DIN(N__7333),
            .DOUT(N__7332),
            .PACKAGEPIN(MA[1]));
    defparam MA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_1_preio (
            .PADOEN(N__7334),
            .PADOUT(N__7333),
            .PADIN(N__7332),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6208),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__7325),
            .DIN(N__7324),
            .DOUT(N__7323),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__7325),
            .PADOUT(N__7324),
            .PADIN(N__7323),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__7316),
            .DIN(N__7315),
            .DOUT(N__7314),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__7316),
            .PADOUT(N__7315),
            .PADIN(N__7314),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__7307),
            .DIN(N__7306),
            .DOUT(N__7305),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__7307),
            .PADOUT(N__7306),
            .PADIN(N__7305),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_4_iopad (
            .OE(N__7298),
            .DIN(N__7297),
            .DOUT(N__7296),
            .PACKAGEPIN(MA[4]));
    defparam MA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_4_preio (
            .PADOEN(N__7298),
            .PADOUT(N__7297),
            .PADIN(N__7296),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6064),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__7289),
            .DIN(N__7288),
            .DOUT(N__7287),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__7289),
            .PADOUT(N__7288),
            .PADIN(N__7287),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__7280),
            .DIN(N__7279),
            .DOUT(N__7278),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__7280),
            .PADOUT(N__7279),
            .PADIN(N__7278),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__7271),
            .DIN(N__7270),
            .DOUT(N__7269),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__7271),
            .PADOUT(N__7270),
            .PADIN(N__7269),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5668),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__7262),
            .DIN(N__7261),
            .DOUT(N__7260),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__7262),
            .PADOUT(N__7261),
            .PADIN(N__7260),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_9_iopad (
            .OE(N__7253),
            .DIN(N__7252),
            .DOUT(N__7251),
            .PACKAGEPIN(MA[9]));
    defparam MA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_9_preio (
            .PADOEN(N__7253),
            .PADOUT(N__7252),
            .PADIN(N__7251),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3442),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__7244),
            .DIN(N__7243),
            .DOUT(N__7242),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__7244),
            .PADOUT(N__7243),
            .PADIN(N__7242),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5659),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__7235),
            .DIN(N__7234),
            .DOUT(N__7233),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__7235),
            .PADOUT(N__7234),
            .PADIN(N__7233),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__7226),
            .DIN(N__7225),
            .DOUT(N__7224),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__7226),
            .PADOUT(N__7225),
            .PADIN(N__7224),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__7217),
            .DIN(N__7216),
            .DOUT(N__7215),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__7217),
            .PADOUT(N__7216),
            .PADIN(N__7215),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4687),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__7208),
            .DIN(N__7207),
            .DOUT(N__7206),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__7208),
            .PADOUT(N__7207),
            .PADIN(N__7206),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__7199),
            .DIN(N__7198),
            .DOUT(N__7197),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__7199),
            .PADOUT(N__7198),
            .PADIN(N__7197),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_3_iopad (
            .OE(N__7190),
            .DIN(N__7189),
            .DOUT(N__7188),
            .PACKAGEPIN(MA[3]));
    defparam MA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_3_preio (
            .PADOEN(N__7190),
            .PADOUT(N__7189),
            .PADIN(N__7188),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6139),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__7181),
            .DIN(N__7180),
            .DOUT(N__7179),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__7181),
            .PADOUT(N__7180),
            .PADIN(N__7179),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__7172),
            .DIN(N__7171),
            .DOUT(N__7170),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__7172),
            .PADOUT(N__7171),
            .PADIN(N__7170),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__7163),
            .DIN(N__7162),
            .DOUT(N__7161),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__7163),
            .PADOUT(N__7162),
            .PADIN(N__7161),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_6_iopad (
            .OE(N__7154),
            .DIN(N__7153),
            .DOUT(N__7152),
            .PACKAGEPIN(MA[6]));
    defparam MA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_6_preio (
            .PADOEN(N__7154),
            .PADOUT(N__7153),
            .PADIN(N__7152),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3136),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__7145),
            .DIN(N__7144),
            .DOUT(N__7143),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__7145),
            .PADOUT(N__7144),
            .PADIN(N__7143),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__7136),
            .DIN(N__7135),
            .DOUT(N__7134),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__7136),
            .PADOUT(N__7135),
            .PADIN(N__7134),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__7127),
            .DIN(N__7126),
            .DOUT(N__7125),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__7127),
            .PADOUT(N__7126),
            .PADIN(N__7125),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__7118),
            .DIN(N__7117),
            .DOUT(N__7116),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__7118),
            .PADOUT(N__7117),
            .PADIN(N__7116),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2986),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__7109),
            .DIN(N__7108),
            .DOUT(N__7107),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__7109),
            .PADOUT(N__7108),
            .PADIN(N__7107),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__7100),
            .DIN(N__7099),
            .DOUT(N__7098),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__7100),
            .PADOUT(N__7099),
            .PADIN(N__7098),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5053),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_11_iopad (
            .OE(N__7091),
            .DIN(N__7090),
            .DOUT(N__7089),
            .PACKAGEPIN(MA[11]));
    defparam MA_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_11_preio (
            .PADOEN(N__7091),
            .PADOUT(N__7090),
            .PADIN(N__7089),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5329),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TAn_obuft_iopad (
            .OE(N__7082),
            .DIN(N__7081),
            .DOUT(N__7080),
            .PACKAGEPIN(TAn));
    defparam TAn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TAn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TAn_obuft_preio (
            .PADOEN(N__7082),
            .PADOUT(N__7081),
            .PADIN(N__7080),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6427),
            .DIN0(),
            .DOUT0(N__5269),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__7073),
            .DIN(N__7072),
            .DOUT(N__7071),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__7073),
            .PADOUT(N__7072),
            .PADIN(N__7071),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_5_iopad (
            .OE(N__7064),
            .DIN(N__7063),
            .DOUT(N__7062),
            .PACKAGEPIN(MA[5]));
    defparam MA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_5_preio (
            .PADOEN(N__7064),
            .PADOUT(N__7063),
            .PADIN(N__7062),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6184),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__7055),
            .DIN(N__7054),
            .DOUT(N__7053),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__7055),
            .PADOUT(N__7054),
            .PADIN(N__7053),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__7046),
            .DIN(N__7045),
            .DOUT(N__7044),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__7046),
            .PADOUT(N__7045),
            .PADIN(N__7044),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LBENn_obuf_iopad.PULLUP=1'b1;
    IO_PAD LBENn_obuf_iopad (
            .OE(N__7037),
            .DIN(N__7036),
            .DOUT(N__7035),
            .PACKAGEPIN(LBENn));
    defparam LBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LBENn_obuf_preio (
            .PADOEN(N__7037),
            .PADOUT(N__7036),
            .PADIN(N__7035),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6454),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__7028),
            .DIN(N__7027),
            .DOUT(N__7026),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__7028),
            .PADOUT(N__7027),
            .PADIN(N__7026),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CS1n_obuf_iopad (
            .OE(N__7019),
            .DIN(N__7018),
            .DOUT(N__7017),
            .PACKAGEPIN(CS1n));
    defparam CS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CS1n_obuf_preio (
            .PADOEN(N__7019),
            .PADOUT(N__7018),
            .PADIN(N__7017),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4174),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__7010),
            .DIN(N__7009),
            .DOUT(N__7008),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__7010),
            .PADOUT(N__7009),
            .PADIN(N__7008),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__7001),
            .DIN(N__7000),
            .DOUT(N__6999),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__7001),
            .PADOUT(N__7000),
            .PADIN(N__6999),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__6992),
            .DIN(N__6991),
            .DOUT(N__6990),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__6992),
            .PADOUT(N__6991),
            .PADIN(N__6990),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__6983),
            .DIN(N__6982),
            .DOUT(N__6981),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__6983),
            .PADOUT(N__6982),
            .PADIN(N__6981),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__6974),
            .DIN(N__6973),
            .DOUT(N__6972),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__6974),
            .PADOUT(N__6973),
            .PADIN(N__6972),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2995),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MA_obuf_0_iopad (
            .OE(N__6965),
            .DIN(N__6964),
            .DOUT(N__6963),
            .PACKAGEPIN(MA[0]));
    defparam MA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam MA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO MA_obuf_0_preio (
            .PADOEN(N__6965),
            .PADOUT(N__6964),
            .PADIN(N__6963),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6808),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__6956),
            .DIN(N__6955),
            .DOUT(N__6954),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__6956),
            .PADOUT(N__6955),
            .PADIN(N__6954),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__6947),
            .DIN(N__6946),
            .DOUT(N__6945),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__6947),
            .PADOUT(N__6946),
            .PADIN(N__6945),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__6938),
            .DIN(N__6937),
            .DOUT(N__6936),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__6938),
            .PADOUT(N__6937),
            .PADIN(N__6936),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CS0n_obuf_iopad (
            .OE(N__6929),
            .DIN(N__6928),
            .DOUT(N__6927),
            .PACKAGEPIN(CS0n));
    defparam CS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CS0n_obuf_preio (
            .PADOEN(N__6929),
            .PADOUT(N__6928),
            .PADIN(N__6927),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3505),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__6920),
            .DIN(N__6919),
            .DOUT(N__6918),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__6920),
            .PADOUT(N__6919),
            .PADIN(N__6918),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__6911),
            .DIN(N__6910),
            .DOUT(N__6909),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__6911),
            .PADOUT(N__6910),
            .PADIN(N__6909),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5614),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__6902),
            .DIN(N__6901),
            .DOUT(N__6900),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__6902),
            .PADOUT(N__6901),
            .PADIN(N__6900),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_ibuf_gb_io_iopad (
            .OE(N__6893),
            .DIN(N__6892),
            .DOUT(N__6891),
            .PACKAGEPIN(CLK40));
    defparam CLK40_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_ibuf_gb_io_preio (
            .PADOEN(N__6893),
            .PADOUT(N__6892),
            .PADIN(N__6891),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__1627 (
            .O(N__6874),
            .I(N__6871));
    InMux I__1626 (
            .O(N__6871),
            .I(N__6868));
    LocalMux I__1625 (
            .O(N__6868),
            .I(N__6865));
    Span4Mux_s1_v I__1624 (
            .O(N__6865),
            .I(N__6862));
    Odrv4 I__1623 (
            .O(N__6862),
            .I(A_c_10));
    InMux I__1622 (
            .O(N__6859),
            .I(N__6853));
    InMux I__1621 (
            .O(N__6858),
            .I(N__6853));
    LocalMux I__1620 (
            .O(N__6853),
            .I(N__6846));
    InMux I__1619 (
            .O(N__6852),
            .I(N__6843));
    InMux I__1618 (
            .O(N__6851),
            .I(N__6836));
    InMux I__1617 (
            .O(N__6850),
            .I(N__6836));
    InMux I__1616 (
            .O(N__6849),
            .I(N__6836));
    Span4Mux_h I__1615 (
            .O(N__6846),
            .I(N__6830));
    LocalMux I__1614 (
            .O(N__6843),
            .I(N__6827));
    LocalMux I__1613 (
            .O(N__6836),
            .I(N__6824));
    InMux I__1612 (
            .O(N__6835),
            .I(N__6817));
    InMux I__1611 (
            .O(N__6834),
            .I(N__6817));
    InMux I__1610 (
            .O(N__6833),
            .I(N__6817));
    Odrv4 I__1609 (
            .O(N__6830),
            .I(\U400_SDRAM.MA19 ));
    Odrv12 I__1608 (
            .O(N__6827),
            .I(\U400_SDRAM.MA19 ));
    Odrv4 I__1607 (
            .O(N__6824),
            .I(\U400_SDRAM.MA19 ));
    LocalMux I__1606 (
            .O(N__6817),
            .I(\U400_SDRAM.MA19 ));
    IoInMux I__1605 (
            .O(N__6808),
            .I(N__6805));
    LocalMux I__1604 (
            .O(N__6805),
            .I(MA_c_0));
    CEMux I__1603 (
            .O(N__6802),
            .I(N__6797));
    CEMux I__1602 (
            .O(N__6801),
            .I(N__6794));
    CEMux I__1601 (
            .O(N__6800),
            .I(N__6791));
    LocalMux I__1600 (
            .O(N__6797),
            .I(N__6787));
    LocalMux I__1599 (
            .O(N__6794),
            .I(N__6784));
    LocalMux I__1598 (
            .O(N__6791),
            .I(N__6781));
    CEMux I__1597 (
            .O(N__6790),
            .I(N__6778));
    Span4Mux_v I__1596 (
            .O(N__6787),
            .I(N__6767));
    Span4Mux_h I__1595 (
            .O(N__6784),
            .I(N__6767));
    Span4Mux_s2_v I__1594 (
            .O(N__6781),
            .I(N__6767));
    LocalMux I__1593 (
            .O(N__6778),
            .I(N__6767));
    CEMux I__1592 (
            .O(N__6777),
            .I(N__6764));
    CEMux I__1591 (
            .O(N__6776),
            .I(N__6761));
    Odrv4 I__1590 (
            .O(N__6767),
            .I(\U400_SDRAM.un1_MA20_0_i_0 ));
    LocalMux I__1589 (
            .O(N__6764),
            .I(\U400_SDRAM.un1_MA20_0_i_0 ));
    LocalMux I__1588 (
            .O(N__6761),
            .I(\U400_SDRAM.un1_MA20_0_i_0 ));
    CascadeMux I__1587 (
            .O(N__6754),
            .I(N__6751));
    InMux I__1586 (
            .O(N__6751),
            .I(N__6748));
    LocalMux I__1585 (
            .O(N__6748),
            .I(N__6743));
    SRMux I__1584 (
            .O(N__6747),
            .I(N__6697));
    SRMux I__1583 (
            .O(N__6746),
            .I(N__6697));
    Glb2LocalMux I__1582 (
            .O(N__6743),
            .I(N__6697));
    SRMux I__1581 (
            .O(N__6742),
            .I(N__6697));
    SRMux I__1580 (
            .O(N__6741),
            .I(N__6697));
    SRMux I__1579 (
            .O(N__6740),
            .I(N__6697));
    SRMux I__1578 (
            .O(N__6739),
            .I(N__6697));
    SRMux I__1577 (
            .O(N__6738),
            .I(N__6697));
    SRMux I__1576 (
            .O(N__6737),
            .I(N__6697));
    SRMux I__1575 (
            .O(N__6736),
            .I(N__6697));
    SRMux I__1574 (
            .O(N__6735),
            .I(N__6697));
    SRMux I__1573 (
            .O(N__6734),
            .I(N__6697));
    SRMux I__1572 (
            .O(N__6733),
            .I(N__6697));
    SRMux I__1571 (
            .O(N__6732),
            .I(N__6697));
    SRMux I__1570 (
            .O(N__6731),
            .I(N__6697));
    SRMux I__1569 (
            .O(N__6730),
            .I(N__6697));
    GlobalMux I__1568 (
            .O(N__6697),
            .I(N__6694));
    gio2CtrlBuf I__1567 (
            .O(N__6694),
            .I(RESETn_c_i_g));
    CascadeMux I__1566 (
            .O(N__6691),
            .I(N__6688));
    InMux I__1565 (
            .O(N__6688),
            .I(N__6682));
    CascadeMux I__1564 (
            .O(N__6687),
            .I(N__6679));
    InMux I__1563 (
            .O(N__6686),
            .I(N__6676));
    InMux I__1562 (
            .O(N__6685),
            .I(N__6673));
    LocalMux I__1561 (
            .O(N__6682),
            .I(N__6670));
    InMux I__1560 (
            .O(N__6679),
            .I(N__6667));
    LocalMux I__1559 (
            .O(N__6676),
            .I(N__6664));
    LocalMux I__1558 (
            .O(N__6673),
            .I(N__6661));
    Span4Mux_h I__1557 (
            .O(N__6670),
            .I(N__6656));
    LocalMux I__1556 (
            .O(N__6667),
            .I(N__6656));
    Span12Mux_s8_h I__1555 (
            .O(N__6664),
            .I(N__6653));
    Span4Mux_v I__1554 (
            .O(N__6661),
            .I(N__6650));
    Span4Mux_v I__1553 (
            .O(N__6656),
            .I(N__6647));
    Odrv12 I__1552 (
            .O(N__6653),
            .I(\U400_ADDRESS_DECODE.N_170_mux ));
    Odrv4 I__1551 (
            .O(N__6650),
            .I(\U400_ADDRESS_DECODE.N_170_mux ));
    Odrv4 I__1550 (
            .O(N__6647),
            .I(\U400_ADDRESS_DECODE.N_170_mux ));
    CascadeMux I__1549 (
            .O(N__6640),
            .I(N__6636));
    InMux I__1548 (
            .O(N__6639),
            .I(N__6632));
    InMux I__1547 (
            .O(N__6636),
            .I(N__6627));
    InMux I__1546 (
            .O(N__6635),
            .I(N__6627));
    LocalMux I__1545 (
            .O(N__6632),
            .I(N__6621));
    LocalMux I__1544 (
            .O(N__6627),
            .I(N__6618));
    InMux I__1543 (
            .O(N__6626),
            .I(N__6613));
    InMux I__1542 (
            .O(N__6625),
            .I(N__6613));
    CascadeMux I__1541 (
            .O(N__6624),
            .I(N__6599));
    Span4Mux_s3_v I__1540 (
            .O(N__6621),
            .I(N__6591));
    Span4Mux_h I__1539 (
            .O(N__6618),
            .I(N__6591));
    LocalMux I__1538 (
            .O(N__6613),
            .I(N__6591));
    InMux I__1537 (
            .O(N__6612),
            .I(N__6588));
    InMux I__1536 (
            .O(N__6611),
            .I(N__6585));
    CascadeMux I__1535 (
            .O(N__6610),
            .I(N__6582));
    InMux I__1534 (
            .O(N__6609),
            .I(N__6575));
    InMux I__1533 (
            .O(N__6608),
            .I(N__6575));
    InMux I__1532 (
            .O(N__6607),
            .I(N__6572));
    InMux I__1531 (
            .O(N__6606),
            .I(N__6569));
    InMux I__1530 (
            .O(N__6605),
            .I(N__6562));
    InMux I__1529 (
            .O(N__6604),
            .I(N__6562));
    InMux I__1528 (
            .O(N__6603),
            .I(N__6562));
    InMux I__1527 (
            .O(N__6602),
            .I(N__6557));
    InMux I__1526 (
            .O(N__6599),
            .I(N__6557));
    CascadeMux I__1525 (
            .O(N__6598),
            .I(N__6552));
    Span4Mux_h I__1524 (
            .O(N__6591),
            .I(N__6547));
    LocalMux I__1523 (
            .O(N__6588),
            .I(N__6547));
    LocalMux I__1522 (
            .O(N__6585),
            .I(N__6544));
    InMux I__1521 (
            .O(N__6582),
            .I(N__6541));
    InMux I__1520 (
            .O(N__6581),
            .I(N__6538));
    InMux I__1519 (
            .O(N__6580),
            .I(N__6535));
    LocalMux I__1518 (
            .O(N__6575),
            .I(N__6530));
    LocalMux I__1517 (
            .O(N__6572),
            .I(N__6530));
    LocalMux I__1516 (
            .O(N__6569),
            .I(N__6523));
    LocalMux I__1515 (
            .O(N__6562),
            .I(N__6523));
    LocalMux I__1514 (
            .O(N__6557),
            .I(N__6523));
    InMux I__1513 (
            .O(N__6556),
            .I(N__6520));
    InMux I__1512 (
            .O(N__6555),
            .I(N__6516));
    InMux I__1511 (
            .O(N__6552),
            .I(N__6513));
    Span4Mux_v I__1510 (
            .O(N__6547),
            .I(N__6510));
    Span4Mux_h I__1509 (
            .O(N__6544),
            .I(N__6505));
    LocalMux I__1508 (
            .O(N__6541),
            .I(N__6505));
    LocalMux I__1507 (
            .O(N__6538),
            .I(N__6500));
    LocalMux I__1506 (
            .O(N__6535),
            .I(N__6500));
    Span4Mux_v I__1505 (
            .O(N__6530),
            .I(N__6493));
    Span4Mux_h I__1504 (
            .O(N__6523),
            .I(N__6493));
    LocalMux I__1503 (
            .O(N__6520),
            .I(N__6493));
    InMux I__1502 (
            .O(N__6519),
            .I(N__6490));
    LocalMux I__1501 (
            .O(N__6516),
            .I(N__6485));
    LocalMux I__1500 (
            .O(N__6513),
            .I(N__6485));
    Span4Mux_h I__1499 (
            .O(N__6510),
            .I(N__6480));
    Span4Mux_h I__1498 (
            .O(N__6505),
            .I(N__6480));
    Span4Mux_v I__1497 (
            .O(N__6500),
            .I(N__6477));
    Span4Mux_h I__1496 (
            .O(N__6493),
            .I(N__6472));
    LocalMux I__1495 (
            .O(N__6490),
            .I(N__6472));
    Span12Mux_s8_v I__1494 (
            .O(N__6485),
            .I(N__6469));
    IoSpan4Mux I__1493 (
            .O(N__6480),
            .I(N__6466));
    Span4Mux_h I__1492 (
            .O(N__6477),
            .I(N__6461));
    Span4Mux_v I__1491 (
            .O(N__6472),
            .I(N__6461));
    Odrv12 I__1490 (
            .O(N__6469),
            .I(RESETn_c));
    Odrv4 I__1489 (
            .O(N__6466),
            .I(RESETn_c));
    Odrv4 I__1488 (
            .O(N__6461),
            .I(RESETn_c));
    IoInMux I__1487 (
            .O(N__6454),
            .I(N__6451));
    LocalMux I__1486 (
            .O(N__6451),
            .I(N__6448));
    Odrv4 I__1485 (
            .O(N__6448),
            .I(N_4_0_i));
    InMux I__1484 (
            .O(N__6445),
            .I(N__6442));
    LocalMux I__1483 (
            .O(N__6442),
            .I(N__6439));
    Span4Mux_v I__1482 (
            .O(N__6439),
            .I(N__6435));
    InMux I__1481 (
            .O(N__6438),
            .I(N__6432));
    Odrv4 I__1480 (
            .O(N__6435),
            .I(TA_EN_i));
    LocalMux I__1479 (
            .O(N__6432),
            .I(TA_EN_i));
    IoInMux I__1478 (
            .O(N__6427),
            .I(N__6424));
    LocalMux I__1477 (
            .O(N__6424),
            .I(N__6421));
    Odrv4 I__1476 (
            .O(N__6421),
            .I(N_304_i));
    InMux I__1475 (
            .O(N__6418),
            .I(N__6415));
    LocalMux I__1474 (
            .O(N__6415),
            .I(N__6412));
    Odrv4 I__1473 (
            .O(N__6412),
            .I(A_c_7));
    CascadeMux I__1472 (
            .O(N__6409),
            .I(N__6404));
    InMux I__1471 (
            .O(N__6408),
            .I(N__6396));
    InMux I__1470 (
            .O(N__6407),
            .I(N__6396));
    InMux I__1469 (
            .O(N__6404),
            .I(N__6391));
    InMux I__1468 (
            .O(N__6403),
            .I(N__6391));
    InMux I__1467 (
            .O(N__6402),
            .I(N__6383));
    InMux I__1466 (
            .O(N__6401),
            .I(N__6383));
    LocalMux I__1465 (
            .O(N__6396),
            .I(N__6380));
    LocalMux I__1464 (
            .O(N__6391),
            .I(N__6377));
    InMux I__1463 (
            .O(N__6390),
            .I(N__6372));
    InMux I__1462 (
            .O(N__6389),
            .I(N__6372));
    InMux I__1461 (
            .O(N__6388),
            .I(N__6368));
    LocalMux I__1460 (
            .O(N__6383),
            .I(N__6358));
    Span4Mux_h I__1459 (
            .O(N__6380),
            .I(N__6358));
    Span4Mux_h I__1458 (
            .O(N__6377),
            .I(N__6358));
    LocalMux I__1457 (
            .O(N__6372),
            .I(N__6358));
    InMux I__1456 (
            .O(N__6371),
            .I(N__6354));
    LocalMux I__1455 (
            .O(N__6368),
            .I(N__6351));
    InMux I__1454 (
            .O(N__6367),
            .I(N__6348));
    Span4Mux_v I__1453 (
            .O(N__6358),
            .I(N__6345));
    InMux I__1452 (
            .O(N__6357),
            .I(N__6342));
    LocalMux I__1451 (
            .O(N__6354),
            .I(N__6339));
    Span4Mux_h I__1450 (
            .O(N__6351),
            .I(N__6334));
    LocalMux I__1449 (
            .O(N__6348),
            .I(N__6334));
    Span4Mux_v I__1448 (
            .O(N__6345),
            .I(N__6331));
    LocalMux I__1447 (
            .O(N__6342),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1446 (
            .O(N__6339),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1445 (
            .O(N__6334),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1444 (
            .O(N__6331),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_1 ));
    CascadeMux I__1443 (
            .O(N__6322),
            .I(N__6319));
    InMux I__1442 (
            .O(N__6319),
            .I(N__6316));
    LocalMux I__1441 (
            .O(N__6316),
            .I(N__6313));
    IoSpan4Mux I__1440 (
            .O(N__6313),
            .I(N__6310));
    Odrv4 I__1439 (
            .O(N__6310),
            .I(A_c_3));
    InMux I__1438 (
            .O(N__6307),
            .I(N__6299));
    InMux I__1437 (
            .O(N__6306),
            .I(N__6299));
    InMux I__1436 (
            .O(N__6305),
            .I(N__6292));
    InMux I__1435 (
            .O(N__6304),
            .I(N__6292));
    LocalMux I__1434 (
            .O(N__6299),
            .I(N__6285));
    InMux I__1433 (
            .O(N__6298),
            .I(N__6280));
    InMux I__1432 (
            .O(N__6297),
            .I(N__6280));
    LocalMux I__1431 (
            .O(N__6292),
            .I(N__6277));
    InMux I__1430 (
            .O(N__6291),
            .I(N__6272));
    InMux I__1429 (
            .O(N__6290),
            .I(N__6272));
    InMux I__1428 (
            .O(N__6289),
            .I(N__6269));
    InMux I__1427 (
            .O(N__6288),
            .I(N__6266));
    Span4Mux_h I__1426 (
            .O(N__6285),
            .I(N__6257));
    LocalMux I__1425 (
            .O(N__6280),
            .I(N__6257));
    Span4Mux_h I__1424 (
            .O(N__6277),
            .I(N__6257));
    LocalMux I__1423 (
            .O(N__6272),
            .I(N__6257));
    LocalMux I__1422 (
            .O(N__6269),
            .I(N__6253));
    LocalMux I__1421 (
            .O(N__6266),
            .I(N__6250));
    Span4Mux_v I__1420 (
            .O(N__6257),
            .I(N__6246));
    InMux I__1419 (
            .O(N__6256),
            .I(N__6243));
    Span4Mux_s3_h I__1418 (
            .O(N__6253),
            .I(N__6238));
    Span4Mux_h I__1417 (
            .O(N__6250),
            .I(N__6238));
    InMux I__1416 (
            .O(N__6249),
            .I(N__6235));
    Span4Mux_h I__1415 (
            .O(N__6246),
            .I(N__6232));
    LocalMux I__1414 (
            .O(N__6243),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1413 (
            .O(N__6238),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1412 (
            .O(N__6235),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1411 (
            .O(N__6232),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_0 ));
    InMux I__1410 (
            .O(N__6223),
            .I(N__6220));
    LocalMux I__1409 (
            .O(N__6220),
            .I(N__6217));
    Odrv4 I__1408 (
            .O(N__6217),
            .I(A_c_11));
    InMux I__1407 (
            .O(N__6214),
            .I(N__6211));
    LocalMux I__1406 (
            .O(N__6211),
            .I(\U400_SDRAM.MA_5_iv_0_1 ));
    IoInMux I__1405 (
            .O(N__6208),
            .I(N__6205));
    LocalMux I__1404 (
            .O(N__6205),
            .I(N__6202));
    Odrv4 I__1403 (
            .O(N__6202),
            .I(MA_c_1));
    InMux I__1402 (
            .O(N__6199),
            .I(N__6196));
    LocalMux I__1401 (
            .O(N__6196),
            .I(N__6193));
    Odrv4 I__1400 (
            .O(N__6193),
            .I(A_c_15));
    InMux I__1399 (
            .O(N__6190),
            .I(N__6187));
    LocalMux I__1398 (
            .O(N__6187),
            .I(\U400_SDRAM.MA_5_iv_0_5 ));
    IoInMux I__1397 (
            .O(N__6184),
            .I(N__6181));
    LocalMux I__1396 (
            .O(N__6181),
            .I(N__6178));
    IoSpan4Mux I__1395 (
            .O(N__6178),
            .I(N__6175));
    Span4Mux_s1_v I__1394 (
            .O(N__6175),
            .I(N__6172));
    Span4Mux_h I__1393 (
            .O(N__6172),
            .I(N__6169));
    Odrv4 I__1392 (
            .O(N__6169),
            .I(MA_c_5));
    InMux I__1391 (
            .O(N__6166),
            .I(N__6163));
    LocalMux I__1390 (
            .O(N__6163),
            .I(N__6160));
    Span4Mux_s3_v I__1389 (
            .O(N__6160),
            .I(N__6157));
    Odrv4 I__1388 (
            .O(N__6157),
            .I(A_c_5));
    CascadeMux I__1387 (
            .O(N__6154),
            .I(N__6151));
    InMux I__1386 (
            .O(N__6151),
            .I(N__6148));
    LocalMux I__1385 (
            .O(N__6148),
            .I(N__6145));
    Span4Mux_v I__1384 (
            .O(N__6145),
            .I(N__6142));
    Odrv4 I__1383 (
            .O(N__6142),
            .I(A_c_13));
    IoInMux I__1382 (
            .O(N__6139),
            .I(N__6136));
    LocalMux I__1381 (
            .O(N__6136),
            .I(N__6133));
    IoSpan4Mux I__1380 (
            .O(N__6133),
            .I(N__6130));
    Span4Mux_s3_h I__1379 (
            .O(N__6130),
            .I(N__6127));
    Span4Mux_h I__1378 (
            .O(N__6127),
            .I(N__6124));
    Odrv4 I__1377 (
            .O(N__6124),
            .I(MA_c_3));
    InMux I__1376 (
            .O(N__6121),
            .I(N__6118));
    LocalMux I__1375 (
            .O(N__6118),
            .I(N__6115));
    Span4Mux_s2_v I__1374 (
            .O(N__6115),
            .I(N__6112));
    IoSpan4Mux I__1373 (
            .O(N__6112),
            .I(N__6109));
    Odrv4 I__1372 (
            .O(N__6109),
            .I(A_c_4));
    CascadeMux I__1371 (
            .O(N__6106),
            .I(N__6103));
    InMux I__1370 (
            .O(N__6103),
            .I(N__6100));
    LocalMux I__1369 (
            .O(N__6100),
            .I(A_c_12));
    IoInMux I__1368 (
            .O(N__6097),
            .I(N__6094));
    LocalMux I__1367 (
            .O(N__6094),
            .I(MA_c_2));
    InMux I__1366 (
            .O(N__6091),
            .I(N__6088));
    LocalMux I__1365 (
            .O(N__6088),
            .I(N__6085));
    Span4Mux_s3_v I__1364 (
            .O(N__6085),
            .I(N__6082));
    Odrv4 I__1363 (
            .O(N__6082),
            .I(A_c_6));
    CascadeMux I__1362 (
            .O(N__6079),
            .I(N__6076));
    InMux I__1361 (
            .O(N__6076),
            .I(N__6073));
    LocalMux I__1360 (
            .O(N__6073),
            .I(N__6070));
    Span4Mux_h I__1359 (
            .O(N__6070),
            .I(N__6067));
    Odrv4 I__1358 (
            .O(N__6067),
            .I(A_c_14));
    IoInMux I__1357 (
            .O(N__6064),
            .I(N__6061));
    LocalMux I__1356 (
            .O(N__6061),
            .I(N__6058));
    IoSpan4Mux I__1355 (
            .O(N__6058),
            .I(N__6055));
    IoSpan4Mux I__1354 (
            .O(N__6055),
            .I(N__6052));
    Odrv4 I__1353 (
            .O(N__6052),
            .I(MA_c_4));
    InMux I__1352 (
            .O(N__6049),
            .I(N__6046));
    LocalMux I__1351 (
            .O(N__6046),
            .I(N__6043));
    Span4Mux_h I__1350 (
            .O(N__6043),
            .I(N__6040));
    Odrv4 I__1349 (
            .O(N__6040),
            .I(A_c_2));
    CascadeMux I__1348 (
            .O(N__6037),
            .I(N__6028));
    InMux I__1347 (
            .O(N__6036),
            .I(N__6020));
    InMux I__1346 (
            .O(N__6035),
            .I(N__6017));
    InMux I__1345 (
            .O(N__6034),
            .I(N__6012));
    InMux I__1344 (
            .O(N__6033),
            .I(N__6012));
    InMux I__1343 (
            .O(N__6032),
            .I(N__6007));
    InMux I__1342 (
            .O(N__6031),
            .I(N__6007));
    InMux I__1341 (
            .O(N__6028),
            .I(N__6001));
    InMux I__1340 (
            .O(N__6027),
            .I(N__6001));
    InMux I__1339 (
            .O(N__6026),
            .I(N__5996));
    InMux I__1338 (
            .O(N__6025),
            .I(N__5996));
    InMux I__1337 (
            .O(N__6024),
            .I(N__5989));
    InMux I__1336 (
            .O(N__6023),
            .I(N__5989));
    LocalMux I__1335 (
            .O(N__6020),
            .I(N__5980));
    LocalMux I__1334 (
            .O(N__6017),
            .I(N__5980));
    LocalMux I__1333 (
            .O(N__6012),
            .I(N__5980));
    LocalMux I__1332 (
            .O(N__6007),
            .I(N__5980));
    InMux I__1331 (
            .O(N__6006),
            .I(N__5975));
    LocalMux I__1330 (
            .O(N__6001),
            .I(N__5972));
    LocalMux I__1329 (
            .O(N__5996),
            .I(N__5969));
    InMux I__1328 (
            .O(N__5995),
            .I(N__5966));
    InMux I__1327 (
            .O(N__5994),
            .I(N__5962));
    LocalMux I__1326 (
            .O(N__5989),
            .I(N__5959));
    Span4Mux_s3_v I__1325 (
            .O(N__5980),
            .I(N__5956));
    InMux I__1324 (
            .O(N__5979),
            .I(N__5953));
    InMux I__1323 (
            .O(N__5978),
            .I(N__5950));
    LocalMux I__1322 (
            .O(N__5975),
            .I(N__5947));
    Span4Mux_s3_v I__1321 (
            .O(N__5972),
            .I(N__5942));
    Span4Mux_s3_v I__1320 (
            .O(N__5969),
            .I(N__5942));
    LocalMux I__1319 (
            .O(N__5966),
            .I(N__5938));
    InMux I__1318 (
            .O(N__5965),
            .I(N__5935));
    LocalMux I__1317 (
            .O(N__5962),
            .I(N__5928));
    Span4Mux_s3_v I__1316 (
            .O(N__5959),
            .I(N__5928));
    Span4Mux_h I__1315 (
            .O(N__5956),
            .I(N__5928));
    LocalMux I__1314 (
            .O(N__5953),
            .I(N__5925));
    LocalMux I__1313 (
            .O(N__5950),
            .I(N__5918));
    Span4Mux_s3_v I__1312 (
            .O(N__5947),
            .I(N__5918));
    Span4Mux_h I__1311 (
            .O(N__5942),
            .I(N__5918));
    InMux I__1310 (
            .O(N__5941),
            .I(N__5915));
    Span4Mux_v I__1309 (
            .O(N__5938),
            .I(N__5912));
    LocalMux I__1308 (
            .O(N__5935),
            .I(N__5907));
    Span4Mux_v I__1307 (
            .O(N__5928),
            .I(N__5907));
    Span4Mux_h I__1306 (
            .O(N__5925),
            .I(N__5902));
    Span4Mux_v I__1305 (
            .O(N__5918),
            .I(N__5902));
    LocalMux I__1304 (
            .O(N__5915),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1303 (
            .O(N__5912),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1302 (
            .O(N__5907),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1301 (
            .O(N__5902),
            .I(\U400_SDRAM.SDRAM_CMDZ0Z_2 ));
    InMux I__1300 (
            .O(N__5893),
            .I(N__5889));
    InMux I__1299 (
            .O(N__5892),
            .I(N__5883));
    LocalMux I__1298 (
            .O(N__5889),
            .I(N__5880));
    InMux I__1297 (
            .O(N__5888),
            .I(N__5875));
    InMux I__1296 (
            .O(N__5887),
            .I(N__5875));
    InMux I__1295 (
            .O(N__5886),
            .I(N__5872));
    LocalMux I__1294 (
            .O(N__5883),
            .I(U400_SDRAM_BURST));
    Odrv4 I__1293 (
            .O(N__5880),
            .I(U400_SDRAM_BURST));
    LocalMux I__1292 (
            .O(N__5875),
            .I(U400_SDRAM_BURST));
    LocalMux I__1291 (
            .O(N__5872),
            .I(U400_SDRAM_BURST));
    InMux I__1290 (
            .O(N__5863),
            .I(N__5860));
    LocalMux I__1289 (
            .O(N__5860),
            .I(\U400_ADDRESS_DECODE.N_114_0 ));
    InMux I__1288 (
            .O(N__5857),
            .I(N__5853));
    InMux I__1287 (
            .O(N__5856),
            .I(N__5848));
    LocalMux I__1286 (
            .O(N__5853),
            .I(N__5843));
    InMux I__1285 (
            .O(N__5852),
            .I(N__5838));
    InMux I__1284 (
            .O(N__5851),
            .I(N__5838));
    LocalMux I__1283 (
            .O(N__5848),
            .I(N__5835));
    InMux I__1282 (
            .O(N__5847),
            .I(N__5830));
    InMux I__1281 (
            .O(N__5846),
            .I(N__5830));
    Span12Mux_s6_h I__1280 (
            .O(N__5843),
            .I(N__5827));
    LocalMux I__1279 (
            .O(N__5838),
            .I(N__5824));
    Span4Mux_h I__1278 (
            .O(N__5835),
            .I(N__5821));
    LocalMux I__1277 (
            .O(N__5830),
            .I(N__5818));
    Odrv12 I__1276 (
            .O(N__5827),
            .I(N_65_0));
    Odrv4 I__1275 (
            .O(N__5824),
            .I(N_65_0));
    Odrv4 I__1274 (
            .O(N__5821),
            .I(N_65_0));
    Odrv4 I__1273 (
            .O(N__5818),
            .I(N_65_0));
    InMux I__1272 (
            .O(N__5809),
            .I(N__5797));
    InMux I__1271 (
            .O(N__5808),
            .I(N__5792));
    InMux I__1270 (
            .O(N__5807),
            .I(N__5792));
    InMux I__1269 (
            .O(N__5806),
            .I(N__5789));
    CascadeMux I__1268 (
            .O(N__5805),
            .I(N__5779));
    InMux I__1267 (
            .O(N__5804),
            .I(N__5776));
    InMux I__1266 (
            .O(N__5803),
            .I(N__5773));
    InMux I__1265 (
            .O(N__5802),
            .I(N__5768));
    InMux I__1264 (
            .O(N__5801),
            .I(N__5768));
    InMux I__1263 (
            .O(N__5800),
            .I(N__5765));
    LocalMux I__1262 (
            .O(N__5797),
            .I(N__5758));
    LocalMux I__1261 (
            .O(N__5792),
            .I(N__5758));
    LocalMux I__1260 (
            .O(N__5789),
            .I(N__5758));
    CascadeMux I__1259 (
            .O(N__5788),
            .I(N__5755));
    InMux I__1258 (
            .O(N__5787),
            .I(N__5752));
    InMux I__1257 (
            .O(N__5786),
            .I(N__5747));
    InMux I__1256 (
            .O(N__5785),
            .I(N__5747));
    InMux I__1255 (
            .O(N__5784),
            .I(N__5742));
    InMux I__1254 (
            .O(N__5783),
            .I(N__5742));
    InMux I__1253 (
            .O(N__5782),
            .I(N__5739));
    InMux I__1252 (
            .O(N__5779),
            .I(N__5736));
    LocalMux I__1251 (
            .O(N__5776),
            .I(N__5733));
    LocalMux I__1250 (
            .O(N__5773),
            .I(N__5728));
    LocalMux I__1249 (
            .O(N__5768),
            .I(N__5728));
    LocalMux I__1248 (
            .O(N__5765),
            .I(N__5720));
    Span4Mux_v I__1247 (
            .O(N__5758),
            .I(N__5720));
    InMux I__1246 (
            .O(N__5755),
            .I(N__5717));
    LocalMux I__1245 (
            .O(N__5752),
            .I(N__5714));
    LocalMux I__1244 (
            .O(N__5747),
            .I(N__5711));
    LocalMux I__1243 (
            .O(N__5742),
            .I(N__5704));
    LocalMux I__1242 (
            .O(N__5739),
            .I(N__5704));
    LocalMux I__1241 (
            .O(N__5736),
            .I(N__5704));
    Span4Mux_v I__1240 (
            .O(N__5733),
            .I(N__5699));
    Span4Mux_v I__1239 (
            .O(N__5728),
            .I(N__5699));
    InMux I__1238 (
            .O(N__5727),
            .I(N__5696));
    InMux I__1237 (
            .O(N__5726),
            .I(N__5691));
    InMux I__1236 (
            .O(N__5725),
            .I(N__5691));
    Span4Mux_h I__1235 (
            .O(N__5720),
            .I(N__5688));
    LocalMux I__1234 (
            .O(N__5717),
            .I(N__5677));
    Span4Mux_v I__1233 (
            .O(N__5714),
            .I(N__5677));
    Span4Mux_v I__1232 (
            .O(N__5711),
            .I(N__5677));
    Span4Mux_v I__1231 (
            .O(N__5704),
            .I(N__5677));
    Span4Mux_h I__1230 (
            .O(N__5699),
            .I(N__5677));
    LocalMux I__1229 (
            .O(N__5696),
            .I(U400_SDRAM_SDRAM_CONFIGURED));
    LocalMux I__1228 (
            .O(N__5691),
            .I(U400_SDRAM_SDRAM_CONFIGURED));
    Odrv4 I__1227 (
            .O(N__5688),
            .I(U400_SDRAM_SDRAM_CONFIGURED));
    Odrv4 I__1226 (
            .O(N__5677),
            .I(U400_SDRAM_SDRAM_CONFIGURED));
    IoInMux I__1225 (
            .O(N__5668),
            .I(N__5665));
    LocalMux I__1224 (
            .O(N__5665),
            .I(N__5662));
    Odrv4 I__1223 (
            .O(N__5662),
            .I(N_129_0));
    IoInMux I__1222 (
            .O(N__5659),
            .I(N__5656));
    LocalMux I__1221 (
            .O(N__5656),
            .I(N__5653));
    Odrv12 I__1220 (
            .O(N__5653),
            .I(N_127_0));
    InMux I__1219 (
            .O(N__5650),
            .I(N__5641));
    InMux I__1218 (
            .O(N__5649),
            .I(N__5641));
    InMux I__1217 (
            .O(N__5648),
            .I(N__5641));
    LocalMux I__1216 (
            .O(N__5641),
            .I(N__5638));
    Span4Mux_v I__1215 (
            .O(N__5638),
            .I(N__5635));
    Span4Mux_v I__1214 (
            .O(N__5635),
            .I(N__5631));
    InMux I__1213 (
            .O(N__5634),
            .I(N__5628));
    Span4Mux_v I__1212 (
            .O(N__5631),
            .I(N__5625));
    LocalMux I__1211 (
            .O(N__5628),
            .I(N__5622));
    Sp12to4 I__1210 (
            .O(N__5625),
            .I(N__5617));
    Span12Mux_v I__1209 (
            .O(N__5622),
            .I(N__5617));
    Odrv12 I__1208 (
            .O(N__5617),
            .I(A_c_1));
    IoInMux I__1207 (
            .O(N__5614),
            .I(N__5611));
    LocalMux I__1206 (
            .O(N__5611),
            .I(N__5608));
    Odrv4 I__1205 (
            .O(N__5608),
            .I(N_128_0));
    CascadeMux I__1204 (
            .O(N__5605),
            .I(N__5600));
    CascadeMux I__1203 (
            .O(N__5604),
            .I(N__5597));
    InMux I__1202 (
            .O(N__5603),
            .I(N__5593));
    InMux I__1201 (
            .O(N__5600),
            .I(N__5586));
    InMux I__1200 (
            .O(N__5597),
            .I(N__5586));
    InMux I__1199 (
            .O(N__5596),
            .I(N__5586));
    LocalMux I__1198 (
            .O(N__5593),
            .I(\U400_ADDRESS_DECODE.N_122_0 ));
    LocalMux I__1197 (
            .O(N__5586),
            .I(\U400_ADDRESS_DECODE.N_122_0 ));
    CascadeMux I__1196 (
            .O(N__5581),
            .I(N__5578));
    InMux I__1195 (
            .O(N__5578),
            .I(N__5573));
    InMux I__1194 (
            .O(N__5577),
            .I(N__5568));
    InMux I__1193 (
            .O(N__5576),
            .I(N__5568));
    LocalMux I__1192 (
            .O(N__5573),
            .I(N__5565));
    LocalMux I__1191 (
            .O(N__5568),
            .I(N__5561));
    Span4Mux_v I__1190 (
            .O(N__5565),
            .I(N__5558));
    InMux I__1189 (
            .O(N__5564),
            .I(N__5555));
    Span4Mux_v I__1188 (
            .O(N__5561),
            .I(N__5552));
    Sp12to4 I__1187 (
            .O(N__5558),
            .I(N__5547));
    LocalMux I__1186 (
            .O(N__5555),
            .I(N__5547));
    Odrv4 I__1185 (
            .O(N__5552),
            .I(SIZ_c_0));
    Odrv12 I__1184 (
            .O(N__5547),
            .I(SIZ_c_0));
    InMux I__1183 (
            .O(N__5542),
            .I(N__5538));
    InMux I__1182 (
            .O(N__5541),
            .I(N__5535));
    LocalMux I__1181 (
            .O(N__5538),
            .I(N__5531));
    LocalMux I__1180 (
            .O(N__5535),
            .I(N__5528));
    InMux I__1179 (
            .O(N__5534),
            .I(N__5525));
    Span4Mux_h I__1178 (
            .O(N__5531),
            .I(N__5520));
    Span4Mux_v I__1177 (
            .O(N__5528),
            .I(N__5520));
    LocalMux I__1176 (
            .O(N__5525),
            .I(N__5517));
    Span4Mux_v I__1175 (
            .O(N__5520),
            .I(N__5514));
    Sp12to4 I__1174 (
            .O(N__5517),
            .I(N__5511));
    Span4Mux_v I__1173 (
            .O(N__5514),
            .I(N__5508));
    Span12Mux_v I__1172 (
            .O(N__5511),
            .I(N__5505));
    Span4Mux_h I__1171 (
            .O(N__5508),
            .I(N__5502));
    Odrv12 I__1170 (
            .O(N__5505),
            .I(A_c_0));
    Odrv4 I__1169 (
            .O(N__5502),
            .I(A_c_0));
    CascadeMux I__1168 (
            .O(N__5497),
            .I(N__5493));
    InMux I__1167 (
            .O(N__5496),
            .I(N__5490));
    InMux I__1166 (
            .O(N__5493),
            .I(N__5486));
    LocalMux I__1165 (
            .O(N__5490),
            .I(N__5483));
    InMux I__1164 (
            .O(N__5489),
            .I(N__5480));
    LocalMux I__1163 (
            .O(N__5486),
            .I(\U400_ADDRESS_DECODE.N_4_0 ));
    Odrv12 I__1162 (
            .O(N__5483),
            .I(\U400_ADDRESS_DECODE.N_4_0 ));
    LocalMux I__1161 (
            .O(N__5480),
            .I(\U400_ADDRESS_DECODE.N_4_0 ));
    InMux I__1160 (
            .O(N__5473),
            .I(N__5470));
    LocalMux I__1159 (
            .O(N__5470),
            .I(N__5466));
    InMux I__1158 (
            .O(N__5469),
            .I(N__5463));
    Span4Mux_v I__1157 (
            .O(N__5466),
            .I(N__5456));
    LocalMux I__1156 (
            .O(N__5463),
            .I(N__5456));
    InMux I__1155 (
            .O(N__5462),
            .I(N__5451));
    InMux I__1154 (
            .O(N__5461),
            .I(N__5451));
    Span4Mux_v I__1153 (
            .O(N__5456),
            .I(N__5448));
    LocalMux I__1152 (
            .O(N__5451),
            .I(N__5445));
    Span4Mux_h I__1151 (
            .O(N__5448),
            .I(N__5442));
    Span4Mux_v I__1150 (
            .O(N__5445),
            .I(N__5439));
    Odrv4 I__1149 (
            .O(N__5442),
            .I(SIZ_c_1));
    Odrv4 I__1148 (
            .O(N__5439),
            .I(SIZ_c_1));
    InMux I__1147 (
            .O(N__5434),
            .I(N__5428));
    InMux I__1146 (
            .O(N__5433),
            .I(N__5428));
    LocalMux I__1145 (
            .O(N__5428),
            .I(\U400_ADDRESS_DECODE.N_186_mux ));
    InMux I__1144 (
            .O(N__5425),
            .I(N__5422));
    LocalMux I__1143 (
            .O(N__5422),
            .I(\U400_ADDRESS_DECODE.N_146_0 ));
    CascadeMux I__1142 (
            .O(N__5419),
            .I(N__5415));
    CascadeMux I__1141 (
            .O(N__5418),
            .I(N__5412));
    InMux I__1140 (
            .O(N__5415),
            .I(N__5407));
    InMux I__1139 (
            .O(N__5412),
            .I(N__5407));
    LocalMux I__1138 (
            .O(N__5407),
            .I(N__5404));
    Span4Mux_h I__1137 (
            .O(N__5404),
            .I(N__5401));
    Span4Mux_v I__1136 (
            .O(N__5401),
            .I(N__5397));
    InMux I__1135 (
            .O(N__5400),
            .I(N__5394));
    Odrv4 I__1134 (
            .O(N__5397),
            .I(N_14_i));
    LocalMux I__1133 (
            .O(N__5394),
            .I(N_14_i));
    CascadeMux I__1132 (
            .O(N__5389),
            .I(\U400_ADDRESS_DECODE.N_147_0_cascade_ ));
    InMux I__1131 (
            .O(N__5386),
            .I(N__5383));
    LocalMux I__1130 (
            .O(N__5383),
            .I(\U400_ADDRESS_DECODE.N_136_0 ));
    InMux I__1129 (
            .O(N__5380),
            .I(N__5377));
    LocalMux I__1128 (
            .O(N__5377),
            .I(N_43));
    InMux I__1127 (
            .O(N__5374),
            .I(N__5371));
    LocalMux I__1126 (
            .O(N__5371),
            .I(N__5368));
    Span4Mux_h I__1125 (
            .O(N__5368),
            .I(N__5365));
    Sp12to4 I__1124 (
            .O(N__5365),
            .I(N__5362));
    Span12Mux_v I__1123 (
            .O(N__5362),
            .I(N__5359));
    Odrv12 I__1122 (
            .O(N__5359),
            .I(A_c_20));
    IoInMux I__1121 (
            .O(N__5356),
            .I(N__5353));
    LocalMux I__1120 (
            .O(N__5353),
            .I(N__5350));
    Span4Mux_s0_v I__1119 (
            .O(N__5350),
            .I(N__5347));
    Odrv4 I__1118 (
            .O(N__5347),
            .I(MA_c_10));
    CascadeMux I__1117 (
            .O(N__5344),
            .I(N__5341));
    InMux I__1116 (
            .O(N__5341),
            .I(N__5338));
    LocalMux I__1115 (
            .O(N__5338),
            .I(N__5335));
    Span12Mux_s11_v I__1114 (
            .O(N__5335),
            .I(N__5332));
    Odrv12 I__1113 (
            .O(N__5332),
            .I(A_c_25));
    IoInMux I__1112 (
            .O(N__5329),
            .I(N__5326));
    LocalMux I__1111 (
            .O(N__5326),
            .I(N__5323));
    Odrv4 I__1110 (
            .O(N__5323),
            .I(MA_c_11));
    CascadeMux I__1109 (
            .O(N__5320),
            .I(\U400_ADDRESS_DECODE.N_4_0_cascade_ ));
    IoInMux I__1108 (
            .O(N__5317),
            .I(N__5314));
    LocalMux I__1107 (
            .O(N__5314),
            .I(N__5311));
    Span12Mux_s3_v I__1106 (
            .O(N__5311),
            .I(N__5308));
    Odrv12 I__1105 (
            .O(N__5308),
            .I(N_124_0));
    InMux I__1104 (
            .O(N__5305),
            .I(N__5302));
    LocalMux I__1103 (
            .O(N__5302),
            .I(\U400_SDRAM.N_252_0_0 ));
    InMux I__1102 (
            .O(N__5299),
            .I(N__5296));
    LocalMux I__1101 (
            .O(N__5296),
            .I(\U400_SDRAM.N_252_0_0_en ));
    InMux I__1100 (
            .O(N__5293),
            .I(N__5289));
    InMux I__1099 (
            .O(N__5292),
            .I(N__5286));
    LocalMux I__1098 (
            .O(N__5289),
            .I(N_174));
    LocalMux I__1097 (
            .O(N__5286),
            .I(N_174));
    InMux I__1096 (
            .O(N__5281),
            .I(N__5278));
    LocalMux I__1095 (
            .O(N__5278),
            .I(U400_SDRAM_TA_OUT_5_0));
    InMux I__1094 (
            .O(N__5275),
            .I(N__5272));
    LocalMux I__1093 (
            .O(N__5272),
            .I(U400_SDRAM_N_252_0));
    IoInMux I__1092 (
            .O(N__5269),
            .I(N__5266));
    LocalMux I__1091 (
            .O(N__5266),
            .I(N__5262));
    CascadeMux I__1090 (
            .O(N__5265),
            .I(N__5259));
    Span4Mux_s3_h I__1089 (
            .O(N__5262),
            .I(N__5256));
    InMux I__1088 (
            .O(N__5259),
            .I(N__5253));
    Odrv4 I__1087 (
            .O(N__5256),
            .I(TA_OUT));
    LocalMux I__1086 (
            .O(N__5253),
            .I(TA_OUT));
    ClkMux I__1085 (
            .O(N__5248),
            .I(N__5167));
    ClkMux I__1084 (
            .O(N__5247),
            .I(N__5167));
    ClkMux I__1083 (
            .O(N__5246),
            .I(N__5167));
    ClkMux I__1082 (
            .O(N__5245),
            .I(N__5167));
    ClkMux I__1081 (
            .O(N__5244),
            .I(N__5167));
    ClkMux I__1080 (
            .O(N__5243),
            .I(N__5167));
    ClkMux I__1079 (
            .O(N__5242),
            .I(N__5167));
    ClkMux I__1078 (
            .O(N__5241),
            .I(N__5167));
    ClkMux I__1077 (
            .O(N__5240),
            .I(N__5167));
    ClkMux I__1076 (
            .O(N__5239),
            .I(N__5167));
    ClkMux I__1075 (
            .O(N__5238),
            .I(N__5167));
    ClkMux I__1074 (
            .O(N__5237),
            .I(N__5167));
    ClkMux I__1073 (
            .O(N__5236),
            .I(N__5167));
    ClkMux I__1072 (
            .O(N__5235),
            .I(N__5167));
    ClkMux I__1071 (
            .O(N__5234),
            .I(N__5167));
    ClkMux I__1070 (
            .O(N__5233),
            .I(N__5167));
    ClkMux I__1069 (
            .O(N__5232),
            .I(N__5167));
    ClkMux I__1068 (
            .O(N__5231),
            .I(N__5167));
    ClkMux I__1067 (
            .O(N__5230),
            .I(N__5167));
    ClkMux I__1066 (
            .O(N__5229),
            .I(N__5167));
    ClkMux I__1065 (
            .O(N__5228),
            .I(N__5167));
    ClkMux I__1064 (
            .O(N__5227),
            .I(N__5167));
    ClkMux I__1063 (
            .O(N__5226),
            .I(N__5167));
    ClkMux I__1062 (
            .O(N__5225),
            .I(N__5167));
    ClkMux I__1061 (
            .O(N__5224),
            .I(N__5167));
    ClkMux I__1060 (
            .O(N__5223),
            .I(N__5167));
    ClkMux I__1059 (
            .O(N__5222),
            .I(N__5167));
    GlobalMux I__1058 (
            .O(N__5167),
            .I(N__5164));
    gio2CtrlBuf I__1057 (
            .O(N__5164),
            .I(CLK40_c_g));
    InMux I__1056 (
            .O(N__5161),
            .I(N__5155));
    InMux I__1055 (
            .O(N__5160),
            .I(N__5155));
    LocalMux I__1054 (
            .O(N__5155),
            .I(U400_SDRAM_TA_COUNTER_5));
    CascadeMux I__1053 (
            .O(N__5152),
            .I(\U400_SDRAM.N_252_0_0_cascade_ ));
    CascadeMux I__1052 (
            .O(N__5149),
            .I(N__5145));
    InMux I__1051 (
            .O(N__5148),
            .I(N__5137));
    InMux I__1050 (
            .O(N__5145),
            .I(N__5137));
    InMux I__1049 (
            .O(N__5144),
            .I(N__5137));
    LocalMux I__1048 (
            .O(N__5137),
            .I(U400_SDRAM_TA_COUNTER_2));
    InMux I__1047 (
            .O(N__5134),
            .I(N__5130));
    InMux I__1046 (
            .O(N__5133),
            .I(N__5127));
    LocalMux I__1045 (
            .O(N__5130),
            .I(U400_SDRAM_TA_COUNTER_3));
    LocalMux I__1044 (
            .O(N__5127),
            .I(U400_SDRAM_TA_COUNTER_3));
    CascadeMux I__1043 (
            .O(N__5122),
            .I(N__5119));
    InMux I__1042 (
            .O(N__5119),
            .I(N__5116));
    LocalMux I__1041 (
            .O(N__5116),
            .I(N__5113));
    Span4Mux_v I__1040 (
            .O(N__5113),
            .I(N__5110));
    Span4Mux_h I__1039 (
            .O(N__5110),
            .I(N__5107));
    Odrv4 I__1038 (
            .O(N__5107),
            .I(A_c_22));
    IoInMux I__1037 (
            .O(N__5104),
            .I(N__5101));
    LocalMux I__1036 (
            .O(N__5101),
            .I(N__5098));
    Span4Mux_s2_h I__1035 (
            .O(N__5098),
            .I(N__5095));
    Span4Mux_h I__1034 (
            .O(N__5095),
            .I(N__5092));
    Span4Mux_v I__1033 (
            .O(N__5092),
            .I(N__5088));
    InMux I__1032 (
            .O(N__5091),
            .I(N__5085));
    Odrv4 I__1031 (
            .O(N__5088),
            .I(BANK1_c));
    LocalMux I__1030 (
            .O(N__5085),
            .I(BANK1_c));
    CascadeMux I__1029 (
            .O(N__5080),
            .I(N__5077));
    InMux I__1028 (
            .O(N__5077),
            .I(N__5074));
    LocalMux I__1027 (
            .O(N__5074),
            .I(N__5071));
    Span4Mux_v I__1026 (
            .O(N__5071),
            .I(N__5068));
    Sp12to4 I__1025 (
            .O(N__5068),
            .I(N__5065));
    Odrv12 I__1024 (
            .O(N__5065),
            .I(A_c_21));
    InMux I__1023 (
            .O(N__5062),
            .I(N__5056));
    InMux I__1022 (
            .O(N__5061),
            .I(N__5056));
    LocalMux I__1021 (
            .O(N__5056),
            .I(U400_SDRAM_un1_SDRAM_COUNTER59_2_0));
    IoInMux I__1020 (
            .O(N__5053),
            .I(N__5050));
    LocalMux I__1019 (
            .O(N__5050),
            .I(N__5047));
    Span4Mux_s2_h I__1018 (
            .O(N__5047),
            .I(N__5044));
    Span4Mux_h I__1017 (
            .O(N__5044),
            .I(N__5041));
    Span4Mux_v I__1016 (
            .O(N__5041),
            .I(N__5037));
    InMux I__1015 (
            .O(N__5040),
            .I(N__5034));
    Odrv4 I__1014 (
            .O(N__5037),
            .I(BANK0_c));
    LocalMux I__1013 (
            .O(N__5034),
            .I(BANK0_c));
    InMux I__1012 (
            .O(N__5029),
            .I(N__5026));
    LocalMux I__1011 (
            .O(N__5026),
            .I(N__5022));
    InMux I__1010 (
            .O(N__5025),
            .I(N__5019));
    Odrv4 I__1009 (
            .O(N__5022),
            .I(U400_SDRAM_SDRAM_CMD_1_sqmuxa_1));
    LocalMux I__1008 (
            .O(N__5019),
            .I(U400_SDRAM_SDRAM_CMD_1_sqmuxa_1));
    InMux I__1007 (
            .O(N__5014),
            .I(N__5007));
    InMux I__1006 (
            .O(N__5013),
            .I(N__5004));
    CascadeMux I__1005 (
            .O(N__5012),
            .I(N__4997));
    CascadeMux I__1004 (
            .O(N__5011),
            .I(N__4993));
    CascadeMux I__1003 (
            .O(N__5010),
            .I(N__4990));
    LocalMux I__1002 (
            .O(N__5007),
            .I(N__4978));
    LocalMux I__1001 (
            .O(N__5004),
            .I(N__4978));
    InMux I__1000 (
            .O(N__5003),
            .I(N__4975));
    InMux I__999 (
            .O(N__5002),
            .I(N__4972));
    InMux I__998 (
            .O(N__5001),
            .I(N__4967));
    InMux I__997 (
            .O(N__5000),
            .I(N__4967));
    InMux I__996 (
            .O(N__4997),
            .I(N__4962));
    InMux I__995 (
            .O(N__4996),
            .I(N__4962));
    InMux I__994 (
            .O(N__4993),
            .I(N__4959));
    InMux I__993 (
            .O(N__4990),
            .I(N__4954));
    InMux I__992 (
            .O(N__4989),
            .I(N__4954));
    CascadeMux I__991 (
            .O(N__4988),
            .I(N__4950));
    CascadeMux I__990 (
            .O(N__4987),
            .I(N__4944));
    InMux I__989 (
            .O(N__4986),
            .I(N__4939));
    InMux I__988 (
            .O(N__4985),
            .I(N__4939));
    CascadeMux I__987 (
            .O(N__4984),
            .I(N__4936));
    InMux I__986 (
            .O(N__4983),
            .I(N__4933));
    Span4Mux_h I__985 (
            .O(N__4978),
            .I(N__4924));
    LocalMux I__984 (
            .O(N__4975),
            .I(N__4924));
    LocalMux I__983 (
            .O(N__4972),
            .I(N__4924));
    LocalMux I__982 (
            .O(N__4967),
            .I(N__4924));
    LocalMux I__981 (
            .O(N__4962),
            .I(N__4919));
    LocalMux I__980 (
            .O(N__4959),
            .I(N__4914));
    LocalMux I__979 (
            .O(N__4954),
            .I(N__4914));
    InMux I__978 (
            .O(N__4953),
            .I(N__4909));
    InMux I__977 (
            .O(N__4950),
            .I(N__4909));
    InMux I__976 (
            .O(N__4949),
            .I(N__4904));
    InMux I__975 (
            .O(N__4948),
            .I(N__4904));
    InMux I__974 (
            .O(N__4947),
            .I(N__4899));
    InMux I__973 (
            .O(N__4944),
            .I(N__4899));
    LocalMux I__972 (
            .O(N__4939),
            .I(N__4896));
    InMux I__971 (
            .O(N__4936),
            .I(N__4893));
    LocalMux I__970 (
            .O(N__4933),
            .I(N__4888));
    Span4Mux_v I__969 (
            .O(N__4924),
            .I(N__4888));
    InMux I__968 (
            .O(N__4923),
            .I(N__4885));
    InMux I__967 (
            .O(N__4922),
            .I(N__4882));
    Span4Mux_h I__966 (
            .O(N__4919),
            .I(N__4871));
    Span4Mux_h I__965 (
            .O(N__4914),
            .I(N__4871));
    LocalMux I__964 (
            .O(N__4909),
            .I(N__4871));
    LocalMux I__963 (
            .O(N__4904),
            .I(N__4871));
    LocalMux I__962 (
            .O(N__4899),
            .I(N__4871));
    Odrv12 I__961 (
            .O(N__4896),
            .I(U400_SDRAM_SDRAM_COUNTER_2));
    LocalMux I__960 (
            .O(N__4893),
            .I(U400_SDRAM_SDRAM_COUNTER_2));
    Odrv4 I__959 (
            .O(N__4888),
            .I(U400_SDRAM_SDRAM_COUNTER_2));
    LocalMux I__958 (
            .O(N__4885),
            .I(U400_SDRAM_SDRAM_COUNTER_2));
    LocalMux I__957 (
            .O(N__4882),
            .I(U400_SDRAM_SDRAM_COUNTER_2));
    Odrv4 I__956 (
            .O(N__4871),
            .I(U400_SDRAM_SDRAM_COUNTER_2));
    InMux I__955 (
            .O(N__4858),
            .I(N__4850));
    InMux I__954 (
            .O(N__4857),
            .I(N__4844));
    InMux I__953 (
            .O(N__4856),
            .I(N__4837));
    InMux I__952 (
            .O(N__4855),
            .I(N__4837));
    InMux I__951 (
            .O(N__4854),
            .I(N__4837));
    InMux I__950 (
            .O(N__4853),
            .I(N__4834));
    LocalMux I__949 (
            .O(N__4850),
            .I(N__4828));
    InMux I__948 (
            .O(N__4849),
            .I(N__4821));
    InMux I__947 (
            .O(N__4848),
            .I(N__4821));
    InMux I__946 (
            .O(N__4847),
            .I(N__4821));
    LocalMux I__945 (
            .O(N__4844),
            .I(N__4815));
    LocalMux I__944 (
            .O(N__4837),
            .I(N__4810));
    LocalMux I__943 (
            .O(N__4834),
            .I(N__4810));
    InMux I__942 (
            .O(N__4833),
            .I(N__4807));
    InMux I__941 (
            .O(N__4832),
            .I(N__4802));
    InMux I__940 (
            .O(N__4831),
            .I(N__4802));
    Span4Mux_v I__939 (
            .O(N__4828),
            .I(N__4792));
    LocalMux I__938 (
            .O(N__4821),
            .I(N__4789));
    InMux I__937 (
            .O(N__4820),
            .I(N__4786));
    InMux I__936 (
            .O(N__4819),
            .I(N__4781));
    InMux I__935 (
            .O(N__4818),
            .I(N__4781));
    Span4Mux_h I__934 (
            .O(N__4815),
            .I(N__4772));
    Span4Mux_v I__933 (
            .O(N__4810),
            .I(N__4772));
    LocalMux I__932 (
            .O(N__4807),
            .I(N__4772));
    LocalMux I__931 (
            .O(N__4802),
            .I(N__4772));
    InMux I__930 (
            .O(N__4801),
            .I(N__4767));
    InMux I__929 (
            .O(N__4800),
            .I(N__4767));
    InMux I__928 (
            .O(N__4799),
            .I(N__4762));
    InMux I__927 (
            .O(N__4798),
            .I(N__4762));
    InMux I__926 (
            .O(N__4797),
            .I(N__4755));
    InMux I__925 (
            .O(N__4796),
            .I(N__4755));
    InMux I__924 (
            .O(N__4795),
            .I(N__4755));
    Odrv4 I__923 (
            .O(N__4792),
            .I(N_60));
    Odrv4 I__922 (
            .O(N__4789),
            .I(N_60));
    LocalMux I__921 (
            .O(N__4786),
            .I(N_60));
    LocalMux I__920 (
            .O(N__4781),
            .I(N_60));
    Odrv4 I__919 (
            .O(N__4772),
            .I(N_60));
    LocalMux I__918 (
            .O(N__4767),
            .I(N_60));
    LocalMux I__917 (
            .O(N__4762),
            .I(N_60));
    LocalMux I__916 (
            .O(N__4755),
            .I(N_60));
    InMux I__915 (
            .O(N__4738),
            .I(N__4735));
    LocalMux I__914 (
            .O(N__4735),
            .I(\U400_ADDRESS_DECODE.m145_nsZ0Z_1 ));
    InMux I__913 (
            .O(N__4732),
            .I(N__4728));
    InMux I__912 (
            .O(N__4731),
            .I(N__4725));
    LocalMux I__911 (
            .O(N__4728),
            .I(N__4716));
    LocalMux I__910 (
            .O(N__4725),
            .I(N__4713));
    InMux I__909 (
            .O(N__4724),
            .I(N__4708));
    InMux I__908 (
            .O(N__4723),
            .I(N__4708));
    InMux I__907 (
            .O(N__4722),
            .I(N__4699));
    InMux I__906 (
            .O(N__4721),
            .I(N__4699));
    InMux I__905 (
            .O(N__4720),
            .I(N__4699));
    InMux I__904 (
            .O(N__4719),
            .I(N__4699));
    Span4Mux_h I__903 (
            .O(N__4716),
            .I(N__4696));
    Odrv4 I__902 (
            .O(N__4713),
            .I(N_100_0_i));
    LocalMux I__901 (
            .O(N__4708),
            .I(N_100_0_i));
    LocalMux I__900 (
            .O(N__4699),
            .I(N_100_0_i));
    Odrv4 I__899 (
            .O(N__4696),
            .I(N_100_0_i));
    IoInMux I__898 (
            .O(N__4687),
            .I(N__4684));
    LocalMux I__897 (
            .O(N__4684),
            .I(N__4681));
    IoSpan4Mux I__896 (
            .O(N__4681),
            .I(N__4678));
    Span4Mux_s1_h I__895 (
            .O(N__4678),
            .I(N__4674));
    CascadeMux I__894 (
            .O(N__4677),
            .I(N__4671));
    Span4Mux_h I__893 (
            .O(N__4674),
            .I(N__4668));
    InMux I__892 (
            .O(N__4671),
            .I(N__4665));
    Odrv4 I__891 (
            .O(N__4668),
            .I(CONSTANT_ONE_NET));
    LocalMux I__890 (
            .O(N__4665),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__889 (
            .O(N__4660),
            .I(N__4649));
    CascadeMux I__888 (
            .O(N__4659),
            .I(N__4641));
    InMux I__887 (
            .O(N__4658),
            .I(N__4638));
    InMux I__886 (
            .O(N__4657),
            .I(N__4635));
    CascadeMux I__885 (
            .O(N__4656),
            .I(N__4632));
    InMux I__884 (
            .O(N__4655),
            .I(N__4627));
    InMux I__883 (
            .O(N__4654),
            .I(N__4624));
    InMux I__882 (
            .O(N__4653),
            .I(N__4619));
    InMux I__881 (
            .O(N__4652),
            .I(N__4619));
    InMux I__880 (
            .O(N__4649),
            .I(N__4612));
    InMux I__879 (
            .O(N__4648),
            .I(N__4612));
    InMux I__878 (
            .O(N__4647),
            .I(N__4612));
    InMux I__877 (
            .O(N__4646),
            .I(N__4609));
    CascadeMux I__876 (
            .O(N__4645),
            .I(N__4604));
    InMux I__875 (
            .O(N__4644),
            .I(N__4593));
    InMux I__874 (
            .O(N__4641),
            .I(N__4593));
    LocalMux I__873 (
            .O(N__4638),
            .I(N__4588));
    LocalMux I__872 (
            .O(N__4635),
            .I(N__4588));
    InMux I__871 (
            .O(N__4632),
            .I(N__4581));
    InMux I__870 (
            .O(N__4631),
            .I(N__4581));
    InMux I__869 (
            .O(N__4630),
            .I(N__4581));
    LocalMux I__868 (
            .O(N__4627),
            .I(N__4576));
    LocalMux I__867 (
            .O(N__4624),
            .I(N__4576));
    LocalMux I__866 (
            .O(N__4619),
            .I(N__4571));
    LocalMux I__865 (
            .O(N__4612),
            .I(N__4571));
    LocalMux I__864 (
            .O(N__4609),
            .I(N__4568));
    InMux I__863 (
            .O(N__4608),
            .I(N__4563));
    InMux I__862 (
            .O(N__4607),
            .I(N__4563));
    InMux I__861 (
            .O(N__4604),
            .I(N__4560));
    InMux I__860 (
            .O(N__4603),
            .I(N__4553));
    InMux I__859 (
            .O(N__4602),
            .I(N__4553));
    InMux I__858 (
            .O(N__4601),
            .I(N__4553));
    InMux I__857 (
            .O(N__4600),
            .I(N__4550));
    InMux I__856 (
            .O(N__4599),
            .I(N__4547));
    InMux I__855 (
            .O(N__4598),
            .I(N__4544));
    LocalMux I__854 (
            .O(N__4593),
            .I(N__4539));
    Span4Mux_v I__853 (
            .O(N__4588),
            .I(N__4539));
    LocalMux I__852 (
            .O(N__4581),
            .I(N__4534));
    Span4Mux_h I__851 (
            .O(N__4576),
            .I(N__4534));
    Span4Mux_h I__850 (
            .O(N__4571),
            .I(N__4531));
    Span4Mux_h I__849 (
            .O(N__4568),
            .I(N__4522));
    LocalMux I__848 (
            .O(N__4563),
            .I(N__4522));
    LocalMux I__847 (
            .O(N__4560),
            .I(N__4522));
    LocalMux I__846 (
            .O(N__4553),
            .I(N__4522));
    LocalMux I__845 (
            .O(N__4550),
            .I(U400_SDRAM_SDRAM_COUNTER_0));
    LocalMux I__844 (
            .O(N__4547),
            .I(U400_SDRAM_SDRAM_COUNTER_0));
    LocalMux I__843 (
            .O(N__4544),
            .I(U400_SDRAM_SDRAM_COUNTER_0));
    Odrv4 I__842 (
            .O(N__4539),
            .I(U400_SDRAM_SDRAM_COUNTER_0));
    Odrv4 I__841 (
            .O(N__4534),
            .I(U400_SDRAM_SDRAM_COUNTER_0));
    Odrv4 I__840 (
            .O(N__4531),
            .I(U400_SDRAM_SDRAM_COUNTER_0));
    Odrv4 I__839 (
            .O(N__4522),
            .I(U400_SDRAM_SDRAM_COUNTER_0));
    CEMux I__838 (
            .O(N__4507),
            .I(N__4504));
    LocalMux I__837 (
            .O(N__4504),
            .I(N__4499));
    CEMux I__836 (
            .O(N__4503),
            .I(N__4496));
    CEMux I__835 (
            .O(N__4502),
            .I(N__4493));
    Span4Mux_h I__834 (
            .O(N__4499),
            .I(N__4490));
    LocalMux I__833 (
            .O(N__4496),
            .I(N__4487));
    LocalMux I__832 (
            .O(N__4493),
            .I(N__4484));
    Odrv4 I__831 (
            .O(N__4490),
            .I(U400_SDRAM_SDRAM_COUNTERe_0_i));
    Odrv4 I__830 (
            .O(N__4487),
            .I(U400_SDRAM_SDRAM_COUNTERe_0_i));
    Odrv4 I__829 (
            .O(N__4484),
            .I(U400_SDRAM_SDRAM_COUNTERe_0_i));
    InMux I__828 (
            .O(N__4477),
            .I(N__4472));
    InMux I__827 (
            .O(N__4476),
            .I(N__4467));
    InMux I__826 (
            .O(N__4475),
            .I(N__4467));
    LocalMux I__825 (
            .O(N__4472),
            .I(N__4464));
    LocalMux I__824 (
            .O(N__4467),
            .I(N__4461));
    Span4Mux_v I__823 (
            .O(N__4464),
            .I(N__4458));
    Odrv12 I__822 (
            .O(N__4461),
            .I(\U400_ADDRESS_DECODE.N_135_0 ));
    Odrv4 I__821 (
            .O(N__4458),
            .I(\U400_ADDRESS_DECODE.N_135_0 ));
    CascadeMux I__820 (
            .O(N__4453),
            .I(N__4449));
    InMux I__819 (
            .O(N__4452),
            .I(N__4441));
    InMux I__818 (
            .O(N__4449),
            .I(N__4441));
    InMux I__817 (
            .O(N__4448),
            .I(N__4441));
    LocalMux I__816 (
            .O(N__4441),
            .I(U400_SDRAM_TA_COUNTER_4));
    InMux I__815 (
            .O(N__4438),
            .I(N__4433));
    InMux I__814 (
            .O(N__4437),
            .I(N__4428));
    InMux I__813 (
            .O(N__4436),
            .I(N__4428));
    LocalMux I__812 (
            .O(N__4433),
            .I(U400_SDRAM_TA_COUNTER_1));
    LocalMux I__811 (
            .O(N__4428),
            .I(U400_SDRAM_TA_COUNTER_1));
    CascadeMux I__810 (
            .O(N__4423),
            .I(\U400_ADDRESS_DECODE.N_177_mux_cascade_ ));
    CascadeMux I__809 (
            .O(N__4420),
            .I(N__4416));
    CascadeMux I__808 (
            .O(N__4419),
            .I(N__4413));
    InMux I__807 (
            .O(N__4416),
            .I(N__4405));
    InMux I__806 (
            .O(N__4413),
            .I(N__4405));
    InMux I__805 (
            .O(N__4412),
            .I(N__4405));
    LocalMux I__804 (
            .O(N__4405),
            .I(U400_SDRAM_TA_COUNTER_0));
    InMux I__803 (
            .O(N__4402),
            .I(N__4389));
    InMux I__802 (
            .O(N__4401),
            .I(N__4389));
    InMux I__801 (
            .O(N__4400),
            .I(N__4389));
    InMux I__800 (
            .O(N__4399),
            .I(N__4389));
    InMux I__799 (
            .O(N__4398),
            .I(N__4386));
    LocalMux I__798 (
            .O(N__4389),
            .I(N__4383));
    LocalMux I__797 (
            .O(N__4386),
            .I(U400_SDRAM_TACK));
    Odrv4 I__796 (
            .O(N__4383),
            .I(U400_SDRAM_TACK));
    InMux I__795 (
            .O(N__4378),
            .I(N__4375));
    LocalMux I__794 (
            .O(N__4375),
            .I(N__4372));
    Span12Mux_v I__793 (
            .O(N__4372),
            .I(N__4369));
    Odrv12 I__792 (
            .O(N__4369),
            .I(RnW_c));
    CascadeMux I__791 (
            .O(N__4366),
            .I(N__4359));
    CascadeMux I__790 (
            .O(N__4365),
            .I(N__4356));
    CascadeMux I__789 (
            .O(N__4364),
            .I(N__4352));
    CascadeMux I__788 (
            .O(N__4363),
            .I(N__4349));
    InMux I__787 (
            .O(N__4362),
            .I(N__4344));
    InMux I__786 (
            .O(N__4359),
            .I(N__4341));
    InMux I__785 (
            .O(N__4356),
            .I(N__4338));
    InMux I__784 (
            .O(N__4355),
            .I(N__4335));
    InMux I__783 (
            .O(N__4352),
            .I(N__4330));
    InMux I__782 (
            .O(N__4349),
            .I(N__4330));
    InMux I__781 (
            .O(N__4348),
            .I(N__4326));
    CascadeMux I__780 (
            .O(N__4347),
            .I(N__4322));
    LocalMux I__779 (
            .O(N__4344),
            .I(N__4317));
    LocalMux I__778 (
            .O(N__4341),
            .I(N__4317));
    LocalMux I__777 (
            .O(N__4338),
            .I(N__4310));
    LocalMux I__776 (
            .O(N__4335),
            .I(N__4310));
    LocalMux I__775 (
            .O(N__4330),
            .I(N__4310));
    InMux I__774 (
            .O(N__4329),
            .I(N__4307));
    LocalMux I__773 (
            .O(N__4326),
            .I(N__4304));
    InMux I__772 (
            .O(N__4325),
            .I(N__4299));
    InMux I__771 (
            .O(N__4322),
            .I(N__4299));
    Span4Mux_h I__770 (
            .O(N__4317),
            .I(N__4296));
    Span4Mux_v I__769 (
            .O(N__4310),
            .I(N__4293));
    LocalMux I__768 (
            .O(N__4307),
            .I(U400_SDRAM_WRITE_CYCLE));
    Odrv4 I__767 (
            .O(N__4304),
            .I(U400_SDRAM_WRITE_CYCLE));
    LocalMux I__766 (
            .O(N__4299),
            .I(U400_SDRAM_WRITE_CYCLE));
    Odrv4 I__765 (
            .O(N__4296),
            .I(U400_SDRAM_WRITE_CYCLE));
    Odrv4 I__764 (
            .O(N__4293),
            .I(U400_SDRAM_WRITE_CYCLE));
    InMux I__763 (
            .O(N__4282),
            .I(N__4279));
    LocalMux I__762 (
            .O(N__4279),
            .I(N_48));
    InMux I__761 (
            .O(N__4276),
            .I(N__4273));
    LocalMux I__760 (
            .O(N__4273),
            .I(N_142_0));
    InMux I__759 (
            .O(N__4270),
            .I(N__4267));
    LocalMux I__758 (
            .O(N__4267),
            .I(N__4263));
    InMux I__757 (
            .O(N__4266),
            .I(N__4260));
    Odrv12 I__756 (
            .O(N__4263),
            .I(\U400_ADDRESS_DECODE.N_12_0 ));
    LocalMux I__755 (
            .O(N__4260),
            .I(\U400_ADDRESS_DECODE.N_12_0 ));
    InMux I__754 (
            .O(N__4255),
            .I(N__4252));
    LocalMux I__753 (
            .O(N__4252),
            .I(N__4249));
    Odrv4 I__752 (
            .O(N__4249),
            .I(\U400_ADDRESS_DECODE.N_21_0 ));
    CascadeMux I__751 (
            .O(N__4246),
            .I(N__4242));
    CascadeMux I__750 (
            .O(N__4245),
            .I(N__4239));
    InMux I__749 (
            .O(N__4242),
            .I(N__4234));
    InMux I__748 (
            .O(N__4239),
            .I(N__4234));
    LocalMux I__747 (
            .O(N__4234),
            .I(N__4231));
    Odrv12 I__746 (
            .O(N__4231),
            .I(A_c_23));
    InMux I__745 (
            .O(N__4228),
            .I(N__4225));
    LocalMux I__744 (
            .O(N__4225),
            .I(N_137_0));
    InMux I__743 (
            .O(N__4222),
            .I(N__4219));
    LocalMux I__742 (
            .O(N__4219),
            .I(N__4215));
    InMux I__741 (
            .O(N__4218),
            .I(N__4212));
    Odrv4 I__740 (
            .O(N__4215),
            .I(N_190_mux));
    LocalMux I__739 (
            .O(N__4212),
            .I(N_190_mux));
    InMux I__738 (
            .O(N__4207),
            .I(N__4204));
    LocalMux I__737 (
            .O(N__4204),
            .I(N_138_0));
    InMux I__736 (
            .O(N__4201),
            .I(N__4197));
    InMux I__735 (
            .O(N__4200),
            .I(N__4194));
    LocalMux I__734 (
            .O(N__4197),
            .I(N_23_0));
    LocalMux I__733 (
            .O(N__4194),
            .I(N_23_0));
    CascadeMux I__732 (
            .O(N__4189),
            .I(N__4185));
    CascadeMux I__731 (
            .O(N__4188),
            .I(N__4182));
    InMux I__730 (
            .O(N__4185),
            .I(N__4177));
    InMux I__729 (
            .O(N__4182),
            .I(N__4177));
    LocalMux I__728 (
            .O(N__4177),
            .I(\U400_SDRAM.CS1_ENZ0 ));
    IoInMux I__727 (
            .O(N__4174),
            .I(N__4171));
    LocalMux I__726 (
            .O(N__4171),
            .I(N__4168));
    Odrv12 I__725 (
            .O(N__4168),
            .I(CS1n_c));
    InMux I__724 (
            .O(N__4165),
            .I(N__4162));
    LocalMux I__723 (
            .O(N__4162),
            .I(\U400_ADDRESS_DECODE.m94_amZ0Z_1 ));
    CascadeMux I__722 (
            .O(N__4159),
            .I(\U400_ADDRESS_DECODE.m94_amZ0_cascade_ ));
    InMux I__721 (
            .O(N__4156),
            .I(N__4153));
    LocalMux I__720 (
            .O(N__4153),
            .I(\U400_ADDRESS_DECODE.N_95_0 ));
    InMux I__719 (
            .O(N__4150),
            .I(N__4141));
    InMux I__718 (
            .O(N__4149),
            .I(N__4136));
    InMux I__717 (
            .O(N__4148),
            .I(N__4136));
    InMux I__716 (
            .O(N__4147),
            .I(N__4131));
    InMux I__715 (
            .O(N__4146),
            .I(N__4131));
    InMux I__714 (
            .O(N__4145),
            .I(N__4126));
    InMux I__713 (
            .O(N__4144),
            .I(N__4126));
    LocalMux I__712 (
            .O(N__4141),
            .I(U400_SDRAM_RAM_CYCLE_START));
    LocalMux I__711 (
            .O(N__4136),
            .I(U400_SDRAM_RAM_CYCLE_START));
    LocalMux I__710 (
            .O(N__4131),
            .I(U400_SDRAM_RAM_CYCLE_START));
    LocalMux I__709 (
            .O(N__4126),
            .I(U400_SDRAM_RAM_CYCLE_START));
    InMux I__708 (
            .O(N__4117),
            .I(N__4112));
    InMux I__707 (
            .O(N__4116),
            .I(N__4107));
    InMux I__706 (
            .O(N__4115),
            .I(N__4107));
    LocalMux I__705 (
            .O(N__4112),
            .I(\U400_ADDRESS_DECODE.N_15_0 ));
    LocalMux I__704 (
            .O(N__4107),
            .I(\U400_ADDRESS_DECODE.N_15_0 ));
    CascadeMux I__703 (
            .O(N__4102),
            .I(N__4097));
    CascadeMux I__702 (
            .O(N__4101),
            .I(N__4094));
    InMux I__701 (
            .O(N__4100),
            .I(N__4091));
    InMux I__700 (
            .O(N__4097),
            .I(N__4088));
    InMux I__699 (
            .O(N__4094),
            .I(N__4085));
    LocalMux I__698 (
            .O(N__4091),
            .I(N_13_0));
    LocalMux I__697 (
            .O(N__4088),
            .I(N_13_0));
    LocalMux I__696 (
            .O(N__4085),
            .I(N_13_0));
    CascadeMux I__695 (
            .O(N__4078),
            .I(N__4072));
    InMux I__694 (
            .O(N__4077),
            .I(N__4068));
    InMux I__693 (
            .O(N__4076),
            .I(N__4065));
    InMux I__692 (
            .O(N__4075),
            .I(N__4062));
    InMux I__691 (
            .O(N__4072),
            .I(N__4056));
    InMux I__690 (
            .O(N__4071),
            .I(N__4056));
    LocalMux I__689 (
            .O(N__4068),
            .I(N__4050));
    LocalMux I__688 (
            .O(N__4065),
            .I(N__4050));
    LocalMux I__687 (
            .O(N__4062),
            .I(N__4047));
    InMux I__686 (
            .O(N__4061),
            .I(N__4044));
    LocalMux I__685 (
            .O(N__4056),
            .I(N__4041));
    InMux I__684 (
            .O(N__4055),
            .I(N__4038));
    Span4Mux_h I__683 (
            .O(N__4050),
            .I(N__4035));
    Span4Mux_v I__682 (
            .O(N__4047),
            .I(N__4026));
    LocalMux I__681 (
            .O(N__4044),
            .I(N__4026));
    Span4Mux_h I__680 (
            .O(N__4041),
            .I(N__4026));
    LocalMux I__679 (
            .O(N__4038),
            .I(N__4026));
    Odrv4 I__678 (
            .O(N__4035),
            .I(U400_SDRAM_SDRAM_CMD11));
    Odrv4 I__677 (
            .O(N__4026),
            .I(U400_SDRAM_SDRAM_CMD11));
    CascadeMux I__676 (
            .O(N__4021),
            .I(\U400_ADDRESS_DECODE.m20_amZ0_cascade_ ));
    CascadeMux I__675 (
            .O(N__4018),
            .I(N__4011));
    InMux I__674 (
            .O(N__4017),
            .I(N__3992));
    InMux I__673 (
            .O(N__4016),
            .I(N__3992));
    InMux I__672 (
            .O(N__4015),
            .I(N__3992));
    InMux I__671 (
            .O(N__4014),
            .I(N__3983));
    InMux I__670 (
            .O(N__4011),
            .I(N__3983));
    InMux I__669 (
            .O(N__4010),
            .I(N__3983));
    InMux I__668 (
            .O(N__4009),
            .I(N__3978));
    InMux I__667 (
            .O(N__4008),
            .I(N__3978));
    InMux I__666 (
            .O(N__4007),
            .I(N__3972));
    InMux I__665 (
            .O(N__4006),
            .I(N__3972));
    InMux I__664 (
            .O(N__4005),
            .I(N__3963));
    InMux I__663 (
            .O(N__4004),
            .I(N__3963));
    InMux I__662 (
            .O(N__4003),
            .I(N__3963));
    InMux I__661 (
            .O(N__4002),
            .I(N__3956));
    InMux I__660 (
            .O(N__4001),
            .I(N__3956));
    InMux I__659 (
            .O(N__4000),
            .I(N__3956));
    InMux I__658 (
            .O(N__3999),
            .I(N__3953));
    LocalMux I__657 (
            .O(N__3992),
            .I(N__3950));
    InMux I__656 (
            .O(N__3991),
            .I(N__3947));
    InMux I__655 (
            .O(N__3990),
            .I(N__3944));
    LocalMux I__654 (
            .O(N__3983),
            .I(N__3941));
    LocalMux I__653 (
            .O(N__3978),
            .I(N__3938));
    InMux I__652 (
            .O(N__3977),
            .I(N__3935));
    LocalMux I__651 (
            .O(N__3972),
            .I(N__3931));
    InMux I__650 (
            .O(N__3971),
            .I(N__3926));
    InMux I__649 (
            .O(N__3970),
            .I(N__3926));
    LocalMux I__648 (
            .O(N__3963),
            .I(N__3921));
    LocalMux I__647 (
            .O(N__3956),
            .I(N__3921));
    LocalMux I__646 (
            .O(N__3953),
            .I(N__3916));
    Span4Mux_v I__645 (
            .O(N__3950),
            .I(N__3916));
    LocalMux I__644 (
            .O(N__3947),
            .I(N__3913));
    LocalMux I__643 (
            .O(N__3944),
            .I(N__3904));
    Span4Mux_h I__642 (
            .O(N__3941),
            .I(N__3904));
    Span4Mux_h I__641 (
            .O(N__3938),
            .I(N__3904));
    LocalMux I__640 (
            .O(N__3935),
            .I(N__3904));
    InMux I__639 (
            .O(N__3934),
            .I(N__3901));
    Span4Mux_h I__638 (
            .O(N__3931),
            .I(N__3898));
    LocalMux I__637 (
            .O(N__3926),
            .I(N__3893));
    Span4Mux_h I__636 (
            .O(N__3921),
            .I(N__3893));
    Odrv4 I__635 (
            .O(N__3916),
            .I(U400_SDRAM_SDRAM_COUNTER_3));
    Odrv12 I__634 (
            .O(N__3913),
            .I(U400_SDRAM_SDRAM_COUNTER_3));
    Odrv4 I__633 (
            .O(N__3904),
            .I(U400_SDRAM_SDRAM_COUNTER_3));
    LocalMux I__632 (
            .O(N__3901),
            .I(U400_SDRAM_SDRAM_COUNTER_3));
    Odrv4 I__631 (
            .O(N__3898),
            .I(U400_SDRAM_SDRAM_COUNTER_3));
    Odrv4 I__630 (
            .O(N__3893),
            .I(U400_SDRAM_SDRAM_COUNTER_3));
    CascadeMux I__629 (
            .O(N__3880),
            .I(N__3876));
    InMux I__628 (
            .O(N__3879),
            .I(N__3872));
    InMux I__627 (
            .O(N__3876),
            .I(N__3867));
    InMux I__626 (
            .O(N__3875),
            .I(N__3867));
    LocalMux I__625 (
            .O(N__3872),
            .I(\U400_ADDRESS_DECODE.N_6_0 ));
    LocalMux I__624 (
            .O(N__3867),
            .I(\U400_ADDRESS_DECODE.N_6_0 ));
    InMux I__623 (
            .O(N__3862),
            .I(N__3859));
    LocalMux I__622 (
            .O(N__3859),
            .I(\U400_ADDRESS_DECODE.m94_bmZ0 ));
    CascadeMux I__621 (
            .O(N__3856),
            .I(N__3852));
    InMux I__620 (
            .O(N__3855),
            .I(N__3843));
    InMux I__619 (
            .O(N__3852),
            .I(N__3840));
    InMux I__618 (
            .O(N__3851),
            .I(N__3837));
    CascadeMux I__617 (
            .O(N__3850),
            .I(N__3834));
    InMux I__616 (
            .O(N__3849),
            .I(N__3831));
    CascadeMux I__615 (
            .O(N__3848),
            .I(N__3827));
    InMux I__614 (
            .O(N__3847),
            .I(N__3819));
    InMux I__613 (
            .O(N__3846),
            .I(N__3816));
    LocalMux I__612 (
            .O(N__3843),
            .I(N__3810));
    LocalMux I__611 (
            .O(N__3840),
            .I(N__3805));
    LocalMux I__610 (
            .O(N__3837),
            .I(N__3805));
    InMux I__609 (
            .O(N__3834),
            .I(N__3802));
    LocalMux I__608 (
            .O(N__3831),
            .I(N__3799));
    InMux I__607 (
            .O(N__3830),
            .I(N__3792));
    InMux I__606 (
            .O(N__3827),
            .I(N__3792));
    InMux I__605 (
            .O(N__3826),
            .I(N__3792));
    InMux I__604 (
            .O(N__3825),
            .I(N__3789));
    InMux I__603 (
            .O(N__3824),
            .I(N__3784));
    InMux I__602 (
            .O(N__3823),
            .I(N__3784));
    InMux I__601 (
            .O(N__3822),
            .I(N__3781));
    LocalMux I__600 (
            .O(N__3819),
            .I(N__3776));
    LocalMux I__599 (
            .O(N__3816),
            .I(N__3776));
    InMux I__598 (
            .O(N__3815),
            .I(N__3769));
    InMux I__597 (
            .O(N__3814),
            .I(N__3769));
    InMux I__596 (
            .O(N__3813),
            .I(N__3769));
    Span4Mux_v I__595 (
            .O(N__3810),
            .I(N__3764));
    Span4Mux_v I__594 (
            .O(N__3805),
            .I(N__3764));
    LocalMux I__593 (
            .O(N__3802),
            .I(N__3753));
    Span4Mux_h I__592 (
            .O(N__3799),
            .I(N__3753));
    LocalMux I__591 (
            .O(N__3792),
            .I(N__3753));
    LocalMux I__590 (
            .O(N__3789),
            .I(N__3753));
    LocalMux I__589 (
            .O(N__3784),
            .I(N__3753));
    LocalMux I__588 (
            .O(N__3781),
            .I(U400_SDRAM_SDRAM_COUNTER_1));
    Odrv12 I__587 (
            .O(N__3776),
            .I(U400_SDRAM_SDRAM_COUNTER_1));
    LocalMux I__586 (
            .O(N__3769),
            .I(U400_SDRAM_SDRAM_COUNTER_1));
    Odrv4 I__585 (
            .O(N__3764),
            .I(U400_SDRAM_SDRAM_COUNTER_1));
    Odrv4 I__584 (
            .O(N__3753),
            .I(U400_SDRAM_SDRAM_COUNTER_1));
    InMux I__583 (
            .O(N__3742),
            .I(N__3739));
    LocalMux I__582 (
            .O(N__3739),
            .I(\U400_ADDRESS_DECODE.m20_bmZ0 ));
    InMux I__581 (
            .O(N__3736),
            .I(N__3733));
    LocalMux I__580 (
            .O(N__3733),
            .I(N__3730));
    Span4Mux_v I__579 (
            .O(N__3730),
            .I(N__3727));
    Span4Mux_h I__578 (
            .O(N__3727),
            .I(N__3723));
    InMux I__577 (
            .O(N__3726),
            .I(N__3720));
    Odrv4 I__576 (
            .O(N__3723),
            .I(\U400_ADDRESS_DECODE.N_20_0 ));
    LocalMux I__575 (
            .O(N__3720),
            .I(\U400_ADDRESS_DECODE.N_20_0 ));
    InMux I__574 (
            .O(N__3715),
            .I(N__3711));
    InMux I__573 (
            .O(N__3714),
            .I(N__3708));
    LocalMux I__572 (
            .O(N__3711),
            .I(\U400_ADDRESS_DECODE.N_179_mux ));
    LocalMux I__571 (
            .O(N__3708),
            .I(\U400_ADDRESS_DECODE.N_179_mux ));
    CascadeMux I__570 (
            .O(N__3703),
            .I(\U400_ADDRESS_DECODE.N_8_0_cascade_ ));
    SRMux I__569 (
            .O(N__3700),
            .I(N__3696));
    SRMux I__568 (
            .O(N__3699),
            .I(N__3692));
    LocalMux I__567 (
            .O(N__3696),
            .I(N__3689));
    SRMux I__566 (
            .O(N__3695),
            .I(N__3686));
    LocalMux I__565 (
            .O(N__3692),
            .I(N__3683));
    Span4Mux_s3_v I__564 (
            .O(N__3689),
            .I(N__3678));
    LocalMux I__563 (
            .O(N__3686),
            .I(N__3678));
    Span4Mux_s2_h I__562 (
            .O(N__3683),
            .I(N__3673));
    Span4Mux_s2_h I__561 (
            .O(N__3678),
            .I(N__3673));
    Odrv4 I__560 (
            .O(N__3673),
            .I(\U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2 ));
    CascadeMux I__559 (
            .O(N__3670),
            .I(N__3667));
    InMux I__558 (
            .O(N__3667),
            .I(N__3661));
    InMux I__557 (
            .O(N__3666),
            .I(N__3661));
    LocalMux I__556 (
            .O(N__3661),
            .I(N__3658));
    Span4Mux_v I__555 (
            .O(N__3658),
            .I(N__3655));
    Span4Mux_h I__554 (
            .O(N__3655),
            .I(N__3652));
    Odrv4 I__553 (
            .O(N__3652),
            .I(TSn_c));
    InMux I__552 (
            .O(N__3649),
            .I(N__3646));
    LocalMux I__551 (
            .O(N__3646),
            .I(\U400_ADDRESS_DECODE.m165_nsZ0Z_1 ));
    CascadeMux I__550 (
            .O(N__3643),
            .I(N_13_0_cascade_));
    InMux I__549 (
            .O(N__3640),
            .I(N__3632));
    InMux I__548 (
            .O(N__3639),
            .I(N__3627));
    InMux I__547 (
            .O(N__3638),
            .I(N__3627));
    InMux I__546 (
            .O(N__3637),
            .I(N__3623));
    InMux I__545 (
            .O(N__3636),
            .I(N__3620));
    InMux I__544 (
            .O(N__3635),
            .I(N__3617));
    LocalMux I__543 (
            .O(N__3632),
            .I(N__3612));
    LocalMux I__542 (
            .O(N__3627),
            .I(N__3612));
    InMux I__541 (
            .O(N__3626),
            .I(N__3609));
    LocalMux I__540 (
            .O(N__3623),
            .I(\U400_ADDRESS_DECODE.N_10_0 ));
    LocalMux I__539 (
            .O(N__3620),
            .I(\U400_ADDRESS_DECODE.N_10_0 ));
    LocalMux I__538 (
            .O(N__3617),
            .I(\U400_ADDRESS_DECODE.N_10_0 ));
    Odrv4 I__537 (
            .O(N__3612),
            .I(\U400_ADDRESS_DECODE.N_10_0 ));
    LocalMux I__536 (
            .O(N__3609),
            .I(\U400_ADDRESS_DECODE.N_10_0 ));
    InMux I__535 (
            .O(N__3598),
            .I(N__3593));
    InMux I__534 (
            .O(N__3597),
            .I(N__3590));
    InMux I__533 (
            .O(N__3596),
            .I(N__3587));
    LocalMux I__532 (
            .O(N__3593),
            .I(N__3584));
    LocalMux I__531 (
            .O(N__3590),
            .I(N__3581));
    LocalMux I__530 (
            .O(N__3587),
            .I(N__3577));
    Span4Mux_v I__529 (
            .O(N__3584),
            .I(N__3572));
    Span4Mux_h I__528 (
            .O(N__3581),
            .I(N__3572));
    InMux I__527 (
            .O(N__3580),
            .I(N__3569));
    Odrv4 I__526 (
            .O(N__3577),
            .I(\U400_ADDRESS_DECODE.N_8_0 ));
    Odrv4 I__525 (
            .O(N__3572),
            .I(\U400_ADDRESS_DECODE.N_8_0 ));
    LocalMux I__524 (
            .O(N__3569),
            .I(\U400_ADDRESS_DECODE.N_8_0 ));
    CascadeMux I__523 (
            .O(N__3562),
            .I(\U400_ADDRESS_DECODE.N_179_mux_cascade_ ));
    InMux I__522 (
            .O(N__3559),
            .I(N__3554));
    InMux I__521 (
            .O(N__3558),
            .I(N__3551));
    InMux I__520 (
            .O(N__3557),
            .I(N__3548));
    LocalMux I__519 (
            .O(N__3554),
            .I(\U400_ADDRESS_DECODE.N_47_0 ));
    LocalMux I__518 (
            .O(N__3551),
            .I(\U400_ADDRESS_DECODE.N_47_0 ));
    LocalMux I__517 (
            .O(N__3548),
            .I(\U400_ADDRESS_DECODE.N_47_0 ));
    InMux I__516 (
            .O(N__3541),
            .I(N__3538));
    LocalMux I__515 (
            .O(N__3538),
            .I(\U400_ADDRESS_DECODE.N_62_0 ));
    CascadeMux I__514 (
            .O(N__3535),
            .I(\U400_ADDRESS_DECODE.N_62_0_cascade_ ));
    CascadeMux I__513 (
            .O(N__3532),
            .I(\U400_ADDRESS_DECODE.m141_bmZ0_cascade_ ));
    InMux I__512 (
            .O(N__3529),
            .I(N__3526));
    LocalMux I__511 (
            .O(N__3526),
            .I(\U400_ADDRESS_DECODE.m141_amZ0 ));
    CascadeMux I__510 (
            .O(N__3523),
            .I(N__3519));
    CascadeMux I__509 (
            .O(N__3522),
            .I(N__3516));
    InMux I__508 (
            .O(N__3519),
            .I(N__3513));
    InMux I__507 (
            .O(N__3516),
            .I(N__3510));
    LocalMux I__506 (
            .O(N__3513),
            .I(\U400_SDRAM.CS0_ENZ0 ));
    LocalMux I__505 (
            .O(N__3510),
            .I(\U400_SDRAM.CS0_ENZ0 ));
    IoInMux I__504 (
            .O(N__3505),
            .I(N__3502));
    LocalMux I__503 (
            .O(N__3502),
            .I(N__3499));
    IoSpan4Mux I__502 (
            .O(N__3499),
            .I(N__3496));
    Span4Mux_s2_h I__501 (
            .O(N__3496),
            .I(N__3493));
    Odrv4 I__500 (
            .O(N__3493),
            .I(CS0n_c));
    CascadeMux I__499 (
            .O(N__3490),
            .I(N__3487));
    InMux I__498 (
            .O(N__3487),
            .I(N__3484));
    LocalMux I__497 (
            .O(N__3484),
            .I(N__3481));
    Span4Mux_v I__496 (
            .O(N__3481),
            .I(N__3478));
    Sp12to4 I__495 (
            .O(N__3478),
            .I(N__3475));
    Span12Mux_s9_h I__494 (
            .O(N__3475),
            .I(N__3472));
    Odrv12 I__493 (
            .O(N__3472),
            .I(A_c_26));
    IoInMux I__492 (
            .O(N__3469),
            .I(N__3466));
    LocalMux I__491 (
            .O(N__3466),
            .I(N__3463));
    Odrv4 I__490 (
            .O(N__3463),
            .I(MA_c_12));
    CascadeMux I__489 (
            .O(N__3460),
            .I(N__3457));
    InMux I__488 (
            .O(N__3457),
            .I(N__3454));
    LocalMux I__487 (
            .O(N__3454),
            .I(N__3451));
    Sp12to4 I__486 (
            .O(N__3451),
            .I(N__3448));
    Span12Mux_s10_v I__485 (
            .O(N__3448),
            .I(N__3445));
    Odrv12 I__484 (
            .O(N__3445),
            .I(A_c_19));
    IoInMux I__483 (
            .O(N__3442),
            .I(N__3439));
    LocalMux I__482 (
            .O(N__3439),
            .I(N__3436));
    Odrv4 I__481 (
            .O(N__3436),
            .I(MA_c_9));
    CascadeMux I__480 (
            .O(N__3433),
            .I(N__3429));
    InMux I__479 (
            .O(N__3432),
            .I(N__3426));
    InMux I__478 (
            .O(N__3429),
            .I(N__3423));
    LocalMux I__477 (
            .O(N__3426),
            .I(N__3420));
    LocalMux I__476 (
            .O(N__3423),
            .I(U400_SDRAM_RAM_CYCLE));
    Odrv12 I__475 (
            .O(N__3420),
            .I(U400_SDRAM_RAM_CYCLE));
    InMux I__474 (
            .O(N__3415),
            .I(N__3412));
    LocalMux I__473 (
            .O(N__3412),
            .I(U400_SDRAM_RAM_CYCLE_START_2_0));
    InMux I__472 (
            .O(N__3409),
            .I(N__3406));
    LocalMux I__471 (
            .O(N__3406),
            .I(\U400_ADDRESS_DECODE.N_33_0 ));
    InMux I__470 (
            .O(N__3403),
            .I(N__3400));
    LocalMux I__469 (
            .O(N__3400),
            .I(\U400_ADDRESS_DECODE.m43_amZ0 ));
    InMux I__468 (
            .O(N__3397),
            .I(N__3394));
    LocalMux I__467 (
            .O(N__3394),
            .I(\U400_ADDRESS_DECODE.m87_nsZ0Z_1 ));
    CascadeMux I__466 (
            .O(N__3391),
            .I(\U400_ADDRESS_DECODE.N_88_0_cascade_ ));
    CascadeMux I__465 (
            .O(N__3388),
            .I(N_96_0_cascade_));
    InMux I__464 (
            .O(N__3385),
            .I(N__3381));
    InMux I__463 (
            .O(N__3384),
            .I(N__3378));
    LocalMux I__462 (
            .O(N__3381),
            .I(N_73_0));
    LocalMux I__461 (
            .O(N__3378),
            .I(N_73_0));
    InMux I__460 (
            .O(N__3373),
            .I(N__3370));
    LocalMux I__459 (
            .O(N__3370),
            .I(\U400_ADDRESS_DECODE.m63_nsZ0Z_1 ));
    CascadeMux I__458 (
            .O(N__3367),
            .I(\U400_ADDRESS_DECODE.N_139_0_cascade_ ));
    CascadeMux I__457 (
            .O(N__3364),
            .I(N__3360));
    CascadeMux I__456 (
            .O(N__3363),
            .I(N__3357));
    InMux I__455 (
            .O(N__3360),
            .I(N__3354));
    InMux I__454 (
            .O(N__3357),
            .I(N__3351));
    LocalMux I__453 (
            .O(N__3354),
            .I(N__3348));
    LocalMux I__452 (
            .O(N__3351),
            .I(\U400_ADDRESS_DECODE.m133Z0Z_0 ));
    Odrv12 I__451 (
            .O(N__3348),
            .I(\U400_ADDRESS_DECODE.m133Z0Z_0 ));
    CascadeMux I__450 (
            .O(N__3343),
            .I(\U400_ADDRESS_DECODE.m41_amZ0_cascade_ ));
    InMux I__449 (
            .O(N__3340),
            .I(N__3337));
    LocalMux I__448 (
            .O(N__3337),
            .I(\U400_ADDRESS_DECODE.m41_bmZ0 ));
    CascadeMux I__447 (
            .O(N__3334),
            .I(\U400_ADDRESS_DECODE.m54Z0Z_0_cascade_ ));
    InMux I__446 (
            .O(N__3331),
            .I(N__3328));
    LocalMux I__445 (
            .O(N__3328),
            .I(\U400_ADDRESS_DECODE.m56_bmZ0 ));
    InMux I__444 (
            .O(N__3325),
            .I(N__3320));
    InMux I__443 (
            .O(N__3324),
            .I(N__3317));
    InMux I__442 (
            .O(N__3323),
            .I(N__3314));
    LocalMux I__441 (
            .O(N__3320),
            .I(\U400_ADDRESS_DECODE.N_185 ));
    LocalMux I__440 (
            .O(N__3317),
            .I(\U400_ADDRESS_DECODE.N_185 ));
    LocalMux I__439 (
            .O(N__3314),
            .I(\U400_ADDRESS_DECODE.N_185 ));
    CascadeMux I__438 (
            .O(N__3307),
            .I(\U400_ADDRESS_DECODE.N_185_mux_cascade_ ));
    InMux I__437 (
            .O(N__3304),
            .I(N__3301));
    LocalMux I__436 (
            .O(N__3301),
            .I(N__3298));
    Odrv4 I__435 (
            .O(N__3298),
            .I(\U400_ADDRESS_DECODE.N_42_0 ));
    CascadeMux I__434 (
            .O(N__3295),
            .I(\U400_ADDRESS_DECODE.m43_bmZ0_cascade_ ));
    InMux I__433 (
            .O(N__3292),
            .I(N__3289));
    LocalMux I__432 (
            .O(N__3289),
            .I(N_44_0));
    InMux I__431 (
            .O(N__3286),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_5 ));
    InMux I__430 (
            .O(N__3283),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_6 ));
    InMux I__429 (
            .O(N__3280),
            .I(N__3276));
    InMux I__428 (
            .O(N__3279),
            .I(N__3273));
    LocalMux I__427 (
            .O(N__3276),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__426 (
            .O(N__3273),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__425 (
            .O(N__3268),
            .I(N__3264));
    InMux I__424 (
            .O(N__3267),
            .I(N__3261));
    LocalMux I__423 (
            .O(N__3264),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__422 (
            .O(N__3261),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__421 (
            .O(N__3256),
            .I(N__3252));
    InMux I__420 (
            .O(N__3255),
            .I(N__3249));
    InMux I__419 (
            .O(N__3252),
            .I(N__3246));
    LocalMux I__418 (
            .O(N__3249),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__417 (
            .O(N__3246),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__416 (
            .O(N__3241),
            .I(N__3237));
    InMux I__415 (
            .O(N__3240),
            .I(N__3234));
    LocalMux I__414 (
            .O(N__3237),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__413 (
            .O(N__3234),
            .I(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__412 (
            .O(N__3229),
            .I(N_60_cascade_));
    CascadeMux I__411 (
            .O(N__3226),
            .I(\U400_ADDRESS_DECODE.N_98_0_cascade_ ));
    InMux I__410 (
            .O(N__3223),
            .I(N__3216));
    InMux I__409 (
            .O(N__3222),
            .I(N__3216));
    InMux I__408 (
            .O(N__3221),
            .I(N__3213));
    LocalMux I__407 (
            .O(N__3216),
            .I(U400_SDRAM_SDRAM_CMD_5_sqmuxa));
    LocalMux I__406 (
            .O(N__3213),
            .I(U400_SDRAM_SDRAM_CMD_5_sqmuxa));
    CascadeMux I__405 (
            .O(N__3208),
            .I(N__3205));
    InMux I__404 (
            .O(N__3205),
            .I(N__3202));
    LocalMux I__403 (
            .O(N__3202),
            .I(N__3199));
    Span12Mux_s10_v I__402 (
            .O(N__3199),
            .I(N__3196));
    Odrv12 I__401 (
            .O(N__3196),
            .I(A_c_18));
    InMux I__400 (
            .O(N__3193),
            .I(N__3190));
    LocalMux I__399 (
            .O(N__3190),
            .I(N__3187));
    Span4Mux_h I__398 (
            .O(N__3187),
            .I(N__3184));
    Sp12to4 I__397 (
            .O(N__3184),
            .I(N__3181));
    Span12Mux_v I__396 (
            .O(N__3181),
            .I(N__3178));
    Odrv12 I__395 (
            .O(N__3178),
            .I(A_c_24));
    IoInMux I__394 (
            .O(N__3175),
            .I(N__3172));
    LocalMux I__393 (
            .O(N__3172),
            .I(N__3169));
    Span4Mux_s1_v I__392 (
            .O(N__3169),
            .I(N__3166));
    Odrv4 I__391 (
            .O(N__3166),
            .I(MA_c_8));
    InMux I__390 (
            .O(N__3163),
            .I(N__3160));
    LocalMux I__389 (
            .O(N__3160),
            .I(N__3157));
    Odrv12 I__388 (
            .O(N__3157),
            .I(A_c_8));
    CascadeMux I__387 (
            .O(N__3154),
            .I(N__3151));
    InMux I__386 (
            .O(N__3151),
            .I(N__3148));
    LocalMux I__385 (
            .O(N__3148),
            .I(N__3145));
    Span4Mux_v I__384 (
            .O(N__3145),
            .I(N__3142));
    Span4Mux_v I__383 (
            .O(N__3142),
            .I(N__3139));
    Odrv4 I__382 (
            .O(N__3139),
            .I(A_c_16));
    IoInMux I__381 (
            .O(N__3136),
            .I(N__3133));
    LocalMux I__380 (
            .O(N__3133),
            .I(N__3130));
    Odrv12 I__379 (
            .O(N__3130),
            .I(MA_c_6));
    InMux I__378 (
            .O(N__3127),
            .I(N__3124));
    LocalMux I__377 (
            .O(N__3124),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_1 ));
    InMux I__376 (
            .O(N__3121),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_0 ));
    InMux I__375 (
            .O(N__3118),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_1 ));
    InMux I__374 (
            .O(N__3115),
            .I(N__3112));
    LocalMux I__373 (
            .O(N__3112),
            .I(\U400_SDRAM.SDRAM_COUNTER_s_3 ));
    InMux I__372 (
            .O(N__3109),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_2 ));
    InMux I__371 (
            .O(N__3106),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_3 ));
    InMux I__370 (
            .O(N__3103),
            .I(\U400_SDRAM.SDRAM_COUNTER_cry_4 ));
    CascadeMux I__369 (
            .O(N__3100),
            .I(\U400_ADDRESS_DECODE.m71_amZ0_cascade_ ));
    InMux I__368 (
            .O(N__3097),
            .I(N__3094));
    LocalMux I__367 (
            .O(N__3094),
            .I(\U400_ADDRESS_DECODE.m71_bmZ0 ));
    CascadeMux I__366 (
            .O(N__3091),
            .I(\U400_ADDRESS_DECODE.N_72_0_cascade_ ));
    CascadeMux I__365 (
            .O(N__3088),
            .I(N_73_0_cascade_));
    InMux I__364 (
            .O(N__3085),
            .I(N__3082));
    LocalMux I__363 (
            .O(N__3082),
            .I(\U400_ADDRESS_DECODE.m56_amZ0 ));
    InMux I__362 (
            .O(N__3079),
            .I(N__3076));
    LocalMux I__361 (
            .O(N__3076),
            .I(N_57_0));
    CascadeMux I__360 (
            .O(N__3073),
            .I(\U400_ADDRESS_DECODE.N_7_0_cascade_ ));
    IoInMux I__359 (
            .O(N__3070),
            .I(N__3067));
    LocalMux I__358 (
            .O(N__3067),
            .I(N__3064));
    Odrv12 I__357 (
            .O(N__3064),
            .I(RESETn_c_i));
    InMux I__356 (
            .O(N__3061),
            .I(N__3058));
    LocalMux I__355 (
            .O(N__3058),
            .I(N__3055));
    Odrv12 I__354 (
            .O(N__3055),
            .I(A_c_9));
    CascadeMux I__353 (
            .O(N__3052),
            .I(N__3049));
    InMux I__352 (
            .O(N__3049),
            .I(N__3046));
    LocalMux I__351 (
            .O(N__3046),
            .I(N__3043));
    Span4Mux_v I__350 (
            .O(N__3043),
            .I(N__3040));
    Odrv4 I__349 (
            .O(N__3040),
            .I(A_c_17));
    IoInMux I__348 (
            .O(N__3037),
            .I(N__3034));
    LocalMux I__347 (
            .O(N__3034),
            .I(N__3031));
    Span4Mux_s1_v I__346 (
            .O(N__3031),
            .I(N__3028));
    Odrv4 I__345 (
            .O(N__3028),
            .I(MA_c_7));
    CascadeMux I__344 (
            .O(N__3025),
            .I(\U400_ADDRESS_DECODE.m84_amZ0_cascade_ ));
    InMux I__343 (
            .O(N__3022),
            .I(N__3019));
    LocalMux I__342 (
            .O(N__3019),
            .I(\U400_ADDRESS_DECODE.m84_bmZ0 ));
    InMux I__341 (
            .O(N__3016),
            .I(N__3013));
    LocalMux I__340 (
            .O(N__3013),
            .I(N_85_0));
    InMux I__339 (
            .O(N__3010),
            .I(N__3007));
    LocalMux I__338 (
            .O(N__3007),
            .I(\U400_ADDRESS_DECODE.N_46_0 ));
    CascadeMux I__337 (
            .O(N__3004),
            .I(\U400_ADDRESS_DECODE.N_47_0_cascade_ ));
    InMux I__336 (
            .O(N__3001),
            .I(N__2998));
    LocalMux I__335 (
            .O(N__2998),
            .I(\U400_ADDRESS_DECODE.m71_amZ0Z_1 ));
    IoInMux I__334 (
            .O(N__2995),
            .I(N__2992));
    LocalMux I__333 (
            .O(N__2992),
            .I(N__2989));
    Odrv12 I__332 (
            .O(N__2989),
            .I(WEn_c));
    IoInMux I__331 (
            .O(N__2986),
            .I(N__2983));
    LocalMux I__330 (
            .O(N__2983),
            .I(N__2980));
    Odrv12 I__329 (
            .O(N__2980),
            .I(RASn_c));
    InMux I__328 (
            .O(N__2977),
            .I(N__2974));
    LocalMux I__327 (
            .O(N__2974),
            .I(N__2971));
    Span4Mux_h I__326 (
            .O(N__2971),
            .I(N__2968));
    Odrv4 I__325 (
            .O(N__2968),
            .I(A_c_30));
    InMux I__324 (
            .O(N__2965),
            .I(N__2962));
    LocalMux I__323 (
            .O(N__2962),
            .I(N__2959));
    Span4Mux_h I__322 (
            .O(N__2959),
            .I(N__2956));
    Odrv4 I__321 (
            .O(N__2956),
            .I(A_c_29));
    CascadeMux I__320 (
            .O(N__2953),
            .I(N__2950));
    InMux I__319 (
            .O(N__2950),
            .I(N__2947));
    LocalMux I__318 (
            .O(N__2947),
            .I(A_c_28));
    InMux I__317 (
            .O(N__2944),
            .I(N__2941));
    LocalMux I__316 (
            .O(N__2941),
            .I(N__2938));
    Odrv4 I__315 (
            .O(N__2938),
            .I(\U400_ADDRESS_DECODE.m2Z0Z_1 ));
    CascadeMux I__314 (
            .O(N__2935),
            .I(\U400_ADDRESS_DECODE.N_185_cascade_ ));
    InMux I__313 (
            .O(N__2932),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_2 ));
    InMux I__312 (
            .O(N__2929),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_3 ));
    InMux I__311 (
            .O(N__2926),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_4 ));
    InMux I__310 (
            .O(N__2923),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_5 ));
    InMux I__309 (
            .O(N__2920),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_6 ));
    InMux I__308 (
            .O(N__2917),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_7 ));
    InMux I__307 (
            .O(N__2914),
            .I(N__2910));
    InMux I__306 (
            .O(N__2913),
            .I(N__2907));
    LocalMux I__305 (
            .O(N__2910),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__304 (
            .O(N__2907),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__303 (
            .O(N__2902),
            .I(N__2898));
    InMux I__302 (
            .O(N__2901),
            .I(N__2895));
    LocalMux I__301 (
            .O(N__2898),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__300 (
            .O(N__2895),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__299 (
            .O(N__2890),
            .I(N__2886));
    InMux I__298 (
            .O(N__2889),
            .I(N__2883));
    LocalMux I__297 (
            .O(N__2886),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__296 (
            .O(N__2883),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__295 (
            .O(N__2878),
            .I(N__2874));
    InMux I__294 (
            .O(N__2877),
            .I(N__2871));
    LocalMux I__293 (
            .O(N__2874),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ));
    LocalMux I__292 (
            .O(N__2871),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ));
    InMux I__291 (
            .O(N__2866),
            .I(N__2862));
    InMux I__290 (
            .O(N__2865),
            .I(N__2859));
    LocalMux I__289 (
            .O(N__2862),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__288 (
            .O(N__2859),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ));
    CascadeMux I__287 (
            .O(N__2854),
            .I(\U400_SDRAM.un1_REFRESH_COUNTERlt7_0_cascade_ ));
    InMux I__286 (
            .O(N__2851),
            .I(N__2847));
    InMux I__285 (
            .O(N__2850),
            .I(N__2844));
    LocalMux I__284 (
            .O(N__2847),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__283 (
            .O(N__2844),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ));
    IoInMux I__282 (
            .O(N__2839),
            .I(N__2836));
    LocalMux I__281 (
            .O(N__2836),
            .I(N__2833));
    Odrv12 I__280 (
            .O(N__2833),
            .I(CASn_c));
    InMux I__279 (
            .O(N__2830),
            .I(N__2827));
    LocalMux I__278 (
            .O(N__2827),
            .I(A_c_31));
    InMux I__277 (
            .O(N__2824),
            .I(N__2821));
    LocalMux I__276 (
            .O(N__2821),
            .I(N__2818));
    Span4Mux_s1_v I__275 (
            .O(N__2818),
            .I(N__2815));
    Odrv4 I__274 (
            .O(N__2815),
            .I(A_c_27));
    InMux I__273 (
            .O(N__2812),
            .I(N__2808));
    InMux I__272 (
            .O(N__2811),
            .I(N__2805));
    LocalMux I__271 (
            .O(N__2808),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__270 (
            .O(N__2805),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ));
    CascadeMux I__269 (
            .O(N__2800),
            .I(N__2795));
    InMux I__268 (
            .O(N__2799),
            .I(N__2792));
    InMux I__267 (
            .O(N__2798),
            .I(N__2789));
    InMux I__266 (
            .O(N__2795),
            .I(N__2786));
    LocalMux I__265 (
            .O(N__2792),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ));
    LocalMux I__264 (
            .O(N__2789),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ));
    LocalMux I__263 (
            .O(N__2786),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ));
    InMux I__262 (
            .O(N__2779),
            .I(N__2776));
    LocalMux I__261 (
            .O(N__2776),
            .I(\U400_SDRAM.REFRESH_COUNTERZ0Z_2 ));
    InMux I__260 (
            .O(N__2773),
            .I(\U400_SDRAM.un3_REFRESH_COUNTER_cry_1 ));
    IoInMux I__259 (
            .O(N__2770),
            .I(N__2767));
    LocalMux I__258 (
            .O(N__2767),
            .I(N__2764));
    IoSpan4Mux I__257 (
            .O(N__2764),
            .I(N__2761));
    Span4Mux_s3_h I__256 (
            .O(N__2761),
            .I(N__2758));
    Span4Mux_h I__255 (
            .O(N__2758),
            .I(N__2755));
    Span4Mux_h I__254 (
            .O(N__2755),
            .I(N__2752));
    Span4Mux_v I__253 (
            .O(N__2752),
            .I(N__2749));
    Odrv4 I__252 (
            .O(N__2749),
            .I(CLK40_ibuf_gb_io_gb_input));
    INV \INVU400_SDRAM.MA_nesr_2C  (
            .O(\INVU400_SDRAM.MA_nesr_2C_net ),
            .I(N__5248));
    INV \INVU400_SDRAM.MA_nesr_1C  (
            .O(\INVU400_SDRAM.MA_nesr_1C_net ),
            .I(N__5247));
    INV \INVU400_SDRAM.SDRAM_CONFIGUREDC  (
            .O(\INVU400_SDRAM.SDRAM_CONFIGUREDC_net ),
            .I(N__5241));
    INV \INVU400_SDRAM.MA_nesr_10C  (
            .O(\INVU400_SDRAM.MA_nesr_10C_net ),
            .I(N__5244));
    INV \INVU400_SDRAM.SDRAM_COUNTER_0C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_0C_net ),
            .I(N__5237));
    INV \INVU400_SDRAM.BANK1C  (
            .O(\INVU400_SDRAM.BANK1C_net ),
            .I(N__5240));
    INV \INVU400_SDRAM.CS1_ENC  (
            .O(\INVU400_SDRAM.CS1_ENC_net ),
            .I(N__5224));
    INV \INVU400_SDRAM.WRITE_CYCLEC  (
            .O(\INVU400_SDRAM.WRITE_CYCLEC_net ),
            .I(N__5233));
    INV \INVU400_SDRAM.MA_nesr_12C  (
            .O(\INVU400_SDRAM.MA_nesr_12C_net ),
            .I(N__5239));
    INV \INVU400_SDRAM.CS0_ENC  (
            .O(\INVU400_SDRAM.CS0_ENC_net ),
            .I(N__5227));
    INV \INVU400_SDRAM.SDRAM_CMD_1C  (
            .O(\INVU400_SDRAM.SDRAM_CMD_1C_net ),
            .I(N__5232));
    INV \INVU400_SDRAM.SDRAM_COUNTER_2C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .I(N__5242));
    INV \INVU400_SDRAM.MA_nesr_6C  (
            .O(\INVU400_SDRAM.MA_nesr_6C_net ),
            .I(N__5234));
    INV \INVU400_SDRAM.MA_nesr_7C  (
            .O(\INVU400_SDRAM.MA_nesr_7C_net ),
            .I(N__5229));
    INV \INVU400_SDRAM.SDRAM_CMD_0C  (
            .O(\INVU400_SDRAM.SDRAM_CMD_0C_net ),
            .I(N__5226));
    INV \INVU400_SDRAM.SDRAM_CMD_2C  (
            .O(\INVU400_SDRAM.SDRAM_CMD_2C_net ),
            .I(N__5230));
    INV \INVU400_SDRAM.RAM_CYCLEC  (
            .O(\INVU400_SDRAM.RAM_CYCLEC_net ),
            .I(N__5235));
    INV \INVU400_SDRAM.SDRAM_COUNTER_1C  (
            .O(\INVU400_SDRAM.SDRAM_COUNTER_1C_net ),
            .I(N__5238));
    INV \INVU400_SDRAM.RASnC  (
            .O(\INVU400_SDRAM.RASnC_net ),
            .I(N__5223));
    INV \INVU400_SDRAM.CASnC  (
            .O(\INVU400_SDRAM.CASnC_net ),
            .I(N__5222));
    INV \INVU400_SDRAM.REFRESH_COUNTER_2C  (
            .O(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .I(N__5228));
    INV \INVU400_SDRAM.REFRESH_COUNTER_1C  (
            .O(\INVU400_SDRAM.REFRESH_COUNTER_1C_net ),
            .I(N__5231));
    INV \INVU400_SDRAM.REFRESH_COUNTER_0C  (
            .O(\INVU400_SDRAM.REFRESH_COUNTER_0C_net ),
            .I(N__5225));
    defparam IN_MUX_bfv_2_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_4_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_3_0_));
    ICE_GB CLK40_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__2770),
            .GLOBALBUFFEROUTPUT(CLK40_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__3070),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_1_4_6 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_1_4_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_0_LC_1_4_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_0_LC_1_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2798),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_0C_net ),
            .ce(),
            .sr(N__3699));
    defparam \U400_ADDRESS_DECODE.m2_1_LC_2_1_3 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m2_1_LC_2_1_3 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m2_1_LC_2_1_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U400_ADDRESS_DECODE.m2_1_LC_2_1_3  (
            .in0(_gnd_net_),
            .in1(N__2830),
            .in2(_gnd_net_),
            .in3(N__2824),
            .lcout(\U400_ADDRESS_DECODE.m2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_2_3_7 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_2_3_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_1_LC_2_3_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_1_LC_2_3_7  (
            .in0(_gnd_net_),
            .in1(N__2799),
            .in2(_gnd_net_),
            .in3(N__2812),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_1C_net ),
            .ce(),
            .sr(N__3700));
    defparam \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_2_4_0 .C_ON=1'b1;
    defparam \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_2_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_2_4_0  (
            .in0(_gnd_net_),
            .in1(N__2811),
            .in2(N__2800),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_4_0_),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_2_4_1 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_2_4_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_2_LC_2_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_2_LC_2_4_1  (
            .in0(_gnd_net_),
            .in1(N__2779),
            .in2(_gnd_net_),
            .in3(N__2773),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_1 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_2 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3695));
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_2_4_2 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_2_4_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_3_LC_2_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_3_LC_2_4_2  (
            .in0(_gnd_net_),
            .in1(N__2890),
            .in2(_gnd_net_),
            .in3(N__2932),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_2 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_3 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3695));
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_2_4_3 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_2_4_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_4_LC_2_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_4_LC_2_4_3  (
            .in0(_gnd_net_),
            .in1(N__2902),
            .in2(_gnd_net_),
            .in3(N__2929),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_3 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_4 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3695));
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_2_4_4 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_2_4_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_5_LC_2_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_5_LC_2_4_4  (
            .in0(_gnd_net_),
            .in1(N__2914),
            .in2(_gnd_net_),
            .in3(N__2926),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_4 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_5 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3695));
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_2_4_5 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_2_4_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_6_LC_2_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_6_LC_2_4_5  (
            .in0(_gnd_net_),
            .in1(N__2851),
            .in2(_gnd_net_),
            .in3(N__2923),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_5 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_6 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3695));
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_2_4_6 .C_ON=1'b1;
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_2_4_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_7_LC_2_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_7_LC_2_4_6  (
            .in0(_gnd_net_),
            .in1(N__2866),
            .in2(_gnd_net_),
            .in3(N__2920),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(\U400_SDRAM.un3_REFRESH_COUNTER_cry_6 ),
            .carryout(\U400_SDRAM.un3_REFRESH_COUNTER_cry_7 ),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3695));
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_2_4_7 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_2_4_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.REFRESH_COUNTER_8_LC_2_4_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_8_LC_2_4_7  (
            .in0(_gnd_net_),
            .in1(N__2878),
            .in2(_gnd_net_),
            .in3(N__2917),
            .lcout(\U400_SDRAM.REFRESH_COUNTERZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.REFRESH_COUNTER_2C_net ),
            .ce(),
            .sr(N__3695));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNILA301_3_LC_2_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNILA301_3_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNILA301_3_LC_2_5_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNILA301_3_LC_2_5_1  (
            .in0(N__2913),
            .in1(N__2901),
            .in2(_gnd_net_),
            .in3(N__2889),
            .lcout(),
            .ltout(\U400_SDRAM.un1_REFRESH_COUNTERlt7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_2_5_2 .C_ON=1'b0;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_2_5_2 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_2_5_2  (
            .in0(N__2877),
            .in1(N__2865),
            .in2(N__2854),
            .in3(N__2850),
            .lcout(U400_SDRAM_SDRAM_CMD11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CASn_LC_2_9_2 .C_ON=1'b0;
    defparam \U400_SDRAM.CASn_LC_2_9_2 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CASn_LC_2_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.CASn_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6388),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CASnC_net ),
            .ce(),
            .sr(N__6730));
    defparam \U400_SDRAM.WEn_LC_2_9_5 .C_ON=1'b0;
    defparam \U400_SDRAM.WEn_LC_2_9_5 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.WEn_LC_2_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.WEn_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6289),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CASnC_net ),
            .ce(),
            .sr(N__6730));
    defparam \U400_SDRAM.RASn_LC_2_10_3 .C_ON=1'b0;
    defparam \U400_SDRAM.RASn_LC_2_10_3 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.RASn_LC_2_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U400_SDRAM.RASn_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5995),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.RASnC_net ),
            .ce(),
            .sr(N__6731));
    defparam \U400_ADDRESS_DECODE.m2_LC_4_1_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m2_LC_4_1_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m2_LC_4_1_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U400_ADDRESS_DECODE.m2_LC_4_1_5  (
            .in0(N__2977),
            .in1(N__2965),
            .in2(N__2953),
            .in3(N__2944),
            .lcout(\U400_ADDRESS_DECODE.N_170_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_4_3_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_4_3_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_1_LC_4_3_3 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_1_LC_4_3_3  (
            .in0(N__3127),
            .in1(N__4723),
            .in2(N__5418),
            .in3(N__3222),
            .lcout(U400_SDRAM_SDRAM_COUNTER_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_1C_net ),
            .ce(N__4502),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_4_3_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_4_3_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_3_LC_4_3_7 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_3_LC_4_3_7  (
            .in0(N__3115),
            .in1(N__4724),
            .in2(N__5419),
            .in3(N__3223),
            .lcout(U400_SDRAM_SDRAM_COUNTER_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_1C_net ),
            .ce(N__4502),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_LC_4_4_6 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_LC_4_4_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.RAM_CYCLE_LC_4_4_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_LC_4_4_6  (
            .in0(N__5809),
            .in1(N__3221),
            .in2(N__3433),
            .in3(N__3016),
            .lcout(U400_SDRAM_RAM_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.RAM_CYCLEC_net ),
            .ce(),
            .sr(N__6736));
    defparam \U400_ADDRESS_DECODE.SDRAM_COUNTERe_0_i_LC_4_4_7 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.SDRAM_COUNTERe_0_i_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.SDRAM_COUNTERe_0_i_LC_4_4_7 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U400_ADDRESS_DECODE.SDRAM_COUNTERe_0_i_LC_4_4_7  (
            .in0(N__5806),
            .in1(N__3596),
            .in2(N__3363),
            .in3(N__3325),
            .lcout(U400_SDRAM_SDRAM_COUNTERe_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m36_e_LC_4_5_1 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m36_e_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m36_e_LC_4_5_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U400_ADDRESS_DECODE.m36_e_LC_4_5_1  (
            .in0(_gnd_net_),
            .in1(N__4055),
            .in2(_gnd_net_),
            .in3(N__4144),
            .lcout(\U400_ADDRESS_DECODE.N_185 ),
            .ltout(\U400_ADDRESS_DECODE.N_185_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m71_am_1_LC_4_5_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m71_am_1_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m71_am_1_LC_4_5_2 .LUT_INIT=16'b0100010111011111;
    LogicCell40 \U400_ADDRESS_DECODE.m71_am_1_LC_4_5_2  (
            .in0(N__5000),
            .in1(N__3826),
            .in2(N__2935),
            .in3(N__3970),
            .lcout(\U400_ADDRESS_DECODE.m71_amZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m45_LC_4_5_3 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m45_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m45_LC_4_5_3 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \U400_ADDRESS_DECODE.m45_LC_4_5_3  (
            .in0(N__3971),
            .in1(N__5001),
            .in2(N__3848),
            .in3(N__4818),
            .lcout(\U400_ADDRESS_DECODE.N_46_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m19_LC_4_5_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m19_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m19_LC_4_5_4 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \U400_ADDRESS_DECODE.m19_LC_4_5_4  (
            .in0(N__4819),
            .in1(N__5003),
            .in2(N__4366),
            .in3(N__3830),
            .lcout(\U400_ADDRESS_DECODE.N_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m84_bm_LC_4_5_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m84_bm_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m84_bm_LC_4_5_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U400_ADDRESS_DECODE.m84_bm_LC_4_5_5  (
            .in0(N__3558),
            .in1(N__3990),
            .in2(_gnd_net_),
            .in3(N__3637),
            .lcout(\U400_ADDRESS_DECODE.m84_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m84_am_LC_4_5_6 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m84_am_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m84_am_LC_4_5_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U400_ADDRESS_DECODE.m84_am_LC_4_5_6  (
            .in0(N__4145),
            .in1(N__3597),
            .in2(_gnd_net_),
            .in3(N__4061),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.m84_amZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m84_ns_LC_4_5_7 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m84_ns_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m84_ns_LC_4_5_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \U400_ADDRESS_DECODE.m84_ns_LC_4_5_7  (
            .in0(N__4655),
            .in1(_gnd_net_),
            .in2(N__3025),
            .in3(N__3022),
            .lcout(N_85_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m71_bm_LC_4_6_0 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m71_bm_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m71_bm_LC_4_6_0 .LUT_INIT=16'b0001000100010101;
    LogicCell40 \U400_ADDRESS_DECODE.m71_bm_LC_4_6_0  (
            .in0(N__4833),
            .in1(N__3847),
            .in2(N__5010),
            .in3(N__3977),
            .lcout(\U400_ADDRESS_DECODE.m71_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m46_LC_4_6_1 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m46_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m46_LC_4_6_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U400_ADDRESS_DECODE.m46_LC_4_6_1  (
            .in0(N__3875),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4989),
            .lcout(\U400_ADDRESS_DECODE.N_47_0 ),
            .ltout(\U400_ADDRESS_DECODE.N_47_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m56_am_LC_4_6_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m56_am_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m56_am_LC_4_6_2 .LUT_INIT=16'b0101000010101010;
    LogicCell40 \U400_ADDRESS_DECODE.m56_am_LC_4_6_2  (
            .in0(N__3010),
            .in1(_gnd_net_),
            .in2(N__3004),
            .in3(N__4652),
            .lcout(\U400_ADDRESS_DECODE.m56_amZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m71_am_LC_4_6_3 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m71_am_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m71_am_LC_4_6_3 .LUT_INIT=16'b0011000001010101;
    LogicCell40 \U400_ADDRESS_DECODE.m71_am_LC_4_6_3  (
            .in0(N__4857),
            .in1(N__3324),
            .in2(N__3880),
            .in3(N__3001),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.m71_amZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m71_ns_LC_4_6_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m71_ns_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m71_ns_LC_4_6_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \U400_ADDRESS_DECODE.m71_ns_LC_4_6_4  (
            .in0(_gnd_net_),
            .in1(N__4653),
            .in2(N__3100),
            .in3(N__3097),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.N_72_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m72_LC_4_6_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m72_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m72_LC_4_6_5 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \U400_ADDRESS_DECODE.m72_LC_4_6_5  (
            .in0(_gnd_net_),
            .in1(N__5807),
            .in2(N__3091),
            .in3(N__5856),
            .lcout(N_73_0),
            .ltout(N_73_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_4_6_6 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_4_6_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_2_LC_4_6_6 .LUT_INIT=16'b0101110111111101;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_2_LC_4_6_6  (
            .in0(N__6555),
            .in1(N__5941),
            .in2(N__3088),
            .in3(N__3079),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m56_ns_LC_4_6_7 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m56_ns_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m56_ns_LC_4_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U400_ADDRESS_DECODE.m56_ns_LC_4_6_7  (
            .in0(N__3085),
            .in1(N__3331),
            .in2(_gnd_net_),
            .in3(N__5808),
            .lcout(N_57_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m6_LC_4_7_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m6_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m6_LC_4_7_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U400_ADDRESS_DECODE.m6_LC_4_7_4  (
            .in0(N__4853),
            .in1(N__5002),
            .in2(_gnd_net_),
            .in3(N__3846),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.N_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m63_ns_1_LC_4_7_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m63_ns_1_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m63_ns_1_LC_4_7_5 .LUT_INIT=16'b0001100101001100;
    LogicCell40 \U400_ADDRESS_DECODE.m63_ns_1_LC_4_7_5  (
            .in0(N__4348),
            .in1(N__3991),
            .in2(N__3073),
            .in3(N__3640),
            .lcout(\U400_ADDRESS_DECODE.m63_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_0_LC_4_7_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_0_LC_4_7_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_0_LC_4_7_7 .LUT_INIT=16'b1100111110101111;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_0_LC_4_7_7  (
            .in0(N__6256),
            .in1(N__3292),
            .in2(N__6598),
            .in3(N__3385),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_4_8_7.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_4_8_7.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_4_8_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_4_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6611),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_7_LC_4_12_4 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_7_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_7_LC_4_12_4 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_7_LC_4_12_4  (
            .in0(N__3061),
            .in1(N__5978),
            .in2(N__3052),
            .in3(N__6858),
            .lcout(MA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_7C_net ),
            .ce(N__6802),
            .sr(N__6735));
    defparam \U400_SDRAM.MA_nesr_8_LC_4_12_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_8_LC_4_12_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_8_LC_4_12_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \U400_SDRAM.MA_nesr_8_LC_4_12_7  (
            .in0(N__6859),
            .in1(N__5994),
            .in2(N__3208),
            .in3(N__3193),
            .lcout(MA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_7C_net ),
            .ce(N__6802),
            .sr(N__6735));
    defparam \U400_SDRAM.MA_nesr_6_LC_4_14_0 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_6_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_6_LC_4_14_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_6_LC_4_14_0  (
            .in0(N__3163),
            .in1(N__6006),
            .in2(N__3154),
            .in3(N__6852),
            .lcout(MA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_6C_net ),
            .ce(N__6801),
            .sr(N__6739));
    defparam \U400_ADDRESS_DECODE.m133_0_LC_5_3_0 .C_ON=1'b1;
    defparam \U400_ADDRESS_DECODE.m133_0_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m133_0_LC_5_3_0 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \U400_ADDRESS_DECODE.m133_0_LC_5_3_0  (
            .in0(N__6639),
            .in1(N__4646),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U400_ADDRESS_DECODE.m133Z0Z_0 ),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_3_1 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_3_1  (
            .in0(_gnd_net_),
            .in1(N__3822),
            .in2(_gnd_net_),
            .in3(N__3121),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_1 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_5_3_2 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_5_3_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_2_LC_5_3_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_2_LC_5_3_2  (
            .in0(N__4719),
            .in1(N__4983),
            .in2(_gnd_net_),
            .in3(N__3118),
            .lcout(U400_SDRAM_SDRAM_COUNTER_2),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_2 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__4503),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_5_3_3 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_5_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_5_3_3  (
            .in0(_gnd_net_),
            .in1(N__3999),
            .in2(_gnd_net_),
            .in3(N__3109),
            .lcout(\U400_SDRAM.SDRAM_COUNTER_s_3 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_5_3_4 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_5_3_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_4_LC_5_3_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_4_LC_5_3_4  (
            .in0(N__4720),
            .in1(N__3241),
            .in2(_gnd_net_),
            .in3(N__3106),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_4 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__4503),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_5_3_5 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_5_3_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_5_LC_5_3_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_5_LC_5_3_5  (
            .in0(N__4731),
            .in1(N__3268),
            .in2(_gnd_net_),
            .in3(N__3103),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_5 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__4503),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_5_3_6 .C_ON=1'b1;
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_5_3_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_6_LC_5_3_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_6_LC_5_3_6  (
            .in0(N__4721),
            .in1(N__3280),
            .in2(_gnd_net_),
            .in3(N__3286),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U400_SDRAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U400_SDRAM.SDRAM_COUNTER_cry_6 ),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__4503),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_5_3_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_5_3_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_7_LC_5_3_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_7_LC_5_3_7  (
            .in0(N__3255),
            .in1(N__4722),
            .in2(_gnd_net_),
            .in3(N__3283),
            .lcout(\U400_SDRAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_2C_net ),
            .ce(N__4503),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m41_bm_LC_5_4_0 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m41_bm_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m41_bm_LC_5_4_0 .LUT_INIT=16'b0000000011111101;
    LogicCell40 \U400_ADDRESS_DECODE.m41_bm_LC_5_4_0  (
            .in0(N__4923),
            .in1(N__3814),
            .in2(N__4364),
            .in3(N__4800),
            .lcout(\U400_ADDRESS_DECODE.m41_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_4_1 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_4_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_4_1  (
            .in0(N__3279),
            .in1(N__3267),
            .in2(N__3256),
            .in3(N__3240),
            .lcout(N_60),
            .ltout(N_60_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m9_LC_5_4_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m9_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m9_LC_5_4_2 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \U400_ADDRESS_DECODE.m9_LC_5_4_2  (
            .in0(_gnd_net_),
            .in1(N__4922),
            .in2(N__3229),
            .in3(N__3813),
            .lcout(\U400_ADDRESS_DECODE.N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m97_LC_5_4_3 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m97_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m97_LC_5_4_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U400_ADDRESS_DECODE.m97_LC_5_4_3  (
            .in0(N__3726),
            .in1(N__4117),
            .in2(_gnd_net_),
            .in3(N__4657),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.N_98_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.N_100_0_i_LC_5_4_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.N_100_0_i_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.N_100_0_i_LC_5_4_4 .LUT_INIT=16'b1111001110111011;
    LogicCell40 \U400_ADDRESS_DECODE.N_100_0_i_LC_5_4_4  (
            .in0(N__4266),
            .in1(N__6635),
            .in2(N__3226),
            .in3(N__5782),
            .lcout(N_100_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m78_LC_5_4_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m78_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m78_LC_5_4_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_ADDRESS_DECODE.m78_LC_5_4_5  (
            .in0(N__4658),
            .in1(N__5802),
            .in2(N__6640),
            .in3(N__3714),
            .lcout(U400_SDRAM_SDRAM_CMD_5_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m41_am_LC_5_4_6 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m41_am_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m41_am_LC_5_4_6 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \U400_ADDRESS_DECODE.m41_am_LC_5_4_6  (
            .in0(N__5801),
            .in1(N__3815),
            .in2(N__4363),
            .in3(N__4801),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.m41_amZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m41_ns_LC_5_4_7 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m41_ns_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m41_ns_LC_5_4_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \U400_ADDRESS_DECODE.m41_ns_LC_5_4_7  (
            .in0(_gnd_net_),
            .in1(N__3934),
            .in2(N__3343),
            .in3(N__3340),
            .lcout(\U400_ADDRESS_DECODE.N_42_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m14_LC_5_5_0 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m14_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m14_LC_5_5_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U400_ADDRESS_DECODE.m14_LC_5_5_0  (
            .in0(N__4796),
            .in1(N__4948),
            .in2(_gnd_net_),
            .in3(N__4003),
            .lcout(\U400_ADDRESS_DECODE.N_15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m5_LC_5_5_1 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m5_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m5_LC_5_5_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U400_ADDRESS_DECODE.m5_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(N__3823),
            .in2(_gnd_net_),
            .in3(N__4795),
            .lcout(\U400_ADDRESS_DECODE.N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m87_ns_1_LC_5_5_3 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m87_ns_1_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m87_ns_1_LC_5_5_3 .LUT_INIT=16'b0001000100011011;
    LogicCell40 \U400_ADDRESS_DECODE.m87_ns_1_LC_5_5_3  (
            .in0(N__4004),
            .in1(N__3635),
            .in2(N__3850),
            .in3(N__4797),
            .lcout(\U400_ADDRESS_DECODE.m87_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m54_0_LC_5_5_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m54_0_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m54_0_LC_5_5_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U400_ADDRESS_DECODE.m54_0_LC_5_5_4  (
            .in0(N__3824),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4949),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.m54Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m56_bm_LC_5_5_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m56_bm_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m56_bm_LC_5_5_5 .LUT_INIT=16'b0011000110010001;
    LogicCell40 \U400_ADDRESS_DECODE.m56_bm_LC_5_5_5  (
            .in0(N__4005),
            .in1(N__4654),
            .in2(N__3334),
            .in3(N__4362),
            .lcout(\U400_ADDRESS_DECODE.m56_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_5_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.RAM_CYCLE_START_LC_5_5_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U400_SDRAM.RAM_CYCLE_START_LC_5_5_6  (
            .in0(N__6606),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3415),
            .lcout(U400_SDRAM_RAM_CYCLE_START),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5236),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m36_LC_5_6_0 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m36_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m36_LC_5_6_0 .LUT_INIT=16'b1000100010001101;
    LogicCell40 \U400_ADDRESS_DECODE.m36_LC_5_6_0  (
            .in0(N__4010),
            .in1(N__3409),
            .in2(N__5011),
            .in3(N__3323),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.N_185_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m43_bm_LC_5_6_1 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m43_bm_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m43_bm_LC_5_6_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \U400_ADDRESS_DECODE.m43_bm_LC_5_6_1  (
            .in0(N__4648),
            .in1(_gnd_net_),
            .in2(N__3307),
            .in3(N__3304),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.m43_bmZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m43_ns_LC_5_6_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m43_ns_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m43_ns_LC_5_6_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \U400_ADDRESS_DECODE.m43_ns_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__5783),
            .in2(N__3295),
            .in3(N__3403),
            .lcout(N_44_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m32_LC_5_6_3 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m32_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m32_LC_5_6_3 .LUT_INIT=16'b0001000010111011;
    LogicCell40 \U400_ADDRESS_DECODE.m32_LC_5_6_3  (
            .in0(N__3825),
            .in1(N__4355),
            .in2(N__4988),
            .in3(N__4831),
            .lcout(\U400_ADDRESS_DECODE.N_33_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m43_am_LC_5_6_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m43_am_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m43_am_LC_5_6_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U400_ADDRESS_DECODE.m43_am_LC_5_6_4  (
            .in0(N__4832),
            .in1(N__4647),
            .in2(N__4018),
            .in3(N__4953),
            .lcout(\U400_ADDRESS_DECODE.m43_amZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m87_ns_LC_5_6_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m87_ns_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m87_ns_LC_5_6_5 .LUT_INIT=16'b1100011011110110;
    LogicCell40 \U400_ADDRESS_DECODE.m87_ns_LC_5_6_5  (
            .in0(N__3397),
            .in1(N__4014),
            .in2(N__4660),
            .in3(N__3559),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.N_88_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m95_ns_LC_5_6_6 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m95_ns_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m95_ns_LC_5_6_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \U400_ADDRESS_DECODE.m95_ns_LC_5_6_6  (
            .in0(N__4156),
            .in1(_gnd_net_),
            .in2(N__3391),
            .in3(N__5784),
            .lcout(),
            .ltout(N_96_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_5_6_7 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CMD_1_LC_5_6_7 .LUT_INIT=16'b1111010111011101;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_1_LC_5_6_7  (
            .in0(N__6612),
            .in1(N__6357),
            .in2(N__3388),
            .in3(N__3384),
            .lcout(\U400_SDRAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CMD_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m63_ns_LC_5_7_0 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m63_ns_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m63_ns_LC_5_7_0 .LUT_INIT=16'b0011011000000110;
    LogicCell40 \U400_ADDRESS_DECODE.m63_ns_LC_5_7_0  (
            .in0(N__3373),
            .in1(N__4017),
            .in2(N__4659),
            .in3(N__3541),
            .lcout(N_48),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m138_LC_5_7_1 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m138_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m138_LC_5_7_1 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \U400_ADDRESS_DECODE.m138_LC_5_7_1  (
            .in0(N__4985),
            .in1(N__3638),
            .in2(N__4347),
            .in3(N__4854),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.N_139_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m141_am_LC_5_7_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m141_am_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m141_am_LC_5_7_2 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \U400_ADDRESS_DECODE.m141_am_LC_5_7_2  (
            .in0(N__4855),
            .in1(N__4986),
            .in2(N__3367),
            .in3(N__4015),
            .lcout(\U400_ADDRESS_DECODE.m141_amZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m133_LC_5_7_3 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m133_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m133_LC_5_7_3 .LUT_INIT=16'b1100000001000000;
    LogicCell40 \U400_ADDRESS_DECODE.m133_LC_5_7_3  (
            .in0(N__5800),
            .in1(N__3598),
            .in2(N__3364),
            .in3(N__4075),
            .lcout(N_190_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m61_LC_5_7_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m61_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m61_LC_5_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U400_ADDRESS_DECODE.m61_LC_5_7_4  (
            .in0(N__3639),
            .in1(N__4325),
            .in2(_gnd_net_),
            .in3(N__3557),
            .lcout(\U400_ADDRESS_DECODE.N_62_0 ),
            .ltout(\U400_ADDRESS_DECODE.N_62_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m141_bm_LC_5_7_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m141_bm_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m141_bm_LC_5_7_5 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \U400_ADDRESS_DECODE.m141_bm_LC_5_7_5  (
            .in0(N__4016),
            .in1(N__5014),
            .in2(N__3535),
            .in3(N__4856),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.m141_bmZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m141_ns_LC_5_7_6 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m141_ns_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m141_ns_LC_5_7_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \U400_ADDRESS_DECODE.m141_ns_LC_5_7_6  (
            .in0(N__4644),
            .in1(_gnd_net_),
            .in2(N__3532),
            .in3(N__3529),
            .lcout(N_142_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS0_EN_LC_5_8_6 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0_EN_LC_5_8_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.CS0_EN_LC_5_8_6 .LUT_INIT=16'b1111101011101110;
    LogicCell40 \U400_SDRAM.CS0_EN_LC_5_8_6  (
            .in0(N__4218),
            .in1(N__4228),
            .in2(N__3523),
            .in3(N__4200),
            .lcout(\U400_SDRAM.CS0_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0_ENC_net ),
            .ce(),
            .sr(N__6732));
    defparam \U400_SDRAM.CS0n_LC_5_8_7 .C_ON=1'b0;
    defparam \U400_SDRAM.CS0n_LC_5_8_7 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CS0n_LC_5_8_7 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \U400_SDRAM.CS0n_LC_5_8_7  (
            .in0(N__5965),
            .in1(N__6367),
            .in2(N__3522),
            .in3(N__6249),
            .lcout(CS0n_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS0_ENC_net ),
            .ce(),
            .sr(N__6732));
    defparam \U400_SDRAM.MA_nesr_12_LC_5_14_2 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_12_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_12_LC_5_14_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.MA_nesr_12_LC_5_14_2  (
            .in0(N__6023),
            .in1(N__6407),
            .in2(N__3490),
            .in3(N__6306),
            .lcout(MA_c_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_12C_net ),
            .ce(N__6790),
            .sr(N__6740));
    defparam \U400_SDRAM.MA_nesr_9_LC_5_14_6 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_9_LC_5_14_6 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_9_LC_5_14_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U400_SDRAM.MA_nesr_9_LC_5_14_6  (
            .in0(N__6024),
            .in1(N__6408),
            .in2(N__3460),
            .in3(N__6307),
            .lcout(MA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_12C_net ),
            .ce(N__6790),
            .sr(N__6740));
    defparam \U400_ADDRESS_DECODE.m165_ns_LC_6_4_0 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m165_ns_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m165_ns_LC_6_4_0 .LUT_INIT=16'b1111011110100010;
    LogicCell40 \U400_ADDRESS_DECODE.m165_ns_LC_6_4_0  (
            .in0(N__3432),
            .in1(N__5496),
            .in2(N__3670),
            .in3(N__3649),
            .lcout(U400_SDRAM_RAM_CYCLE_START_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m7_LC_6_4_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m7_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m7_LC_6_4_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U400_ADDRESS_DECODE.m7_LC_6_4_2  (
            .in0(N__3855),
            .in1(N__4820),
            .in2(N__4984),
            .in3(N__4006),
            .lcout(\U400_ADDRESS_DECODE.N_8_0 ),
            .ltout(\U400_ADDRESS_DECODE.N_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m11_LC_6_4_3 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m11_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m11_LC_6_4_3 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U400_ADDRESS_DECODE.m11_LC_6_4_3  (
            .in0(N__4007),
            .in1(N__4607),
            .in2(N__3703),
            .in3(N__3636),
            .lcout(\U400_ADDRESS_DECODE.N_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCA2_LC_6_4_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCA2_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCA2_LC_6_4_4 .LUT_INIT=16'b0111001100110011;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCA2_LC_6_4_4  (
            .in0(N__4608),
            .in1(N__6626),
            .in2(N__5805),
            .in3(N__4100),
            .lcout(\U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m165_ns_1_LC_6_4_7 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m165_ns_1_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m165_ns_1_LC_6_4_7 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \U400_ADDRESS_DECODE.m165_ns_1_LC_6_4_7  (
            .in0(N__6625),
            .in1(N__3666),
            .in2(N__6687),
            .in3(N__4150),
            .lcout(\U400_ADDRESS_DECODE.m165_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m12_LC_6_5_0 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m12_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m12_LC_6_5_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U400_ADDRESS_DECODE.m12_LC_6_5_0  (
            .in0(N__3851),
            .in1(N__4000),
            .in2(N__4987),
            .in3(N__4798),
            .lcout(N_13_0),
            .ltout(N_13_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m134_LC_6_5_1 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m134_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m134_LC_6_5_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \U400_ADDRESS_DECODE.m134_LC_6_5_1  (
            .in0(N__4799),
            .in1(N__4602),
            .in2(N__3643),
            .in3(N__4947),
            .lcout(\U400_ADDRESS_DECODE.N_135_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m64_LC_6_5_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m64_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m64_LC_6_5_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U400_ADDRESS_DECODE.m64_LC_6_5_2  (
            .in0(N__4601),
            .in1(N__4002),
            .in2(_gnd_net_),
            .in3(N__3626),
            .lcout(N_65_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m75_LC_6_5_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m75_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m75_LC_6_5_4 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \U400_ADDRESS_DECODE.m75_LC_6_5_4  (
            .in0(N__4147),
            .in1(_gnd_net_),
            .in2(N__4078),
            .in3(N__3580),
            .lcout(\U400_ADDRESS_DECODE.N_179_mux ),
            .ltout(\U400_ADDRESS_DECODE.N_179_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m77_LC_6_5_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m77_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m77_LC_6_5_5 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \U400_ADDRESS_DECODE.m77_LC_6_5_5  (
            .in0(_gnd_net_),
            .in1(N__4603),
            .in2(N__3562),
            .in3(N__5803),
            .lcout(U400_SDRAM_SDRAM_CMD_1_sqmuxa_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m94_am_1_LC_6_5_7 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m94_am_1_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m94_am_1_LC_6_5_7 .LUT_INIT=16'b0000101100001010;
    LogicCell40 \U400_ADDRESS_DECODE.m94_am_1_LC_6_5_7  (
            .in0(N__4001),
            .in1(N__4071),
            .in2(N__3856),
            .in3(N__4146),
            .lcout(\U400_ADDRESS_DECODE.m94_amZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m94_am_LC_6_6_0 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m94_am_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m94_am_LC_6_6_0 .LUT_INIT=16'b1011000100110010;
    LogicCell40 \U400_ADDRESS_DECODE.m94_am_LC_6_6_0  (
            .in0(N__4009),
            .in1(N__4848),
            .in2(N__5012),
            .in3(N__4165),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.m94_amZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m94_ns_LC_6_6_1 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m94_ns_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m94_ns_LC_6_6_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \U400_ADDRESS_DECODE.m94_ns_LC_6_6_1  (
            .in0(N__4631),
            .in1(_gnd_net_),
            .in2(N__4159),
            .in3(N__3862),
            .lcout(\U400_ADDRESS_DECODE.N_95_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m145_ns_1_LC_6_6_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m145_ns_1_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m145_ns_1_LC_6_6_2 .LUT_INIT=16'b0001110100001111;
    LogicCell40 \U400_ADDRESS_DECODE.m145_ns_1_LC_6_6_2  (
            .in0(N__4115),
            .in1(N__4076),
            .in2(N__4101),
            .in3(N__4148),
            .lcout(\U400_ADDRESS_DECODE.m145_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m20_am_LC_6_6_3 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m20_am_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m20_am_LC_6_6_3 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \U400_ADDRESS_DECODE.m20_am_LC_6_6_3  (
            .in0(N__4149),
            .in1(N__4116),
            .in2(N__4102),
            .in3(N__4077),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.m20_amZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m20_ns_LC_6_6_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m20_ns_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m20_ns_LC_6_6_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \U400_ADDRESS_DECODE.m20_ns_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(N__4630),
            .in2(N__4021),
            .in3(N__3742),
            .lcout(\U400_ADDRESS_DECODE.N_21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m94_bm_LC_6_6_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m94_bm_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m94_bm_LC_6_6_5 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \U400_ADDRESS_DECODE.m94_bm_LC_6_6_5  (
            .in0(N__4849),
            .in1(N__4008),
            .in2(_gnd_net_),
            .in3(N__3879),
            .lcout(\U400_ADDRESS_DECODE.m94_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m20_bm_LC_6_6_6 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m20_bm_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m20_bm_LC_6_6_6 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \U400_ADDRESS_DECODE.m20_bm_LC_6_6_6  (
            .in0(N__4996),
            .in1(N__3849),
            .in2(N__4365),
            .in3(N__4847),
            .lcout(\U400_ADDRESS_DECODE.m20_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m153_LC_6_6_7 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m153_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m153_LC_6_6_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U400_ADDRESS_DECODE.m153_LC_6_6_7  (
            .in0(N__5804),
            .in1(N__3736),
            .in2(N__4656),
            .in3(N__3715),
            .lcout(U400_SDRAM_un1_SDRAM_COUNTER59_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.WRITE_CYCLE_LC_6_7_5 .C_ON=1'b0;
    defparam \U400_SDRAM.WRITE_CYCLE_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.WRITE_CYCLE_LC_6_7_5 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U400_SDRAM.WRITE_CYCLE_LC_6_7_5  (
            .in0(N__4378),
            .in1(N__4329),
            .in2(_gnd_net_),
            .in3(N__5029),
            .lcout(U400_SDRAM_WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.WRITE_CYCLEC_net ),
            .ce(),
            .sr(N__6733));
    defparam \U400_SDRAM.TACK_LC_6_7_7 .C_ON=1'b0;
    defparam \U400_SDRAM.TACK_LC_6_7_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TACK_LC_6_7_7 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \U400_SDRAM.TACK_LC_6_7_7  (
            .in0(N__4398),
            .in1(N__4282),
            .in2(N__5788),
            .in3(N__4276),
            .lcout(U400_SDRAM_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.WRITE_CYCLEC_net ),
            .ce(),
            .sr(N__6733));
    defparam \U400_ADDRESS_DECODE.m22_LC_6_8_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m22_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m22_LC_6_8_2 .LUT_INIT=16'b0001000010110000;
    LogicCell40 \U400_ADDRESS_DECODE.m22_LC_6_8_2  (
            .in0(N__5787),
            .in1(N__4270),
            .in2(N__6610),
            .in3(N__4255),
            .lcout(N_23_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m137_LC_6_8_3 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m137_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m137_LC_6_8_3 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \U400_ADDRESS_DECODE.m137_LC_6_8_3  (
            .in0(N__5786),
            .in1(N__4476),
            .in2(N__4246),
            .in3(N__5852),
            .lcout(N_138_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_6_8_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_8_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_8_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m136_LC_6_8_7 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m136_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m136_LC_6_8_7 .LUT_INIT=16'b0010000001110000;
    LogicCell40 \U400_ADDRESS_DECODE.m136_LC_6_8_7  (
            .in0(N__5785),
            .in1(N__4475),
            .in2(N__4245),
            .in3(N__5851),
            .lcout(N_137_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.CS1_EN_LC_6_9_1 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1_EN_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.CS1_EN_LC_6_9_1 .LUT_INIT=16'b1111101011101110;
    LogicCell40 \U400_SDRAM.CS1_EN_LC_6_9_1  (
            .in0(N__4222),
            .in1(N__4207),
            .in2(N__4189),
            .in3(N__4201),
            .lcout(\U400_SDRAM.CS1_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS1_ENC_net ),
            .ce(),
            .sr(N__6734));
    defparam \U400_SDRAM.CS1n_LC_6_9_3 .C_ON=1'b0;
    defparam \U400_SDRAM.CS1n_LC_6_9_3 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.CS1n_LC_6_9_3 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \U400_SDRAM.CS1n_LC_6_9_3  (
            .in0(N__6371),
            .in1(N__5979),
            .in2(N__4188),
            .in3(N__6288),
            .lcout(CS1n_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.CS1_ENC_net ),
            .ce(),
            .sr(N__6734));
    defparam \U400_SDRAM.TA_COUNTER_4_LC_7_4_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_4_LC_7_4_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_4_LC_7_4_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_4_LC_7_4_1  (
            .in0(_gnd_net_),
            .in1(N__6608),
            .in2(_gnd_net_),
            .in3(N__5134),
            .lcout(U400_SDRAM_TA_COUNTER_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5245),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_5_LC_7_4_2 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_5_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_5_LC_7_4_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_5_LC_7_4_2  (
            .in0(N__6609),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4452),
            .lcout(U400_SDRAM_TA_COUNTER_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5245),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m111_e_LC_7_4_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m111_e_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m111_e_LC_7_4_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U400_ADDRESS_DECODE.m111_e_LC_7_4_4  (
            .in0(_gnd_net_),
            .in1(N__4448),
            .in2(_gnd_net_),
            .in3(N__4436),
            .lcout(N_174),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m102_LC_7_4_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m102_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m102_LC_7_4_5 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \U400_ADDRESS_DECODE.m102_LC_7_4_5  (
            .in0(N__4437),
            .in1(_gnd_net_),
            .in2(N__4453),
            .in3(N__5893),
            .lcout(U400_SDRAM_TA_OUT_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_1_LC_7_5_0 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_1_LC_7_5_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_1_LC_7_5_0 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_1_LC_7_5_0  (
            .in0(N__4402),
            .in1(_gnd_net_),
            .in2(N__4420),
            .in3(N__6603),
            .lcout(U400_SDRAM_TA_COUNTER_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5243),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_2_LC_7_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_2_LC_7_5_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_2_LC_7_5_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_2_LC_7_5_1  (
            .in0(N__6604),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4438),
            .lcout(U400_SDRAM_TA_COUNTER_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5243),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m112_LC_7_5_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m112_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m112_LC_7_5_2 .LUT_INIT=16'b0001111100001111;
    LogicCell40 \U400_ADDRESS_DECODE.m112_LC_7_5_2  (
            .in0(N__4401),
            .in1(N__5133),
            .in2(N__6624),
            .in3(N__5292),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.N_177_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_0_LC_7_5_3 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_0_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_0_LC_7_5_3 .LUT_INIT=16'b1101110011111110;
    LogicCell40 \U400_SDRAM.TA_COUNTER_0_LC_7_5_3  (
            .in0(N__5148),
            .in1(N__5161),
            .in2(N__4423),
            .in3(N__5863),
            .lcout(U400_SDRAM_TA_COUNTER_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5243),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m26_LC_7_5_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m26_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m26_LC_7_5_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U400_ADDRESS_DECODE.m26_LC_7_5_4  (
            .in0(N__4400),
            .in1(_gnd_net_),
            .in2(N__4419),
            .in3(_gnd_net_),
            .lcout(U400_SDRAM_N_252_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_RNIF6C61_0_LC_7_5_5 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_RNIF6C61_0_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_COUNTER_RNIF6C61_0_LC_7_5_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_RNIF6C61_0_LC_7_5_5  (
            .in0(N__6605),
            .in1(N__4412),
            .in2(_gnd_net_),
            .in3(N__4399),
            .lcout(\U400_SDRAM.N_252_0_0 ),
            .ltout(\U400_SDRAM.N_252_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_EN_i_RNO_0_LC_7_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_EN_i_RNO_0_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.TA_EN_i_RNO_0_LC_7_5_6 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \U400_SDRAM.TA_EN_i_RNO_0_LC_7_5_6  (
            .in0(N__5160),
            .in1(N__5144),
            .in2(N__5152),
            .in3(N__5887),
            .lcout(\U400_SDRAM.N_252_0_0_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_COUNTER_3_LC_7_5_7 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_COUNTER_3_LC_7_5_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.TA_COUNTER_3_LC_7_5_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U400_SDRAM.TA_COUNTER_3_LC_7_5_7  (
            .in0(N__5888),
            .in1(_gnd_net_),
            .in2(N__5149),
            .in3(N__6602),
            .lcout(U400_SDRAM_TA_COUNTER_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5243),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.BANK1_LC_7_6_0 .C_ON=1'b0;
    defparam \U400_SDRAM.BANK1_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BANK1_LC_7_6_0 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \U400_SDRAM.BANK1_LC_7_6_0  (
            .in0(N__5062),
            .in1(N__5091),
            .in2(N__5122),
            .in3(N__4600),
            .lcout(BANK1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK1C_net ),
            .ce(),
            .sr(N__6737));
    defparam \U400_SDRAM.BANK0_LC_7_6_1 .C_ON=1'b0;
    defparam \U400_SDRAM.BANK0_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BANK0_LC_7_6_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \U400_SDRAM.BANK0_LC_7_6_1  (
            .in0(N__5040),
            .in1(N__4599),
            .in2(N__5080),
            .in3(N__5061),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK1C_net ),
            .ce(),
            .sr(N__6737));
    defparam \U400_SDRAM.BURST_LC_7_6_2 .C_ON=1'b0;
    defparam \U400_SDRAM.BURST_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.BURST_LC_7_6_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U400_SDRAM.BURST_LC_7_6_2  (
            .in0(N__5473),
            .in1(N__5892),
            .in2(N__5581),
            .in3(N__5025),
            .lcout(U400_SDRAM_BURST),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.BANK1C_net ),
            .ce(),
            .sr(N__6737));
    defparam \U400_ADDRESS_DECODE.m145_ns_LC_7_7_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m145_ns_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m145_ns_LC_7_7_2 .LUT_INIT=16'b0010000000101111;
    LogicCell40 \U400_ADDRESS_DECODE.m145_ns_LC_7_7_2  (
            .in0(N__5013),
            .in1(N__4858),
            .in2(N__4645),
            .in3(N__4738),
            .lcout(\U400_ADDRESS_DECODE.N_146_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_7_7_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_COUNTER_0_LC_7_7_5 .LUT_INIT=16'b0001001011011110;
    LogicCell40 \U400_SDRAM.SDRAM_COUNTER_0_LC_7_7_5  (
            .in0(N__4598),
            .in1(N__4732),
            .in2(N__4677),
            .in3(N__5380),
            .lcout(U400_SDRAM_SDRAM_COUNTER_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_COUNTER_0C_net ),
            .ce(N__4507),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m149_e_LC_7_8_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m149_e_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m149_e_LC_7_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U400_ADDRESS_DECODE.m149_e_LC_7_8_2  (
            .in0(_gnd_net_),
            .in1(N__5564),
            .in2(_gnd_net_),
            .in3(N__5469),
            .lcout(N_14_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m135_LC_7_8_3 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m135_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m135_LC_7_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U400_ADDRESS_DECODE.m135_LC_7_8_3  (
            .in0(N__5725),
            .in1(N__5846),
            .in2(_gnd_net_),
            .in3(N__4477),
            .lcout(\U400_ADDRESS_DECODE.N_136_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m146_LC_7_8_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m146_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m146_LC_7_8_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U400_ADDRESS_DECODE.m146_LC_7_8_4  (
            .in0(N__5847),
            .in1(N__5726),
            .in2(_gnd_net_),
            .in3(N__5425),
            .lcout(),
            .ltout(\U400_ADDRESS_DECODE.N_147_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m149_LC_7_8_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m149_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m149_LC_7_8_5 .LUT_INIT=16'b1111011111010101;
    LogicCell40 \U400_ADDRESS_DECODE.m149_LC_7_8_5  (
            .in0(N__6580),
            .in1(N__5400),
            .in2(N__5389),
            .in3(N__5386),
            .lcout(N_43),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_10_LC_7_14_0 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_10_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_10_LC_7_14_0 .LUT_INIT=16'b0000100000001010;
    LogicCell40 \U400_SDRAM.MA_nesr_10_LC_7_14_0  (
            .in0(N__6401),
            .in1(N__5374),
            .in2(N__6037),
            .in3(N__6297),
            .lcout(MA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_10C_net ),
            .ce(N__6776),
            .sr(N__6742));
    defparam \U400_SDRAM.MA_nesr_11_LC_7_14_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_11_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_11_LC_7_14_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U400_SDRAM.MA_nesr_11_LC_7_14_7  (
            .in0(N__6298),
            .in1(N__6027),
            .in2(N__5344),
            .in3(N__6402),
            .lcout(MA_c_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_10C_net ),
            .ce(N__6776),
            .sr(N__6742));
    defparam \U400_ADDRESS_DECODE.m3_LC_8_4_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m3_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m3_LC_8_4_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U400_ADDRESS_DECODE.m3_LC_8_4_4  (
            .in0(N__6685),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6607),
            .lcout(\U400_ADDRESS_DECODE.N_4_0 ),
            .ltout(\U400_ADDRESS_DECODE.N_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m123_LC_8_4_5 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m123_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m123_LC_8_4_5 .LUT_INIT=16'b0101010101000111;
    LogicCell40 \U400_ADDRESS_DECODE.m123_LC_8_4_5  (
            .in0(N__5603),
            .in1(N__5634),
            .in2(N__5320),
            .in3(N__5541),
            .lcout(N_124_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.TA_EN_i_LC_8_5_1 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_EN_i_LC_8_5_1 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.TA_EN_i_LC_8_5_1 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \U400_SDRAM.TA_EN_i_LC_8_5_1  (
            .in0(N__6438),
            .in1(N__5305),
            .in2(_gnd_net_),
            .in3(N__5299),
            .lcout(TA_EN_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5246),
            .ce(),
            .sr(N__6741));
    defparam \U400_SDRAM.TA_OUT_LC_8_5_6 .C_ON=1'b0;
    defparam \U400_SDRAM.TA_OUT_LC_8_5_6 .SEQ_MODE=4'b1001;
    defparam \U400_SDRAM.TA_OUT_LC_8_5_6 .LUT_INIT=16'b0011001110110001;
    LogicCell40 \U400_SDRAM.TA_OUT_LC_8_5_6  (
            .in0(N__5293),
            .in1(N__5281),
            .in2(N__5265),
            .in3(N__5275),
            .lcout(TA_OUT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5246),
            .ce(),
            .sr(N__6741));
    defparam \U400_ADDRESS_DECODE.m113_LC_8_6_3 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m113_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m113_LC_8_6_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U400_ADDRESS_DECODE.m113_LC_8_6_3  (
            .in0(N__6581),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5886),
            .lcout(\U400_ADDRESS_DECODE.N_114_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_8_7_4 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.SDRAM_CONFIGURED_LC_8_7_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U400_SDRAM.SDRAM_CONFIGURED_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__5727),
            .in2(_gnd_net_),
            .in3(N__5857),
            .lcout(U400_SDRAM_SDRAM_CONFIGURED),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.SDRAM_CONFIGUREDC_net ),
            .ce(),
            .sr(N__6738));
    defparam \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_8_14_3 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_8_14_3 .LUT_INIT=16'b1111011011110111;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_8_14_3  (
            .in0(N__6026),
            .in1(N__6390),
            .in2(N__6754),
            .in3(N__6291),
            .lcout(\U400_SDRAM.un1_MA20_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_8_14_5 .C_ON=1'b0;
    defparam \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_8_14_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_8_14_5  (
            .in0(N__6025),
            .in1(N__6389),
            .in2(_gnd_net_),
            .in3(N__6290),
            .lcout(\U400_SDRAM.MA19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m128_LC_9_4_0 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m128_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m128_LC_9_4_0 .LUT_INIT=16'b0101010100001111;
    LogicCell40 \U400_ADDRESS_DECODE.m128_LC_9_4_0  (
            .in0(N__5434),
            .in1(_gnd_net_),
            .in2(N__5605),
            .in3(N__5650),
            .lcout(N_129_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m126_LC_9_4_1 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m126_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m126_LC_9_4_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \U400_ADDRESS_DECODE.m126_LC_9_4_1  (
            .in0(N__5648),
            .in1(N__5433),
            .in2(_gnd_net_),
            .in3(N__5596),
            .lcout(N_127_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m127_LC_9_4_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m127_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m127_LC_9_4_4 .LUT_INIT=16'b0000101101001111;
    LogicCell40 \U400_ADDRESS_DECODE.m127_LC_9_4_4  (
            .in0(N__5534),
            .in1(N__5649),
            .in2(N__5604),
            .in3(N__5489),
            .lcout(N_128_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m121_LC_9_5_4 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m121_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m121_LC_9_5_4 .LUT_INIT=16'b1000000001000000;
    LogicCell40 \U400_ADDRESS_DECODE.m121_LC_9_5_4  (
            .in0(N__5461),
            .in1(N__6556),
            .in2(N__6691),
            .in3(N__5576),
            .lcout(\U400_ADDRESS_DECODE.N_122_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_ADDRESS_DECODE.m125_LC_9_5_7 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.m125_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.m125_LC_9_5_7 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \U400_ADDRESS_DECODE.m125_LC_9_5_7  (
            .in0(N__5577),
            .in1(N__5542),
            .in2(N__5497),
            .in3(N__5462),
            .lcout(\U400_ADDRESS_DECODE.N_186_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_RNO_0_5_LC_9_14_5 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_RNO_0_5_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.MA_nesr_RNO_0_5_LC_9_14_5 .LUT_INIT=16'b0011001111111010;
    LogicCell40 \U400_SDRAM.MA_nesr_RNO_0_5_LC_9_14_5  (
            .in0(N__6305),
            .in1(N__6418),
            .in2(N__6409),
            .in3(N__6032),
            .lcout(\U400_SDRAM.MA_5_iv_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_RNO_0_1_LC_9_14_6 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_RNO_0_1_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \U400_SDRAM.MA_nesr_RNO_0_1_LC_9_14_6 .LUT_INIT=16'b0101111101001110;
    LogicCell40 \U400_SDRAM.MA_nesr_RNO_0_1_LC_9_14_6  (
            .in0(N__6031),
            .in1(N__6403),
            .in2(N__6322),
            .in3(N__6304),
            .lcout(\U400_SDRAM.MA_5_iv_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U400_SDRAM.MA_nesr_1_LC_9_15_2 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_1_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_1_LC_9_15_2 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \U400_SDRAM.MA_nesr_1_LC_9_15_2  (
            .in0(N__6223),
            .in1(N__6214),
            .in2(_gnd_net_),
            .in3(N__6833),
            .lcout(MA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_1C_net ),
            .ce(N__6777),
            .sr(N__6746));
    defparam \U400_SDRAM.MA_nesr_5_LC_9_15_3 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_5_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_5_LC_9_15_3 .LUT_INIT=16'b1000100011111111;
    LogicCell40 \U400_SDRAM.MA_nesr_5_LC_9_15_3  (
            .in0(N__6834),
            .in1(N__6199),
            .in2(_gnd_net_),
            .in3(N__6190),
            .lcout(MA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_1C_net ),
            .ce(N__6777),
            .sr(N__6746));
    defparam \U400_SDRAM.MA_nesr_3_LC_9_15_7 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_3_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_3_LC_9_15_7 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \U400_SDRAM.MA_nesr_3_LC_9_15_7  (
            .in0(N__6835),
            .in1(N__6166),
            .in2(N__6154),
            .in3(N__6035),
            .lcout(MA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_1C_net ),
            .ce(N__6777),
            .sr(N__6746));
    defparam \U400_SDRAM.MA_nesr_2_LC_9_16_0 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_2_LC_9_16_0 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_2_LC_9_16_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_2_LC_9_16_0  (
            .in0(N__6121),
            .in1(N__6034),
            .in2(N__6106),
            .in3(N__6850),
            .lcout(MA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_2C_net ),
            .ce(N__6800),
            .sr(N__6747));
    defparam \U400_SDRAM.MA_nesr_4_LC_9_16_1 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_4_LC_9_16_1 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_4_LC_9_16_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \U400_SDRAM.MA_nesr_4_LC_9_16_1  (
            .in0(N__6851),
            .in1(N__6091),
            .in2(N__6079),
            .in3(N__6036),
            .lcout(MA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_2C_net ),
            .ce(N__6800),
            .sr(N__6747));
    defparam \U400_SDRAM.MA_nesr_0_LC_9_16_2 .C_ON=1'b0;
    defparam \U400_SDRAM.MA_nesr_0_LC_9_16_2 .SEQ_MODE=4'b1000;
    defparam \U400_SDRAM.MA_nesr_0_LC_9_16_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U400_SDRAM.MA_nesr_0_LC_9_16_2  (
            .in0(N__6049),
            .in1(N__6033),
            .in2(N__6874),
            .in3(N__6849),
            .lcout(MA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU400_SDRAM.MA_nesr_2C_net ),
            .ce(N__6800),
            .sr(N__6747));
    defparam \U400_ADDRESS_DECODE.N_4_0_i_LC_11_6_2 .C_ON=1'b0;
    defparam \U400_ADDRESS_DECODE.N_4_0_i_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \U400_ADDRESS_DECODE.N_4_0_i_LC_11_6_2 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U400_ADDRESS_DECODE.N_4_0_i_LC_11_6_2  (
            .in0(N__6686),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6519),
            .lcout(N_4_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TAn_obuft_RNO_LC_11_6_3.C_ON=1'b0;
    defparam TAn_obuft_RNO_LC_11_6_3.SEQ_MODE=4'b0000;
    defparam TAn_obuft_RNO_LC_11_6_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 TAn_obuft_RNO_LC_11_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6445),
            .lcout(N_304_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U400_TOP

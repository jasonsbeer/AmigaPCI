// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 7 2025 17:55:14

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    DRA,
    SIZ,
    CMA,
    A,
    TSn,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    VBENn,
    CUMBEn,
    CLKRAM,
    C3,
    ASn,
    LDSn,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    DBRn,
    CLK40C,
    CLK40_IN,
    REGSPACEn,
    RAMENn,
    RASn,
    TACKn,
    C1);

    input [8:0] DRA;
    input [1:0] SIZ;
    output [10:0] CMA;
    input [20:0] A;
    input TSn;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    input C3;
    output ASn;
    output LDSn;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    input DBRn;
    output CLK40C;
    input CLK40_IN;
    input REGSPACEn;
    output RAMENn;
    output RASn;
    output TACKn;
    input C1;

    wire N__10415;
    wire N__10414;
    wire N__10413;
    wire N__10406;
    wire N__10405;
    wire N__10404;
    wire N__10397;
    wire N__10396;
    wire N__10395;
    wire N__10388;
    wire N__10387;
    wire N__10386;
    wire N__10379;
    wire N__10378;
    wire N__10377;
    wire N__10370;
    wire N__10369;
    wire N__10368;
    wire N__10361;
    wire N__10360;
    wire N__10359;
    wire N__10352;
    wire N__10351;
    wire N__10350;
    wire N__10343;
    wire N__10342;
    wire N__10341;
    wire N__10334;
    wire N__10333;
    wire N__10332;
    wire N__10325;
    wire N__10324;
    wire N__10323;
    wire N__10316;
    wire N__10315;
    wire N__10314;
    wire N__10307;
    wire N__10306;
    wire N__10305;
    wire N__10298;
    wire N__10297;
    wire N__10296;
    wire N__10289;
    wire N__10288;
    wire N__10287;
    wire N__10280;
    wire N__10279;
    wire N__10278;
    wire N__10271;
    wire N__10270;
    wire N__10269;
    wire N__10262;
    wire N__10261;
    wire N__10260;
    wire N__10253;
    wire N__10252;
    wire N__10251;
    wire N__10244;
    wire N__10243;
    wire N__10242;
    wire N__10235;
    wire N__10234;
    wire N__10233;
    wire N__10226;
    wire N__10225;
    wire N__10224;
    wire N__10217;
    wire N__10216;
    wire N__10215;
    wire N__10208;
    wire N__10207;
    wire N__10206;
    wire N__10199;
    wire N__10198;
    wire N__10197;
    wire N__10190;
    wire N__10189;
    wire N__10188;
    wire N__10181;
    wire N__10180;
    wire N__10179;
    wire N__10172;
    wire N__10171;
    wire N__10170;
    wire N__10163;
    wire N__10162;
    wire N__10161;
    wire N__10154;
    wire N__10153;
    wire N__10152;
    wire N__10145;
    wire N__10144;
    wire N__10143;
    wire N__10136;
    wire N__10135;
    wire N__10134;
    wire N__10127;
    wire N__10126;
    wire N__10125;
    wire N__10118;
    wire N__10117;
    wire N__10116;
    wire N__10109;
    wire N__10108;
    wire N__10107;
    wire N__10100;
    wire N__10099;
    wire N__10098;
    wire N__10091;
    wire N__10090;
    wire N__10089;
    wire N__10082;
    wire N__10081;
    wire N__10080;
    wire N__10073;
    wire N__10072;
    wire N__10071;
    wire N__10064;
    wire N__10063;
    wire N__10062;
    wire N__10055;
    wire N__10054;
    wire N__10053;
    wire N__10046;
    wire N__10045;
    wire N__10044;
    wire N__10037;
    wire N__10036;
    wire N__10035;
    wire N__10028;
    wire N__10027;
    wire N__10026;
    wire N__10019;
    wire N__10018;
    wire N__10017;
    wire N__10010;
    wire N__10009;
    wire N__10008;
    wire N__10001;
    wire N__10000;
    wire N__9999;
    wire N__9992;
    wire N__9991;
    wire N__9990;
    wire N__9983;
    wire N__9982;
    wire N__9981;
    wire N__9974;
    wire N__9973;
    wire N__9972;
    wire N__9965;
    wire N__9964;
    wire N__9963;
    wire N__9956;
    wire N__9955;
    wire N__9954;
    wire N__9947;
    wire N__9946;
    wire N__9945;
    wire N__9938;
    wire N__9937;
    wire N__9936;
    wire N__9929;
    wire N__9928;
    wire N__9927;
    wire N__9920;
    wire N__9919;
    wire N__9918;
    wire N__9911;
    wire N__9910;
    wire N__9909;
    wire N__9902;
    wire N__9901;
    wire N__9900;
    wire N__9893;
    wire N__9892;
    wire N__9891;
    wire N__9884;
    wire N__9883;
    wire N__9882;
    wire N__9875;
    wire N__9874;
    wire N__9873;
    wire N__9866;
    wire N__9865;
    wire N__9864;
    wire N__9857;
    wire N__9856;
    wire N__9855;
    wire N__9848;
    wire N__9847;
    wire N__9846;
    wire N__9839;
    wire N__9838;
    wire N__9837;
    wire N__9830;
    wire N__9829;
    wire N__9828;
    wire N__9821;
    wire N__9820;
    wire N__9819;
    wire N__9812;
    wire N__9811;
    wire N__9810;
    wire N__9803;
    wire N__9802;
    wire N__9801;
    wire N__9794;
    wire N__9793;
    wire N__9792;
    wire N__9785;
    wire N__9784;
    wire N__9783;
    wire N__9776;
    wire N__9775;
    wire N__9774;
    wire N__9767;
    wire N__9766;
    wire N__9765;
    wire N__9758;
    wire N__9757;
    wire N__9756;
    wire N__9749;
    wire N__9748;
    wire N__9747;
    wire N__9740;
    wire N__9739;
    wire N__9738;
    wire N__9731;
    wire N__9730;
    wire N__9729;
    wire N__9722;
    wire N__9721;
    wire N__9720;
    wire N__9713;
    wire N__9712;
    wire N__9711;
    wire N__9694;
    wire N__9693;
    wire N__9692;
    wire N__9691;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9679;
    wire N__9678;
    wire N__9675;
    wire N__9672;
    wire N__9669;
    wire N__9668;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9642;
    wire N__9631;
    wire N__9630;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9601;
    wire N__9598;
    wire N__9595;
    wire N__9592;
    wire N__9589;
    wire N__9588;
    wire N__9587;
    wire N__9586;
    wire N__9585;
    wire N__9582;
    wire N__9579;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9544;
    wire N__9541;
    wire N__9536;
    wire N__9533;
    wire N__9526;
    wire N__9525;
    wire N__9524;
    wire N__9523;
    wire N__9522;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9502;
    wire N__9501;
    wire N__9500;
    wire N__9499;
    wire N__9498;
    wire N__9497;
    wire N__9496;
    wire N__9495;
    wire N__9494;
    wire N__9493;
    wire N__9492;
    wire N__9491;
    wire N__9490;
    wire N__9489;
    wire N__9488;
    wire N__9487;
    wire N__9486;
    wire N__9485;
    wire N__9484;
    wire N__9483;
    wire N__9482;
    wire N__9479;
    wire N__9478;
    wire N__9477;
    wire N__9476;
    wire N__9475;
    wire N__9474;
    wire N__9473;
    wire N__9472;
    wire N__9471;
    wire N__9470;
    wire N__9469;
    wire N__9468;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9460;
    wire N__9457;
    wire N__9454;
    wire N__9453;
    wire N__9452;
    wire N__9451;
    wire N__9450;
    wire N__9449;
    wire N__9448;
    wire N__9447;
    wire N__9446;
    wire N__9445;
    wire N__9442;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9319;
    wire N__9316;
    wire N__9313;
    wire N__9310;
    wire N__9309;
    wire N__9308;
    wire N__9307;
    wire N__9306;
    wire N__9305;
    wire N__9304;
    wire N__9303;
    wire N__9300;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9276;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9234;
    wire N__9231;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9138;
    wire N__9135;
    wire N__9132;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9114;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9100;
    wire N__9097;
    wire N__9096;
    wire N__9095;
    wire N__9094;
    wire N__9093;
    wire N__9092;
    wire N__9091;
    wire N__9090;
    wire N__9087;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9063;
    wire N__9062;
    wire N__9059;
    wire N__9054;
    wire N__9049;
    wire N__9048;
    wire N__9045;
    wire N__9042;
    wire N__9039;
    wire N__9034;
    wire N__9033;
    wire N__9030;
    wire N__9027;
    wire N__9026;
    wire N__9025;
    wire N__9022;
    wire N__9021;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9003;
    wire N__8996;
    wire N__8989;
    wire N__8986;
    wire N__8983;
    wire N__8980;
    wire N__8977;
    wire N__8974;
    wire N__8971;
    wire N__8968;
    wire N__8965;
    wire N__8962;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8949;
    wire N__8946;
    wire N__8943;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8912;
    wire N__8911;
    wire N__8910;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8890;
    wire N__8889;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8877;
    wire N__8872;
    wire N__8867;
    wire N__8864;
    wire N__8851;
    wire N__8850;
    wire N__8849;
    wire N__8846;
    wire N__8845;
    wire N__8844;
    wire N__8841;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8826;
    wire N__8821;
    wire N__8818;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8784;
    wire N__8783;
    wire N__8782;
    wire N__8781;
    wire N__8780;
    wire N__8779;
    wire N__8778;
    wire N__8777;
    wire N__8776;
    wire N__8775;
    wire N__8774;
    wire N__8773;
    wire N__8772;
    wire N__8771;
    wire N__8770;
    wire N__8769;
    wire N__8768;
    wire N__8767;
    wire N__8766;
    wire N__8765;
    wire N__8764;
    wire N__8763;
    wire N__8762;
    wire N__8761;
    wire N__8760;
    wire N__8759;
    wire N__8758;
    wire N__8755;
    wire N__8754;
    wire N__8753;
    wire N__8752;
    wire N__8751;
    wire N__8750;
    wire N__8749;
    wire N__8748;
    wire N__8747;
    wire N__8674;
    wire N__8671;
    wire N__8670;
    wire N__8669;
    wire N__8668;
    wire N__8665;
    wire N__8664;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8620;
    wire N__8617;
    wire N__8608;
    wire N__8605;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8587;
    wire N__8584;
    wire N__8581;
    wire N__8578;
    wire N__8575;
    wire N__8572;
    wire N__8571;
    wire N__8570;
    wire N__8569;
    wire N__8566;
    wire N__8565;
    wire N__8564;
    wire N__8563;
    wire N__8562;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8554;
    wire N__8553;
    wire N__8552;
    wire N__8549;
    wire N__8548;
    wire N__8547;
    wire N__8546;
    wire N__8545;
    wire N__8542;
    wire N__8539;
    wire N__8536;
    wire N__8529;
    wire N__8528;
    wire N__8527;
    wire N__8526;
    wire N__8525;
    wire N__8524;
    wire N__8523;
    wire N__8516;
    wire N__8511;
    wire N__8508;
    wire N__8505;
    wire N__8500;
    wire N__8499;
    wire N__8496;
    wire N__8487;
    wire N__8484;
    wire N__8473;
    wire N__8468;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8452;
    wire N__8447;
    wire N__8438;
    wire N__8431;
    wire N__8430;
    wire N__8429;
    wire N__8424;
    wire N__8423;
    wire N__8422;
    wire N__8421;
    wire N__8420;
    wire N__8419;
    wire N__8418;
    wire N__8417;
    wire N__8416;
    wire N__8415;
    wire N__8412;
    wire N__8409;
    wire N__8406;
    wire N__8403;
    wire N__8402;
    wire N__8401;
    wire N__8400;
    wire N__8397;
    wire N__8396;
    wire N__8395;
    wire N__8394;
    wire N__8391;
    wire N__8390;
    wire N__8389;
    wire N__8388;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8371;
    wire N__8366;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8346;
    wire N__8343;
    wire N__8336;
    wire N__8331;
    wire N__8330;
    wire N__8327;
    wire N__8318;
    wire N__8311;
    wire N__8304;
    wire N__8301;
    wire N__8296;
    wire N__8293;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8259;
    wire N__8256;
    wire N__8253;
    wire N__8250;
    wire N__8245;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8233;
    wire N__8230;
    wire N__8227;
    wire N__8226;
    wire N__8223;
    wire N__8220;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8185;
    wire N__8182;
    wire N__8179;
    wire N__8178;
    wire N__8175;
    wire N__8172;
    wire N__8167;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8155;
    wire N__8154;
    wire N__8149;
    wire N__8146;
    wire N__8143;
    wire N__8140;
    wire N__8137;
    wire N__8136;
    wire N__8135;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8122;
    wire N__8117;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8103;
    wire N__8100;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8083;
    wire N__8082;
    wire N__8077;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8064;
    wire N__8063;
    wire N__8062;
    wire N__8059;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8043;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8031;
    wire N__8030;
    wire N__8029;
    wire N__8026;
    wire N__8019;
    wire N__8014;
    wire N__8011;
    wire N__8008;
    wire N__8005;
    wire N__8002;
    wire N__7999;
    wire N__7998;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7981;
    wire N__7980;
    wire N__7979;
    wire N__7978;
    wire N__7977;
    wire N__7974;
    wire N__7971;
    wire N__7966;
    wire N__7965;
    wire N__7962;
    wire N__7961;
    wire N__7960;
    wire N__7959;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7938;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7920;
    wire N__7915;
    wire N__7912;
    wire N__7897;
    wire N__7896;
    wire N__7893;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7885;
    wire N__7884;
    wire N__7883;
    wire N__7880;
    wire N__7875;
    wire N__7872;
    wire N__7867;
    wire N__7858;
    wire N__7855;
    wire N__7852;
    wire N__7849;
    wire N__7846;
    wire N__7845;
    wire N__7844;
    wire N__7843;
    wire N__7842;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7825;
    wire N__7824;
    wire N__7823;
    wire N__7822;
    wire N__7821;
    wire N__7812;
    wire N__7809;
    wire N__7806;
    wire N__7803;
    wire N__7800;
    wire N__7797;
    wire N__7788;
    wire N__7785;
    wire N__7782;
    wire N__7779;
    wire N__7776;
    wire N__7771;
    wire N__7768;
    wire N__7765;
    wire N__7762;
    wire N__7759;
    wire N__7756;
    wire N__7753;
    wire N__7750;
    wire N__7747;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7739;
    wire N__7734;
    wire N__7733;
    wire N__7732;
    wire N__7729;
    wire N__7728;
    wire N__7725;
    wire N__7722;
    wire N__7719;
    wire N__7716;
    wire N__7713;
    wire N__7710;
    wire N__7705;
    wire N__7702;
    wire N__7699;
    wire N__7692;
    wire N__7687;
    wire N__7684;
    wire N__7683;
    wire N__7680;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7654;
    wire N__7651;
    wire N__7648;
    wire N__7645;
    wire N__7642;
    wire N__7639;
    wire N__7636;
    wire N__7633;
    wire N__7630;
    wire N__7627;
    wire N__7624;
    wire N__7621;
    wire N__7618;
    wire N__7615;
    wire N__7612;
    wire N__7609;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7591;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7570;
    wire N__7567;
    wire N__7564;
    wire N__7561;
    wire N__7558;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7537;
    wire N__7536;
    wire N__7535;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7527;
    wire N__7526;
    wire N__7525;
    wire N__7524;
    wire N__7523;
    wire N__7522;
    wire N__7517;
    wire N__7516;
    wire N__7513;
    wire N__7510;
    wire N__7509;
    wire N__7506;
    wire N__7505;
    wire N__7504;
    wire N__7503;
    wire N__7500;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7479;
    wire N__7476;
    wire N__7473;
    wire N__7468;
    wire N__7465;
    wire N__7460;
    wire N__7441;
    wire N__7440;
    wire N__7437;
    wire N__7434;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7419;
    wire N__7416;
    wire N__7413;
    wire N__7408;
    wire N__7407;
    wire N__7404;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7391;
    wire N__7388;
    wire N__7381;
    wire N__7378;
    wire N__7375;
    wire N__7374;
    wire N__7373;
    wire N__7370;
    wire N__7369;
    wire N__7366;
    wire N__7363;
    wire N__7360;
    wire N__7357;
    wire N__7348;
    wire N__7345;
    wire N__7344;
    wire N__7341;
    wire N__7338;
    wire N__7337;
    wire N__7336;
    wire N__7333;
    wire N__7330;
    wire N__7325;
    wire N__7322;
    wire N__7319;
    wire N__7312;
    wire N__7311;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7291;
    wire N__7288;
    wire N__7285;
    wire N__7282;
    wire N__7279;
    wire N__7276;
    wire N__7273;
    wire N__7272;
    wire N__7271;
    wire N__7270;
    wire N__7269;
    wire N__7268;
    wire N__7267;
    wire N__7266;
    wire N__7259;
    wire N__7254;
    wire N__7247;
    wire N__7240;
    wire N__7239;
    wire N__7238;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7224;
    wire N__7221;
    wire N__7220;
    wire N__7219;
    wire N__7218;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7204;
    wire N__7195;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7182;
    wire N__7179;
    wire N__7176;
    wire N__7173;
    wire N__7170;
    wire N__7167;
    wire N__7162;
    wire N__7161;
    wire N__7158;
    wire N__7157;
    wire N__7156;
    wire N__7155;
    wire N__7152;
    wire N__7151;
    wire N__7146;
    wire N__7141;
    wire N__7140;
    wire N__7139;
    wire N__7138;
    wire N__7137;
    wire N__7136;
    wire N__7135;
    wire N__7134;
    wire N__7133;
    wire N__7132;
    wire N__7131;
    wire N__7130;
    wire N__7125;
    wire N__7122;
    wire N__7119;
    wire N__7110;
    wire N__7107;
    wire N__7104;
    wire N__7099;
    wire N__7096;
    wire N__7091;
    wire N__7086;
    wire N__7083;
    wire N__7080;
    wire N__7063;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7050;
    wire N__7049;
    wire N__7048;
    wire N__7047;
    wire N__7046;
    wire N__7045;
    wire N__7044;
    wire N__7043;
    wire N__7042;
    wire N__7041;
    wire N__7040;
    wire N__7039;
    wire N__7034;
    wire N__7031;
    wire N__7030;
    wire N__7029;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7013;
    wire N__7008;
    wire N__7007;
    wire N__7004;
    wire N__7003;
    wire N__7002;
    wire N__7001;
    wire N__7000;
    wire N__6999;
    wire N__6998;
    wire N__6995;
    wire N__6994;
    wire N__6993;
    wire N__6992;
    wire N__6991;
    wire N__6988;
    wire N__6985;
    wire N__6978;
    wire N__6975;
    wire N__6968;
    wire N__6965;
    wire N__6962;
    wire N__6959;
    wire N__6954;
    wire N__6949;
    wire N__6944;
    wire N__6941;
    wire N__6934;
    wire N__6927;
    wire N__6922;
    wire N__6901;
    wire N__6900;
    wire N__6899;
    wire N__6898;
    wire N__6897;
    wire N__6894;
    wire N__6893;
    wire N__6890;
    wire N__6889;
    wire N__6886;
    wire N__6885;
    wire N__6882;
    wire N__6881;
    wire N__6880;
    wire N__6879;
    wire N__6876;
    wire N__6873;
    wire N__6870;
    wire N__6869;
    wire N__6866;
    wire N__6861;
    wire N__6856;
    wire N__6849;
    wire N__6846;
    wire N__6845;
    wire N__6844;
    wire N__6839;
    wire N__6836;
    wire N__6829;
    wire N__6828;
    wire N__6823;
    wire N__6820;
    wire N__6817;
    wire N__6810;
    wire N__6807;
    wire N__6796;
    wire N__6793;
    wire N__6790;
    wire N__6787;
    wire N__6784;
    wire N__6781;
    wire N__6778;
    wire N__6775;
    wire N__6772;
    wire N__6769;
    wire N__6766;
    wire N__6763;
    wire N__6760;
    wire N__6757;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6745;
    wire N__6742;
    wire N__6741;
    wire N__6736;
    wire N__6733;
    wire N__6732;
    wire N__6731;
    wire N__6728;
    wire N__6723;
    wire N__6718;
    wire N__6715;
    wire N__6714;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6694;
    wire N__6691;
    wire N__6688;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6678;
    wire N__6677;
    wire N__6676;
    wire N__6675;
    wire N__6674;
    wire N__6673;
    wire N__6670;
    wire N__6667;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6630;
    wire N__6627;
    wire N__6626;
    wire N__6623;
    wire N__6622;
    wire N__6621;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6606;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6582;
    wire N__6581;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6529;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6502;
    wire N__6499;
    wire N__6496;
    wire N__6493;
    wire N__6490;
    wire N__6487;
    wire N__6484;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6349;
    wire N__6346;
    wire N__6343;
    wire N__6340;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6325;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6286;
    wire N__6283;
    wire N__6280;
    wire N__6277;
    wire N__6274;
    wire N__6271;
    wire N__6268;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6247;
    wire N__6246;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6236;
    wire N__6235;
    wire N__6230;
    wire N__6227;
    wire N__6224;
    wire N__6221;
    wire N__6216;
    wire N__6211;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6203;
    wire N__6200;
    wire N__6197;
    wire N__6196;
    wire N__6193;
    wire N__6192;
    wire N__6187;
    wire N__6186;
    wire N__6185;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6173;
    wire N__6168;
    wire N__6165;
    wire N__6162;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6129;
    wire N__6126;
    wire N__6123;
    wire N__6118;
    wire N__6117;
    wire N__6114;
    wire N__6111;
    wire N__6106;
    wire N__6103;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6093;
    wire N__6092;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6080;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6066;
    wire N__6063;
    wire N__6062;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6030;
    wire N__6027;
    wire N__6024;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6005;
    wire N__6004;
    wire N__6003;
    wire N__6002;
    wire N__6001;
    wire N__5998;
    wire N__5995;
    wire N__5992;
    wire N__5991;
    wire N__5990;
    wire N__5989;
    wire N__5980;
    wire N__5979;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5967;
    wire N__5964;
    wire N__5961;
    wire N__5958;
    wire N__5955;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5929;
    wire N__5926;
    wire N__5925;
    wire N__5920;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5910;
    wire N__5907;
    wire N__5904;
    wire N__5901;
    wire N__5898;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5881;
    wire N__5878;
    wire N__5875;
    wire N__5874;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5857;
    wire N__5856;
    wire N__5853;
    wire N__5850;
    wire N__5845;
    wire N__5842;
    wire N__5839;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5815;
    wire N__5812;
    wire N__5809;
    wire N__5806;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5788;
    wire N__5785;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5739;
    wire N__5736;
    wire N__5733;
    wire N__5728;
    wire N__5725;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5704;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5692;
    wire N__5689;
    wire N__5686;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5665;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5644;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5575;
    wire N__5574;
    wire N__5571;
    wire N__5568;
    wire N__5565;
    wire N__5560;
    wire N__5557;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5545;
    wire N__5542;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5487;
    wire N__5484;
    wire N__5481;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5445;
    wire N__5444;
    wire N__5443;
    wire N__5438;
    wire N__5433;
    wire N__5428;
    wire N__5427;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5401;
    wire N__5398;
    wire N__5397;
    wire N__5394;
    wire N__5391;
    wire N__5386;
    wire N__5383;
    wire N__5382;
    wire N__5379;
    wire N__5376;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5314;
    wire N__5311;
    wire N__5310;
    wire N__5309;
    wire N__5304;
    wire N__5301;
    wire N__5296;
    wire N__5293;
    wire N__5292;
    wire N__5291;
    wire N__5286;
    wire N__5283;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5268;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5230;
    wire N__5227;
    wire N__5224;
    wire N__5221;
    wire N__5218;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5187;
    wire N__5182;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5167;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5154;
    wire N__5149;
    wire N__5146;
    wire N__5145;
    wire N__5142;
    wire N__5139;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5115;
    wire N__5110;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5074;
    wire N__5073;
    wire N__5068;
    wire N__5065;
    wire N__5062;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5047;
    wire N__5046;
    wire N__5043;
    wire N__5040;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5023;
    wire N__5020;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5010;
    wire N__5007;
    wire N__5002;
    wire N__4999;
    wire N__4996;
    wire N__4993;
    wire N__4990;
    wire N__4987;
    wire N__4986;
    wire N__4985;
    wire N__4980;
    wire N__4977;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4969;
    wire N__4966;
    wire N__4963;
    wire N__4960;
    wire N__4957;
    wire N__4954;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4927;
    wire N__4924;
    wire N__4921;
    wire N__4918;
    wire N__4915;
    wire N__4912;
    wire N__4909;
    wire N__4906;
    wire N__4905;
    wire N__4902;
    wire N__4899;
    wire N__4894;
    wire N__4893;
    wire N__4890;
    wire N__4887;
    wire N__4882;
    wire N__4881;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4867;
    wire N__4864;
    wire N__4861;
    wire N__4858;
    wire N__4857;
    wire N__4856;
    wire N__4855;
    wire N__4854;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4831;
    wire N__4830;
    wire N__4825;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4809;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4780;
    wire N__4777;
    wire N__4776;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4759;
    wire N__4758;
    wire N__4757;
    wire N__4756;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4744;
    wire N__4735;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4725;
    wire N__4720;
    wire N__4717;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4702;
    wire N__4699;
    wire N__4696;
    wire N__4693;
    wire N__4692;
    wire N__4689;
    wire N__4688;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4672;
    wire N__4669;
    wire N__4666;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4651;
    wire N__4648;
    wire N__4645;
    wire N__4644;
    wire N__4641;
    wire N__4638;
    wire N__4633;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4573;
    wire N__4570;
    wire N__4567;
    wire N__4564;
    wire N__4561;
    wire N__4560;
    wire N__4557;
    wire N__4556;
    wire N__4555;
    wire N__4552;
    wire N__4549;
    wire N__4546;
    wire N__4543;
    wire N__4540;
    wire N__4531;
    wire N__4530;
    wire N__4527;
    wire N__4524;
    wire N__4519;
    wire N__4516;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4501;
    wire N__4500;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4482;
    wire N__4471;
    wire N__4468;
    wire N__4467;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4441;
    wire N__4440;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4405;
    wire N__4404;
    wire N__4403;
    wire N__4400;
    wire N__4399;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4378;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4368;
    wire N__4363;
    wire N__4360;
    wire N__4357;
    wire N__4354;
    wire N__4351;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4338;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4300;
    wire N__4299;
    wire N__4296;
    wire N__4293;
    wire N__4288;
    wire N__4287;
    wire N__4286;
    wire N__4281;
    wire N__4278;
    wire N__4273;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4261;
    wire N__4258;
    wire N__4257;
    wire N__4256;
    wire N__4255;
    wire N__4254;
    wire N__4253;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4241;
    wire N__4238;
    wire N__4231;
    wire N__4222;
    wire N__4219;
    wire N__4216;
    wire N__4213;
    wire N__4210;
    wire N__4209;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4192;
    wire N__4191;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4174;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4144;
    wire N__4143;
    wire N__4142;
    wire N__4135;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4127;
    wire N__4126;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4110;
    wire N__4107;
    wire N__4104;
    wire N__4099;
    wire N__4096;
    wire N__4095;
    wire N__4094;
    wire N__4093;
    wire N__4086;
    wire N__4083;
    wire N__4078;
    wire N__4075;
    wire N__4072;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4055;
    wire N__4052;
    wire N__4047;
    wire N__4042;
    wire N__4039;
    wire N__4036;
    wire N__4033;
    wire N__4030;
    wire N__4027;
    wire N__4024;
    wire N__4023;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4006;
    wire N__4003;
    wire N__4000;
    wire N__3997;
    wire N__3996;
    wire N__3995;
    wire N__3994;
    wire N__3985;
    wire N__3982;
    wire N__3979;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3963;
    wire N__3960;
    wire N__3957;
    wire N__3954;
    wire N__3949;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3937;
    wire N__3934;
    wire N__3931;
    wire N__3928;
    wire N__3925;
    wire N__3922;
    wire N__3919;
    wire N__3916;
    wire N__3913;
    wire N__3910;
    wire N__3907;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3889;
    wire N__3886;
    wire N__3883;
    wire N__3880;
    wire N__3877;
    wire N__3874;
    wire N__3871;
    wire N__3868;
    wire N__3865;
    wire N__3862;
    wire N__3859;
    wire N__3856;
    wire N__3853;
    wire N__3850;
    wire N__3847;
    wire N__3844;
    wire N__3841;
    wire N__3838;
    wire N__3835;
    wire N__3832;
    wire N__3829;
    wire N__3826;
    wire N__3825;
    wire N__3822;
    wire N__3819;
    wire N__3814;
    wire N__3811;
    wire N__3808;
    wire N__3805;
    wire N__3804;
    wire N__3801;
    wire N__3798;
    wire N__3795;
    wire N__3792;
    wire N__3787;
    wire N__3784;
    wire N__3781;
    wire N__3778;
    wire N__3775;
    wire N__3774;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3760;
    wire N__3759;
    wire N__3758;
    wire N__3757;
    wire N__3750;
    wire N__3747;
    wire N__3744;
    wire N__3739;
    wire N__3736;
    wire N__3733;
    wire N__3730;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3715;
    wire N__3712;
    wire N__3709;
    wire N__3706;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3694;
    wire N__3691;
    wire N__3688;
    wire N__3685;
    wire N__3682;
    wire N__3679;
    wire N__3676;
    wire N__3673;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_OUT_i_i;
    wire CLK40_OUT_i_i;
    wire REGSPACEn_c;
    wire \U712_REG_SM.REG_CYCLE_GOZ0 ;
    wire \U712_REG_SM.UDS_OUT_2_0_a2_0_a3_0 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.LDS_OUT_2_0_a2_0_a3_0 ;
    wire \U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1 ;
    wire N_944_i;
    wire VBENn_c;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_cascade_ ;
    wire N_41_i;
    wire \U712_BYTE_ENABLE.N_273 ;
    wire N_43_i;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0 ;
    wire \U712_BYTE_ENABLE.N_275_cascade_ ;
    wire N_42_i;
    wire \U712_BYTE_ENABLE.N_271_cascade_ ;
    wire N_44_i;
    wire A_c_0;
    wire A_c_1;
    wire \U712_BYTE_ENABLE.N_277 ;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire \U712_BYTE_ENABLE.N_270 ;
    wire ASn_c;
    wire \U712_REG_SM.N_266_cascade_ ;
    wire \U712_REG_SM.N_215 ;
    wire \U712_REG_SM.N_215_cascade_ ;
    wire \U712_REG_SM.N_200_cascade_ ;
    wire \U712_REG_SM.C1_SYNCZ0Z_2 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_6 ;
    wire \U712_REG_SM.N_200 ;
    wire \U712_REG_SM.N_219 ;
    wire \U712_REG_SM.N_325_cascade_ ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_198 ;
    wire \U712_REG_SM.N_212 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_REG_SM.N_198_cascade_ ;
    wire \U712_REG_SM.DS_EN_RNOZ0Z_0_cascade_ ;
    wire C3_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.LDS_OUTZ0 ;
    wire U712_REG_SM_un1_LDSn_i;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0 ;
    wire bfn_9_9_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire TSn_c;
    wire RAMSPACEn_c;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.N_325 ;
    wire \U712_REG_SM.N_201 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_RNOZ0Z_0 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.N_265 ;
    wire \U712_REG_SM.N_183 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_2 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire U712_REG_SM_DBR_SYNC_1;
    wire \U712_CHIP_RAM.DBR_SYNCZ0Z_2 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_177_cascade_ ;
    wire \U712_CHIP_RAM.N_197 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ;
    wire \U712_CHIP_RAM.N_307_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_cascade_ ;
    wire CASUn_c;
    wire CASLn_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire U712_REG_SM_DBR_SYNC_0;
    wire \U712_REG_SM.DS_ENZ0 ;
    wire \U712_REG_SM.UDS_OUTZ0 ;
    wire U712_REG_SM_un1_UDSn_i;
    wire RnW_c;
    wire DRDDIR_i_m4_i_m2;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire \U712_CHIP_RAM.REFRESH5lto2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH5lto1 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire A_c_4;
    wire A_c_11;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.N_209 ;
    wire AWEn_c;
    wire DBDIR_c;
    wire \U712_CHIP_RAM.N_323_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a2_0_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a3_3_2_0_cascade_ ;
    wire \U712_CHIP_RAM.N_242_cascade_ ;
    wire \U712_CHIP_RAM.N_188_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0_0 ;
    wire \U712_CHIP_RAM.N_306 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0 ;
    wire \U712_CHIP_RAM.N_238 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_323 ;
    wire \U712_CHIP_RAM.N_240 ;
    wire \U712_CHIP_RAM.N_10_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER16_cascade_ ;
    wire \U712_CHIP_RAM.N_328 ;
    wire \U712_CHIP_RAM.N_307 ;
    wire \U712_CHIP_RAM.N_328_cascade_ ;
    wire \U712_CHIP_RAM.N_177 ;
    wire \U712_CHIP_RAM.N_251_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_cascade_ ;
    wire bfn_10_14_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire TACK_EN_i_ess;
    wire A_c_18;
    wire A_c_16;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CMA_c_2;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.un1_CMA30_0_i_cascade_ ;
    wire A_c_5;
    wire A_c_12;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire A_c_3;
    wire A_c_10;
    wire A_c_9;
    wire A_c_2;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_2_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_66_0_i_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNI9MVM2Z0Z_1 ;
    wire \U712_CHIP_RAM.N_222 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_9_0_cascade_ ;
    wire DBENn_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_3_0 ;
    wire \U712_CHIP_RAM.N_305_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_2_cascade_ ;
    wire \U712_CHIP_RAM.N_221 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ;
    wire \U712_CHIP_RAM.N_305 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_cascade_ ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.N_10 ;
    wire \U712_CHIP_RAM.N_260 ;
    wire \U712_CYCLE_TERM.N_214_i_0_en_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_3 ;
    wire CONSTANT_ONE_NET;
    wire CRCSn_c;
    wire WEn_c;
    wire A_c_19;
    wire RAS0n_c;
    wire CMA_c_9;
    wire A_c_17;
    wire CMA_c_8;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire A_c_15;
    wire A_c_8;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire CMA_c_1;
    wire CMA_c_5;
    wire A_c_7;
    wire \U712_CHIP_RAM.N_316_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire A_c_14;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_3_0_0 ;
    wire \U712_CHIP_RAM.N_180 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a3_2_1_0 ;
    wire \U712_CHIP_RAM.N_254_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1Z0Z_1 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_0 ;
    wire CPU_TACKm;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.N_187 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_5 ;
    wire REG_TACK;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_0_a3_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a3_0_a3_0 ;
    wire \U712_CHIP_RAM.N_96 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER16 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_0_a3_0 ;
    wire \U712_CYCLE_TERM.N_214_i_0_en ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.N_312 ;
    wire \U712_CHIP_RAM.N_243 ;
    wire RESETn_c;
    wire RESETn_c_i;
    wire RAMENn_c;
    wire REG_CYCLEm;
    wire DRDENn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire CLK40_OUT_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire TACK_OUTn;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire CASn_c;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ;
    wire CMA_c_4;
    wire CLK80_OUT;
    wire \U712_CHIP_RAM.un1_CMA30_0_i_0 ;
    wire A_c_13;
    wire A_c_6;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CPU_CYCLEm;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire C1_c_g;
    wire DBRn_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_8C_net ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire C3_c_g;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire _gnd_net_;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ;
    wire RESETn_c_i_g;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_OUT_i),
            .REFERENCECLK(N__3691),
            .RESETB(N__6424),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_OUT),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__10415),
            .DIN(N__10414),
            .DOUT(N__10413),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__10415),
            .PADOUT(N__10414),
            .PADIN(N__10413),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5890),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__10406),
            .DIN(N__10405),
            .DOUT(N__10404),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__10406),
            .PADOUT(N__10405),
            .PADIN(N__10404),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__10397),
            .DIN(N__10396),
            .DOUT(N__10395),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__10397),
            .PADOUT(N__10396),
            .PADIN(N__10395),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8977),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__10388),
            .DIN(N__10387),
            .DOUT(N__10386),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__10388),
            .PADOUT(N__10387),
            .PADIN(N__10386),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4927),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__10379),
            .DIN(N__10378),
            .DOUT(N__10377),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__10379),
            .PADOUT(N__10378),
            .PADIN(N__10377),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__10370),
            .DIN(N__10369),
            .DOUT(N__10368),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__10370),
            .PADOUT(N__10369),
            .PADIN(N__10368),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__10361),
            .DIN(N__10360),
            .DOUT(N__10359),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__10361),
            .PADOUT(N__10360),
            .PADIN(N__10359),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__10352),
            .DIN(N__10351),
            .DOUT(N__10350),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__10352),
            .PADOUT(N__10351),
            .PADIN(N__10350),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__10343),
            .DIN(N__10342),
            .DOUT(N__10341),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__10343),
            .PADOUT(N__10342),
            .PADIN(N__10341),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__10334),
            .DIN(N__10333),
            .DOUT(N__10332),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__10334),
            .PADOUT(N__10333),
            .PADIN(N__10332),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6553),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__10325),
            .DIN(N__10324),
            .DOUT(N__10323),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__10325),
            .PADOUT(N__10324),
            .PADIN(N__10323),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7759),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__10316),
            .DIN(N__10315),
            .DOUT(N__10314),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__10316),
            .PADOUT(N__10315),
            .PADIN(N__10314),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__10307),
            .DIN(N__10306),
            .DOUT(N__10305),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__10307),
            .PADOUT(N__10306),
            .PADIN(N__10305),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__10298),
            .DIN(N__10297),
            .DOUT(N__10296),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__10298),
            .PADOUT(N__10297),
            .PADIN(N__10296),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3907),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__10289),
            .DIN(N__10288),
            .DOUT(N__10287),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__10289),
            .PADOUT(N__10288),
            .PADIN(N__10287),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__10280),
            .DIN(N__10279),
            .DOUT(N__10278),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__10280),
            .PADOUT(N__10279),
            .PADIN(N__10278),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__10271),
            .DIN(N__10270),
            .DOUT(N__10269),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__10271),
            .PADOUT(N__10270),
            .PADIN(N__10269),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7627),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__10262),
            .DIN(N__10261),
            .DOUT(N__10260),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__10262),
            .PADOUT(N__10261),
            .PADIN(N__10260),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__10253),
            .DIN(N__10252),
            .DOUT(N__10251),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__10253),
            .PADOUT(N__10252),
            .PADIN(N__10251),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6409),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__10244),
            .DIN(N__10243),
            .DOUT(N__10242),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__10244),
            .PADOUT(N__10243),
            .PADIN(N__10242),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__10235),
            .DIN(N__10234),
            .DOUT(N__10233),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__10235),
            .PADOUT(N__10234),
            .PADIN(N__10233),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__10226),
            .DIN(N__10225),
            .DOUT(N__10224),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__10226),
            .PADOUT(N__10225),
            .PADIN(N__10224),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__10217),
            .DIN(N__10216),
            .DOUT(N__10215),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__10217),
            .PADOUT(N__10216),
            .PADIN(N__10215),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__10208),
            .DIN(N__10207),
            .DOUT(N__10206),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__10208),
            .PADOUT(N__10207),
            .PADIN(N__10206),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__10199),
            .DIN(N__10198),
            .DOUT(N__10197),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__10199),
            .PADOUT(N__10198),
            .PADIN(N__10197),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__10190),
            .DIN(N__10189),
            .DOUT(N__10188),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__10190),
            .PADOUT(N__10189),
            .PADIN(N__10188),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__10181),
            .DIN(N__10180),
            .DOUT(N__10179),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__10181),
            .PADOUT(N__10180),
            .PADIN(N__10179),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__10172),
            .DIN(N__10171),
            .DOUT(N__10170),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__10172),
            .PADOUT(N__10171),
            .PADIN(N__10170),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__10163),
            .DIN(N__10162),
            .DOUT(N__10161),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__10163),
            .PADOUT(N__10162),
            .PADIN(N__10161),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6271),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__10154),
            .DIN(N__10153),
            .DOUT(N__10152),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__10154),
            .PADOUT(N__10153),
            .PADIN(N__10152),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__10145),
            .DIN(N__10144),
            .DOUT(N__10143),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__10145),
            .PADOUT(N__10144),
            .PADIN(N__10143),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__10136),
            .DIN(N__10135),
            .DOUT(N__10134),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__10136),
            .PADOUT(N__10135),
            .PADIN(N__10134),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__10127),
            .DIN(N__10126),
            .DOUT(N__10125),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__10127),
            .PADOUT(N__10126),
            .PADIN(N__10125),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__10118),
            .DIN(N__10117),
            .DOUT(N__10116),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__10118),
            .PADOUT(N__10117),
            .PADIN(N__10116),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3724),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__10109),
            .DIN(N__10108),
            .DOUT(N__10107),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__10109),
            .PADOUT(N__10108),
            .PADIN(N__10107),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4363),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__10100),
            .DIN(N__10099),
            .DOUT(N__10098),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__10100),
            .PADOUT(N__10099),
            .PADIN(N__10098),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__10091),
            .DIN(N__10090),
            .DOUT(N__10089),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__10091),
            .PADOUT(N__10090),
            .PADIN(N__10089),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8989),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__10082),
            .DIN(N__10081),
            .DOUT(N__10080),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__10082),
            .PADOUT(N__10081),
            .PADIN(N__10080),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__10073),
            .DIN(N__10072),
            .DOUT(N__10071),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__10073),
            .PADOUT(N__10072),
            .PADIN(N__10071),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__10064),
            .DIN(N__10063),
            .DOUT(N__10062),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__10064),
            .PADOUT(N__10063),
            .PADIN(N__10062),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3739),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__10055),
            .DIN(N__10054),
            .DOUT(N__10053),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__10055),
            .PADOUT(N__10054),
            .PADIN(N__10053),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__10046),
            .DIN(N__10045),
            .DOUT(N__10044),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__10046),
            .PADOUT(N__10045),
            .PADIN(N__10044),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3982),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__10037),
            .DIN(N__10036),
            .DOUT(N__10035),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__10037),
            .PADOUT(N__10036),
            .PADIN(N__10035),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5647),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__10028),
            .DIN(N__10027),
            .DOUT(N__10026),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__10028),
            .PADOUT(N__10027),
            .PADIN(N__10026),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__10019),
            .DIN(N__10018),
            .DOUT(N__10017),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__10019),
            .PADOUT(N__10018),
            .PADIN(N__10017),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_0_iopad (
            .OE(N__10010),
            .DIN(N__10009),
            .DOUT(N__10008),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__10010),
            .PADOUT(N__10009),
            .PADIN(N__10008),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__10001),
            .DIN(N__10000),
            .DOUT(N__9999),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__10001),
            .PADOUT(N__10000),
            .PADIN(N__9999),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6151),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__9992),
            .DIN(N__9991),
            .DOUT(N__9990),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__9992),
            .PADOUT(N__9991),
            .PADIN(N__9990),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__9983),
            .DIN(N__9982),
            .DOUT(N__9981),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__9983),
            .PADOUT(N__9982),
            .PADIN(N__9981),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8809),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__9974),
            .DIN(N__9973),
            .DOUT(N__9972),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__9974),
            .PADOUT(N__9973),
            .PADIN(N__9972),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7654),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__9965),
            .DIN(N__9964),
            .DOUT(N__9963),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__9965),
            .PADOUT(N__9964),
            .PADIN(N__9963),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3892),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__9956),
            .DIN(N__9955),
            .DOUT(N__9954),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__9956),
            .PADOUT(N__9955),
            .PADIN(N__9954),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6331),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__9947),
            .DIN(N__9946),
            .DOUT(N__9945),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__9947),
            .PADOUT(N__9946),
            .PADIN(N__9945),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3978),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__9938),
            .DIN(N__9937),
            .DOUT(N__9936),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__9938),
            .PADOUT(N__9937),
            .PADIN(N__9936),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__9929),
            .DIN(N__9928),
            .DOUT(N__9927),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__9929),
            .PADOUT(N__9928),
            .PADIN(N__9927),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__9920),
            .DIN(N__9919),
            .DOUT(N__9918),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__9920),
            .PADOUT(N__9919),
            .PADIN(N__9918),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3844),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__9911),
            .DIN(N__9910),
            .DOUT(N__9909),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__9911),
            .PADOUT(N__9910),
            .PADIN(N__9909),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6388),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__9902),
            .DIN(N__9901),
            .DOUT(N__9900),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__9902),
            .PADOUT(N__9901),
            .PADIN(N__9900),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5230),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__9893),
            .DIN(N__9892),
            .DOUT(N__9891),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__9893),
            .PADOUT(N__9892),
            .PADIN(N__9891),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3871),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__9884),
            .DIN(N__9883),
            .DOUT(N__9882),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__9884),
            .PADOUT(N__9883),
            .PADIN(N__9882),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__9875),
            .DIN(N__9874),
            .DOUT(N__9873),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__9875),
            .PADOUT(N__9874),
            .PADIN(N__9873),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__9866),
            .DIN(N__9865),
            .DOUT(N__9864),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__9866),
            .PADOUT(N__9865),
            .PADIN(N__9864),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__9857),
            .DIN(N__9856),
            .DOUT(N__9855),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__9857),
            .PADOUT(N__9856),
            .PADIN(N__9855),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__9848),
            .DIN(N__9847),
            .DOUT(N__9846),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__9848),
            .PADOUT(N__9847),
            .PADIN(N__9846),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6463),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__9839),
            .DIN(N__9838),
            .DOUT(N__9837),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__9839),
            .PADOUT(N__9838),
            .PADIN(N__9837),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__9830),
            .DIN(N__9829),
            .DOUT(N__9828),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__9830),
            .PADOUT(N__9829),
            .PADIN(N__9828),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4165),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__9821),
            .DIN(N__9820),
            .DOUT(N__9819),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__9821),
            .PADOUT(N__9820),
            .PADIN(N__9819),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3928),
            .DIN0(),
            .DOUT0(N__8014),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__9812),
            .DIN(N__9811),
            .DOUT(N__9810),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__9812),
            .PADOUT(N__9811),
            .PADIN(N__9810),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5659),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__9803),
            .DIN(N__9802),
            .DOUT(N__9801),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__9803),
            .PADOUT(N__9802),
            .PADIN(N__9801),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__9794),
            .DIN(N__9793),
            .DOUT(N__9792),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__9794),
            .PADOUT(N__9793),
            .PADIN(N__9792),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__9785),
            .DIN(N__9784),
            .DOUT(N__9783),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__9785),
            .PADOUT(N__9784),
            .PADIN(N__9783),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6295),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__9776),
            .DIN(N__9775),
            .DOUT(N__9774),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__9776),
            .PADOUT(N__9775),
            .PADIN(N__9774),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__9767),
            .DIN(N__9766),
            .DOUT(N__9765),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__9767),
            .PADOUT(N__9766),
            .PADIN(N__9765),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__9758),
            .DIN(N__9757),
            .DOUT(N__9756),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__9758),
            .PADOUT(N__9757),
            .PADIN(N__9756),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__9749),
            .DIN(N__9748),
            .DOUT(N__9747),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__9749),
            .PADOUT(N__9748),
            .PADIN(N__9747),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__9740),
            .DIN(N__9739),
            .DOUT(N__9738),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__9740),
            .PADOUT(N__9739),
            .PADIN(N__9738),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6796),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__9731),
            .DIN(N__9730),
            .DOUT(N__9729),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__9731),
            .PADOUT(N__9730),
            .PADIN(N__9729),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5002),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__9722),
            .DIN(N__9721),
            .DOUT(N__9720),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__9722),
            .PADOUT(N__9721),
            .PADIN(N__9720),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6046),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__9713),
            .DIN(N__9712),
            .DOUT(N__9711),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__9713),
            .PADOUT(N__9712),
            .PADIN(N__9711),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CEMux I__2323 (
            .O(N__9694),
            .I(N__9688));
    CEMux I__2322 (
            .O(N__9693),
            .I(N__9685));
    CEMux I__2321 (
            .O(N__9692),
            .I(N__9682));
    CEMux I__2320 (
            .O(N__9691),
            .I(N__9679));
    LocalMux I__2319 (
            .O(N__9688),
            .I(N__9675));
    LocalMux I__2318 (
            .O(N__9685),
            .I(N__9672));
    LocalMux I__2317 (
            .O(N__9682),
            .I(N__9669));
    LocalMux I__2316 (
            .O(N__9679),
            .I(N__9664));
    CEMux I__2315 (
            .O(N__9678),
            .I(N__9661));
    Span4Mux_v I__2314 (
            .O(N__9675),
            .I(N__9658));
    Span4Mux_h I__2313 (
            .O(N__9672),
            .I(N__9653));
    Span4Mux_h I__2312 (
            .O(N__9669),
            .I(N__9653));
    CEMux I__2311 (
            .O(N__9668),
            .I(N__9650));
    CEMux I__2310 (
            .O(N__9667),
            .I(N__9647));
    Sp12to4 I__2309 (
            .O(N__9664),
            .I(N__9642));
    LocalMux I__2308 (
            .O(N__9661),
            .I(N__9642));
    Odrv4 I__2307 (
            .O(N__9658),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    Odrv4 I__2306 (
            .O(N__9653),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    LocalMux I__2305 (
            .O(N__9650),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    LocalMux I__2304 (
            .O(N__9647),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    Odrv12 I__2303 (
            .O(N__9642),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    InMux I__2302 (
            .O(N__9631),
            .I(N__9627));
    InMux I__2301 (
            .O(N__9630),
            .I(N__9624));
    LocalMux I__2300 (
            .O(N__9627),
            .I(N__9621));
    LocalMux I__2299 (
            .O(N__9624),
            .I(N__9618));
    Span4Mux_h I__2298 (
            .O(N__9621),
            .I(N__9615));
    Span4Mux_v I__2297 (
            .O(N__9618),
            .I(N__9612));
    Sp12to4 I__2296 (
            .O(N__9615),
            .I(N__9609));
    Span4Mux_v I__2295 (
            .O(N__9612),
            .I(N__9606));
    Span12Mux_v I__2294 (
            .O(N__9609),
            .I(N__9601));
    Sp12to4 I__2293 (
            .O(N__9606),
            .I(N__9601));
    Odrv12 I__2292 (
            .O(N__9601),
            .I(DRA_c_4));
    InMux I__2291 (
            .O(N__9598),
            .I(N__9595));
    LocalMux I__2290 (
            .O(N__9595),
            .I(N__9592));
    Odrv12 I__2289 (
            .O(N__9592),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    CEMux I__2288 (
            .O(N__9589),
            .I(N__9582));
    CEMux I__2287 (
            .O(N__9588),
            .I(N__9579));
    CEMux I__2286 (
            .O(N__9587),
            .I(N__9575));
    CEMux I__2285 (
            .O(N__9586),
            .I(N__9572));
    CEMux I__2284 (
            .O(N__9585),
            .I(N__9569));
    LocalMux I__2283 (
            .O(N__9582),
            .I(N__9566));
    LocalMux I__2282 (
            .O(N__9579),
            .I(N__9563));
    CEMux I__2281 (
            .O(N__9578),
            .I(N__9560));
    LocalMux I__2280 (
            .O(N__9575),
            .I(N__9557));
    LocalMux I__2279 (
            .O(N__9572),
            .I(N__9554));
    LocalMux I__2278 (
            .O(N__9569),
            .I(N__9551));
    Span4Mux_h I__2277 (
            .O(N__9566),
            .I(N__9544));
    Span4Mux_v I__2276 (
            .O(N__9563),
            .I(N__9544));
    LocalMux I__2275 (
            .O(N__9560),
            .I(N__9544));
    Span4Mux_h I__2274 (
            .O(N__9557),
            .I(N__9541));
    Span4Mux_v I__2273 (
            .O(N__9554),
            .I(N__9536));
    Span4Mux_h I__2272 (
            .O(N__9551),
            .I(N__9536));
    Sp12to4 I__2271 (
            .O(N__9544),
            .I(N__9533));
    Odrv4 I__2270 (
            .O(N__9541),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    Odrv4 I__2269 (
            .O(N__9536),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    Odrv12 I__2268 (
            .O(N__9533),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    InMux I__2267 (
            .O(N__9526),
            .I(N__9518));
    InMux I__2266 (
            .O(N__9525),
            .I(N__9515));
    InMux I__2265 (
            .O(N__9524),
            .I(N__9512));
    InMux I__2264 (
            .O(N__9523),
            .I(N__9509));
    InMux I__2263 (
            .O(N__9522),
            .I(N__9506));
    InMux I__2262 (
            .O(N__9521),
            .I(N__9503));
    LocalMux I__2261 (
            .O(N__9518),
            .I(N__9479));
    LocalMux I__2260 (
            .O(N__9515),
            .I(N__9464));
    LocalMux I__2259 (
            .O(N__9512),
            .I(N__9461));
    LocalMux I__2258 (
            .O(N__9509),
            .I(N__9457));
    LocalMux I__2257 (
            .O(N__9506),
            .I(N__9454));
    LocalMux I__2256 (
            .O(N__9503),
            .I(N__9442));
    SRMux I__2255 (
            .O(N__9502),
            .I(N__9343));
    SRMux I__2254 (
            .O(N__9501),
            .I(N__9343));
    SRMux I__2253 (
            .O(N__9500),
            .I(N__9343));
    SRMux I__2252 (
            .O(N__9499),
            .I(N__9343));
    SRMux I__2251 (
            .O(N__9498),
            .I(N__9343));
    SRMux I__2250 (
            .O(N__9497),
            .I(N__9343));
    SRMux I__2249 (
            .O(N__9496),
            .I(N__9343));
    SRMux I__2248 (
            .O(N__9495),
            .I(N__9343));
    SRMux I__2247 (
            .O(N__9494),
            .I(N__9343));
    SRMux I__2246 (
            .O(N__9493),
            .I(N__9343));
    SRMux I__2245 (
            .O(N__9492),
            .I(N__9343));
    SRMux I__2244 (
            .O(N__9491),
            .I(N__9343));
    SRMux I__2243 (
            .O(N__9490),
            .I(N__9343));
    SRMux I__2242 (
            .O(N__9489),
            .I(N__9343));
    SRMux I__2241 (
            .O(N__9488),
            .I(N__9343));
    SRMux I__2240 (
            .O(N__9487),
            .I(N__9343));
    SRMux I__2239 (
            .O(N__9486),
            .I(N__9343));
    SRMux I__2238 (
            .O(N__9485),
            .I(N__9343));
    SRMux I__2237 (
            .O(N__9484),
            .I(N__9343));
    SRMux I__2236 (
            .O(N__9483),
            .I(N__9343));
    SRMux I__2235 (
            .O(N__9482),
            .I(N__9343));
    Glb2LocalMux I__2234 (
            .O(N__9479),
            .I(N__9343));
    SRMux I__2233 (
            .O(N__9478),
            .I(N__9343));
    SRMux I__2232 (
            .O(N__9477),
            .I(N__9343));
    SRMux I__2231 (
            .O(N__9476),
            .I(N__9343));
    SRMux I__2230 (
            .O(N__9475),
            .I(N__9343));
    SRMux I__2229 (
            .O(N__9474),
            .I(N__9343));
    SRMux I__2228 (
            .O(N__9473),
            .I(N__9343));
    SRMux I__2227 (
            .O(N__9472),
            .I(N__9343));
    SRMux I__2226 (
            .O(N__9471),
            .I(N__9343));
    SRMux I__2225 (
            .O(N__9470),
            .I(N__9343));
    SRMux I__2224 (
            .O(N__9469),
            .I(N__9343));
    SRMux I__2223 (
            .O(N__9468),
            .I(N__9343));
    SRMux I__2222 (
            .O(N__9467),
            .I(N__9343));
    Glb2LocalMux I__2221 (
            .O(N__9464),
            .I(N__9343));
    Glb2LocalMux I__2220 (
            .O(N__9461),
            .I(N__9343));
    SRMux I__2219 (
            .O(N__9460),
            .I(N__9343));
    Glb2LocalMux I__2218 (
            .O(N__9457),
            .I(N__9343));
    Glb2LocalMux I__2217 (
            .O(N__9454),
            .I(N__9343));
    SRMux I__2216 (
            .O(N__9453),
            .I(N__9343));
    SRMux I__2215 (
            .O(N__9452),
            .I(N__9343));
    SRMux I__2214 (
            .O(N__9451),
            .I(N__9343));
    SRMux I__2213 (
            .O(N__9450),
            .I(N__9343));
    SRMux I__2212 (
            .O(N__9449),
            .I(N__9343));
    SRMux I__2211 (
            .O(N__9448),
            .I(N__9343));
    SRMux I__2210 (
            .O(N__9447),
            .I(N__9343));
    SRMux I__2209 (
            .O(N__9446),
            .I(N__9343));
    SRMux I__2208 (
            .O(N__9445),
            .I(N__9343));
    Glb2LocalMux I__2207 (
            .O(N__9442),
            .I(N__9343));
    GlobalMux I__2206 (
            .O(N__9343),
            .I(N__9340));
    gio2CtrlBuf I__2205 (
            .O(N__9340),
            .I(RESETn_c_i_g));
    CascadeMux I__2204 (
            .O(N__9337),
            .I(N__9334));
    InMux I__2203 (
            .O(N__9334),
            .I(N__9331));
    LocalMux I__2202 (
            .O(N__9331),
            .I(N__9328));
    Span4Mux_h I__2201 (
            .O(N__9328),
            .I(N__9325));
    Odrv4 I__2200 (
            .O(N__9325),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2199 (
            .O(N__9322),
            .I(N__9319));
    LocalMux I__2198 (
            .O(N__9319),
            .I(N__9316));
    Odrv4 I__2197 (
            .O(N__9316),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2196 (
            .O(N__9313),
            .I(N__9310));
    LocalMux I__2195 (
            .O(N__9310),
            .I(N__9300));
    ClkMux I__2194 (
            .O(N__9309),
            .I(N__9283));
    ClkMux I__2193 (
            .O(N__9308),
            .I(N__9283));
    ClkMux I__2192 (
            .O(N__9307),
            .I(N__9283));
    ClkMux I__2191 (
            .O(N__9306),
            .I(N__9283));
    ClkMux I__2190 (
            .O(N__9305),
            .I(N__9283));
    ClkMux I__2189 (
            .O(N__9304),
            .I(N__9283));
    ClkMux I__2188 (
            .O(N__9303),
            .I(N__9283));
    Glb2LocalMux I__2187 (
            .O(N__9300),
            .I(N__9283));
    GlobalMux I__2186 (
            .O(N__9283),
            .I(N__9280));
    gio2CtrlBuf I__2185 (
            .O(N__9280),
            .I(C1_c_g));
    InMux I__2184 (
            .O(N__9277),
            .I(N__9272));
    InMux I__2183 (
            .O(N__9276),
            .I(N__9269));
    InMux I__2182 (
            .O(N__9275),
            .I(N__9266));
    LocalMux I__2181 (
            .O(N__9272),
            .I(N__9263));
    LocalMux I__2180 (
            .O(N__9269),
            .I(N__9260));
    LocalMux I__2179 (
            .O(N__9266),
            .I(N__9257));
    Sp12to4 I__2178 (
            .O(N__9263),
            .I(N__9254));
    Sp12to4 I__2177 (
            .O(N__9260),
            .I(N__9251));
    Span4Mux_v I__2176 (
            .O(N__9257),
            .I(N__9248));
    Span12Mux_v I__2175 (
            .O(N__9254),
            .I(N__9245));
    Span12Mux_h I__2174 (
            .O(N__9251),
            .I(N__9242));
    Sp12to4 I__2173 (
            .O(N__9248),
            .I(N__9239));
    Span12Mux_h I__2172 (
            .O(N__9245),
            .I(N__9234));
    Span12Mux_v I__2171 (
            .O(N__9242),
            .I(N__9234));
    Span12Mux_h I__2170 (
            .O(N__9239),
            .I(N__9231));
    Odrv12 I__2169 (
            .O(N__9234),
            .I(DBRn_c));
    Odrv12 I__2168 (
            .O(N__9231),
            .I(DBRn_c));
    InMux I__2167 (
            .O(N__9226),
            .I(N__9223));
    LocalMux I__2166 (
            .O(N__9223),
            .I(N__9220));
    Odrv12 I__2165 (
            .O(N__9220),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2164 (
            .O(N__9217),
            .I(N__9214));
    LocalMux I__2163 (
            .O(N__9214),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2162 (
            .O(N__9211),
            .I(N__9208));
    LocalMux I__2161 (
            .O(N__9208),
            .I(N__9205));
    Span4Mux_v I__2160 (
            .O(N__9205),
            .I(N__9201));
    InMux I__2159 (
            .O(N__9204),
            .I(N__9198));
    Sp12to4 I__2158 (
            .O(N__9201),
            .I(N__9193));
    LocalMux I__2157 (
            .O(N__9198),
            .I(N__9193));
    Span12Mux_h I__2156 (
            .O(N__9193),
            .I(N__9190));
    Odrv12 I__2155 (
            .O(N__9190),
            .I(DRA_c_7));
    InMux I__2154 (
            .O(N__9187),
            .I(N__9184));
    LocalMux I__2153 (
            .O(N__9184),
            .I(N__9181));
    Span4Mux_h I__2152 (
            .O(N__9181),
            .I(N__9178));
    Odrv4 I__2151 (
            .O(N__9178),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__2150 (
            .O(N__9175),
            .I(N__9171));
    InMux I__2149 (
            .O(N__9174),
            .I(N__9168));
    LocalMux I__2148 (
            .O(N__9171),
            .I(N__9163));
    LocalMux I__2147 (
            .O(N__9168),
            .I(N__9163));
    Span4Mux_h I__2146 (
            .O(N__9163),
            .I(N__9160));
    Sp12to4 I__2145 (
            .O(N__9160),
            .I(N__9157));
    Span12Mux_v I__2144 (
            .O(N__9157),
            .I(N__9154));
    Odrv12 I__2143 (
            .O(N__9154),
            .I(DRA_c_8));
    InMux I__2142 (
            .O(N__9151),
            .I(N__9148));
    LocalMux I__2141 (
            .O(N__9148),
            .I(N__9145));
    Span4Mux_h I__2140 (
            .O(N__9145),
            .I(N__9142));
    Odrv4 I__2139 (
            .O(N__9142),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    InMux I__2138 (
            .O(N__9139),
            .I(N__9135));
    InMux I__2137 (
            .O(N__9138),
            .I(N__9132));
    LocalMux I__2136 (
            .O(N__9135),
            .I(N__9127));
    LocalMux I__2135 (
            .O(N__9132),
            .I(N__9127));
    Span4Mux_v I__2134 (
            .O(N__9127),
            .I(N__9124));
    Sp12to4 I__2133 (
            .O(N__9124),
            .I(N__9121));
    Span12Mux_h I__2132 (
            .O(N__9121),
            .I(N__9118));
    Odrv12 I__2131 (
            .O(N__9118),
            .I(DRA_c_5));
    InMux I__2130 (
            .O(N__9115),
            .I(N__9109));
    InMux I__2129 (
            .O(N__9114),
            .I(N__9109));
    LocalMux I__2128 (
            .O(N__9109),
            .I(N__9106));
    Span4Mux_h I__2127 (
            .O(N__9106),
            .I(N__9103));
    Odrv4 I__2126 (
            .O(N__9103),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__2125 (
            .O(N__9100),
            .I(N__9097));
    LocalMux I__2124 (
            .O(N__9097),
            .I(N__9087));
    ClkMux I__2123 (
            .O(N__9096),
            .I(N__9070));
    ClkMux I__2122 (
            .O(N__9095),
            .I(N__9070));
    ClkMux I__2121 (
            .O(N__9094),
            .I(N__9070));
    ClkMux I__2120 (
            .O(N__9093),
            .I(N__9070));
    ClkMux I__2119 (
            .O(N__9092),
            .I(N__9070));
    ClkMux I__2118 (
            .O(N__9091),
            .I(N__9070));
    ClkMux I__2117 (
            .O(N__9090),
            .I(N__9070));
    Glb2LocalMux I__2116 (
            .O(N__9087),
            .I(N__9070));
    GlobalMux I__2115 (
            .O(N__9070),
            .I(N__9067));
    gio2CtrlBuf I__2114 (
            .O(N__9067),
            .I(C3_c_g));
    InMux I__2113 (
            .O(N__9064),
            .I(N__9059));
    InMux I__2112 (
            .O(N__9063),
            .I(N__9054));
    InMux I__2111 (
            .O(N__9062),
            .I(N__9054));
    LocalMux I__2110 (
            .O(N__9059),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__2109 (
            .O(N__9054),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    CascadeMux I__2108 (
            .O(N__9049),
            .I(N__9045));
    InMux I__2107 (
            .O(N__9048),
            .I(N__9042));
    InMux I__2106 (
            .O(N__9045),
            .I(N__9039));
    LocalMux I__2105 (
            .O(N__9042),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__2104 (
            .O(N__9039),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    InMux I__2103 (
            .O(N__9034),
            .I(N__9030));
    InMux I__2102 (
            .O(N__9033),
            .I(N__9027));
    LocalMux I__2101 (
            .O(N__9030),
            .I(N__9022));
    LocalMux I__2100 (
            .O(N__9027),
            .I(N__9017));
    InMux I__2099 (
            .O(N__9026),
            .I(N__9014));
    InMux I__2098 (
            .O(N__9025),
            .I(N__9011));
    Span12Mux_v I__2097 (
            .O(N__9022),
            .I(N__9008));
    InMux I__2096 (
            .O(N__9021),
            .I(N__9003));
    InMux I__2095 (
            .O(N__9020),
            .I(N__9003));
    Span4Mux_h I__2094 (
            .O(N__9017),
            .I(N__8996));
    LocalMux I__2093 (
            .O(N__9014),
            .I(N__8996));
    LocalMux I__2092 (
            .O(N__9011),
            .I(N__8996));
    Odrv12 I__2091 (
            .O(N__9008),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__2090 (
            .O(N__9003),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2089 (
            .O(N__8996),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__2088 (
            .O(N__8989),
            .I(N__8986));
    LocalMux I__2087 (
            .O(N__8986),
            .I(N__8983));
    Span12Mux_s8_v I__2086 (
            .O(N__8983),
            .I(N__8980));
    Odrv12 I__2085 (
            .O(N__8980),
            .I(RASn_c));
    IoInMux I__2084 (
            .O(N__8977),
            .I(N__8974));
    LocalMux I__2083 (
            .O(N__8974),
            .I(N__8971));
    IoSpan4Mux I__2082 (
            .O(N__8971),
            .I(N__8968));
    Span4Mux_s2_v I__2081 (
            .O(N__8968),
            .I(N__8965));
    Sp12to4 I__2080 (
            .O(N__8965),
            .I(N__8962));
    Span12Mux_s10_v I__2079 (
            .O(N__8962),
            .I(N__8959));
    Odrv12 I__2078 (
            .O(N__8959),
            .I(CASn_c));
    InMux I__2077 (
            .O(N__8956),
            .I(N__8953));
    LocalMux I__2076 (
            .O(N__8953),
            .I(N__8950));
    Span4Mux_v I__2075 (
            .O(N__8950),
            .I(N__8946));
    InMux I__2074 (
            .O(N__8949),
            .I(N__8943));
    Sp12to4 I__2073 (
            .O(N__8946),
            .I(N__8938));
    LocalMux I__2072 (
            .O(N__8943),
            .I(N__8938));
    Span12Mux_h I__2071 (
            .O(N__8938),
            .I(N__8935));
    Odrv12 I__2070 (
            .O(N__8935),
            .I(DRA_c_6));
    CascadeMux I__2069 (
            .O(N__8932),
            .I(N__8929));
    InMux I__2068 (
            .O(N__8929),
            .I(N__8926));
    LocalMux I__2067 (
            .O(N__8926),
            .I(N__8923));
    Odrv4 I__2066 (
            .O(N__8923),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2065 (
            .O(N__8920),
            .I(N__8916));
    InMux I__2064 (
            .O(N__8919),
            .I(N__8913));
    LocalMux I__2063 (
            .O(N__8916),
            .I(N__8906));
    LocalMux I__2062 (
            .O(N__8913),
            .I(N__8903));
    InMux I__2061 (
            .O(N__8912),
            .I(N__8900));
    InMux I__2060 (
            .O(N__8911),
            .I(N__8897));
    InMux I__2059 (
            .O(N__8910),
            .I(N__8894));
    InMux I__2058 (
            .O(N__8909),
            .I(N__8891));
    Span4Mux_h I__2057 (
            .O(N__8906),
            .I(N__8885));
    Span4Mux_v I__2056 (
            .O(N__8903),
            .I(N__8882));
    LocalMux I__2055 (
            .O(N__8900),
            .I(N__8877));
    LocalMux I__2054 (
            .O(N__8897),
            .I(N__8877));
    LocalMux I__2053 (
            .O(N__8894),
            .I(N__8872));
    LocalMux I__2052 (
            .O(N__8891),
            .I(N__8872));
    InMux I__2051 (
            .O(N__8890),
            .I(N__8867));
    InMux I__2050 (
            .O(N__8889),
            .I(N__8867));
    InMux I__2049 (
            .O(N__8888),
            .I(N__8864));
    Odrv4 I__2048 (
            .O(N__8885),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__2047 (
            .O(N__8882),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__2046 (
            .O(N__8877),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__2045 (
            .O(N__8872),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__2044 (
            .O(N__8867),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__2043 (
            .O(N__8864),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    CascadeMux I__2042 (
            .O(N__8851),
            .I(N__8846));
    CascadeMux I__2041 (
            .O(N__8850),
            .I(N__8841));
    CascadeMux I__2040 (
            .O(N__8849),
            .I(N__8837));
    InMux I__2039 (
            .O(N__8846),
            .I(N__8834));
    InMux I__2038 (
            .O(N__8845),
            .I(N__8831));
    InMux I__2037 (
            .O(N__8844),
            .I(N__8826));
    InMux I__2036 (
            .O(N__8841),
            .I(N__8826));
    InMux I__2035 (
            .O(N__8840),
            .I(N__8821));
    InMux I__2034 (
            .O(N__8837),
            .I(N__8821));
    LocalMux I__2033 (
            .O(N__8834),
            .I(N__8818));
    LocalMux I__2032 (
            .O(N__8831),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    LocalMux I__2031 (
            .O(N__8826),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    LocalMux I__2030 (
            .O(N__8821),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    Odrv4 I__2029 (
            .O(N__8818),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    IoInMux I__2028 (
            .O(N__8809),
            .I(N__8806));
    LocalMux I__2027 (
            .O(N__8806),
            .I(N__8803));
    IoSpan4Mux I__2026 (
            .O(N__8803),
            .I(N__8800));
    Sp12to4 I__2025 (
            .O(N__8800),
            .I(N__8797));
    Span12Mux_s9_h I__2024 (
            .O(N__8797),
            .I(N__8794));
    Span12Mux_v I__2023 (
            .O(N__8794),
            .I(N__8791));
    Odrv12 I__2022 (
            .O(N__8791),
            .I(CMA_c_4));
    InMux I__2021 (
            .O(N__8788),
            .I(N__8785));
    LocalMux I__2020 (
            .O(N__8785),
            .I(N__8755));
    ClkMux I__2019 (
            .O(N__8784),
            .I(N__8674));
    ClkMux I__2018 (
            .O(N__8783),
            .I(N__8674));
    ClkMux I__2017 (
            .O(N__8782),
            .I(N__8674));
    ClkMux I__2016 (
            .O(N__8781),
            .I(N__8674));
    ClkMux I__2015 (
            .O(N__8780),
            .I(N__8674));
    ClkMux I__2014 (
            .O(N__8779),
            .I(N__8674));
    ClkMux I__2013 (
            .O(N__8778),
            .I(N__8674));
    ClkMux I__2012 (
            .O(N__8777),
            .I(N__8674));
    ClkMux I__2011 (
            .O(N__8776),
            .I(N__8674));
    ClkMux I__2010 (
            .O(N__8775),
            .I(N__8674));
    ClkMux I__2009 (
            .O(N__8774),
            .I(N__8674));
    ClkMux I__2008 (
            .O(N__8773),
            .I(N__8674));
    ClkMux I__2007 (
            .O(N__8772),
            .I(N__8674));
    ClkMux I__2006 (
            .O(N__8771),
            .I(N__8674));
    ClkMux I__2005 (
            .O(N__8770),
            .I(N__8674));
    ClkMux I__2004 (
            .O(N__8769),
            .I(N__8674));
    ClkMux I__2003 (
            .O(N__8768),
            .I(N__8674));
    ClkMux I__2002 (
            .O(N__8767),
            .I(N__8674));
    ClkMux I__2001 (
            .O(N__8766),
            .I(N__8674));
    ClkMux I__2000 (
            .O(N__8765),
            .I(N__8674));
    ClkMux I__1999 (
            .O(N__8764),
            .I(N__8674));
    ClkMux I__1998 (
            .O(N__8763),
            .I(N__8674));
    ClkMux I__1997 (
            .O(N__8762),
            .I(N__8674));
    ClkMux I__1996 (
            .O(N__8761),
            .I(N__8674));
    ClkMux I__1995 (
            .O(N__8760),
            .I(N__8674));
    ClkMux I__1994 (
            .O(N__8759),
            .I(N__8674));
    ClkMux I__1993 (
            .O(N__8758),
            .I(N__8674));
    Glb2LocalMux I__1992 (
            .O(N__8755),
            .I(N__8674));
    ClkMux I__1991 (
            .O(N__8754),
            .I(N__8674));
    ClkMux I__1990 (
            .O(N__8753),
            .I(N__8674));
    ClkMux I__1989 (
            .O(N__8752),
            .I(N__8674));
    ClkMux I__1988 (
            .O(N__8751),
            .I(N__8674));
    ClkMux I__1987 (
            .O(N__8750),
            .I(N__8674));
    ClkMux I__1986 (
            .O(N__8749),
            .I(N__8674));
    ClkMux I__1985 (
            .O(N__8748),
            .I(N__8674));
    ClkMux I__1984 (
            .O(N__8747),
            .I(N__8674));
    GlobalMux I__1983 (
            .O(N__8674),
            .I(CLK80_OUT));
    CEMux I__1982 (
            .O(N__8671),
            .I(N__8665));
    CEMux I__1981 (
            .O(N__8670),
            .I(N__8661));
    CEMux I__1980 (
            .O(N__8669),
            .I(N__8658));
    CEMux I__1979 (
            .O(N__8668),
            .I(N__8655));
    LocalMux I__1978 (
            .O(N__8665),
            .I(N__8651));
    CEMux I__1977 (
            .O(N__8664),
            .I(N__8648));
    LocalMux I__1976 (
            .O(N__8661),
            .I(N__8645));
    LocalMux I__1975 (
            .O(N__8658),
            .I(N__8642));
    LocalMux I__1974 (
            .O(N__8655),
            .I(N__8639));
    CEMux I__1973 (
            .O(N__8654),
            .I(N__8636));
    Span4Mux_h I__1972 (
            .O(N__8651),
            .I(N__8631));
    LocalMux I__1971 (
            .O(N__8648),
            .I(N__8631));
    Span4Mux_v I__1970 (
            .O(N__8645),
            .I(N__8628));
    Span4Mux_v I__1969 (
            .O(N__8642),
            .I(N__8625));
    Span4Mux_h I__1968 (
            .O(N__8639),
            .I(N__8620));
    LocalMux I__1967 (
            .O(N__8636),
            .I(N__8620));
    Span4Mux_v I__1966 (
            .O(N__8631),
            .I(N__8617));
    Odrv4 I__1965 (
            .O(N__8628),
            .I(\U712_CHIP_RAM.un1_CMA30_0_i_0 ));
    Odrv4 I__1964 (
            .O(N__8625),
            .I(\U712_CHIP_RAM.un1_CMA30_0_i_0 ));
    Odrv4 I__1963 (
            .O(N__8620),
            .I(\U712_CHIP_RAM.un1_CMA30_0_i_0 ));
    Odrv4 I__1962 (
            .O(N__8617),
            .I(\U712_CHIP_RAM.un1_CMA30_0_i_0 ));
    InMux I__1961 (
            .O(N__8608),
            .I(N__8605));
    LocalMux I__1960 (
            .O(N__8605),
            .I(N__8602));
    Span4Mux_v I__1959 (
            .O(N__8602),
            .I(N__8599));
    Sp12to4 I__1958 (
            .O(N__8599),
            .I(N__8596));
    Span12Mux_h I__1957 (
            .O(N__8596),
            .I(N__8593));
    Odrv12 I__1956 (
            .O(N__8593),
            .I(A_c_13));
    InMux I__1955 (
            .O(N__8590),
            .I(N__8587));
    LocalMux I__1954 (
            .O(N__8587),
            .I(N__8584));
    Span4Mux_v I__1953 (
            .O(N__8584),
            .I(N__8581));
    Sp12to4 I__1952 (
            .O(N__8581),
            .I(N__8578));
    Span12Mux_h I__1951 (
            .O(N__8578),
            .I(N__8575));
    Odrv12 I__1950 (
            .O(N__8575),
            .I(A_c_6));
    CascadeMux I__1949 (
            .O(N__8572),
            .I(N__8566));
    CascadeMux I__1948 (
            .O(N__8571),
            .I(N__8558));
    CascadeMux I__1947 (
            .O(N__8570),
            .I(N__8555));
    InMux I__1946 (
            .O(N__8569),
            .I(N__8549));
    InMux I__1945 (
            .O(N__8566),
            .I(N__8542));
    InMux I__1944 (
            .O(N__8565),
            .I(N__8539));
    InMux I__1943 (
            .O(N__8564),
            .I(N__8536));
    InMux I__1942 (
            .O(N__8563),
            .I(N__8529));
    InMux I__1941 (
            .O(N__8562),
            .I(N__8529));
    InMux I__1940 (
            .O(N__8561),
            .I(N__8529));
    InMux I__1939 (
            .O(N__8558),
            .I(N__8516));
    InMux I__1938 (
            .O(N__8555),
            .I(N__8516));
    InMux I__1937 (
            .O(N__8554),
            .I(N__8516));
    InMux I__1936 (
            .O(N__8553),
            .I(N__8511));
    InMux I__1935 (
            .O(N__8552),
            .I(N__8511));
    LocalMux I__1934 (
            .O(N__8549),
            .I(N__8508));
    InMux I__1933 (
            .O(N__8548),
            .I(N__8505));
    InMux I__1932 (
            .O(N__8547),
            .I(N__8500));
    InMux I__1931 (
            .O(N__8546),
            .I(N__8500));
    InMux I__1930 (
            .O(N__8545),
            .I(N__8496));
    LocalMux I__1929 (
            .O(N__8542),
            .I(N__8487));
    LocalMux I__1928 (
            .O(N__8539),
            .I(N__8487));
    LocalMux I__1927 (
            .O(N__8536),
            .I(N__8487));
    LocalMux I__1926 (
            .O(N__8529),
            .I(N__8487));
    InMux I__1925 (
            .O(N__8528),
            .I(N__8484));
    InMux I__1924 (
            .O(N__8527),
            .I(N__8473));
    InMux I__1923 (
            .O(N__8526),
            .I(N__8473));
    InMux I__1922 (
            .O(N__8525),
            .I(N__8473));
    InMux I__1921 (
            .O(N__8524),
            .I(N__8473));
    InMux I__1920 (
            .O(N__8523),
            .I(N__8473));
    LocalMux I__1919 (
            .O(N__8516),
            .I(N__8468));
    LocalMux I__1918 (
            .O(N__8511),
            .I(N__8468));
    Span4Mux_h I__1917 (
            .O(N__8508),
            .I(N__8461));
    LocalMux I__1916 (
            .O(N__8505),
            .I(N__8461));
    LocalMux I__1915 (
            .O(N__8500),
            .I(N__8461));
    InMux I__1914 (
            .O(N__8499),
            .I(N__8458));
    LocalMux I__1913 (
            .O(N__8496),
            .I(N__8455));
    Span4Mux_v I__1912 (
            .O(N__8487),
            .I(N__8452));
    LocalMux I__1911 (
            .O(N__8484),
            .I(N__8447));
    LocalMux I__1910 (
            .O(N__8473),
            .I(N__8447));
    Span4Mux_h I__1909 (
            .O(N__8468),
            .I(N__8438));
    Span4Mux_v I__1908 (
            .O(N__8461),
            .I(N__8438));
    LocalMux I__1907 (
            .O(N__8458),
            .I(N__8438));
    Span4Mux_h I__1906 (
            .O(N__8455),
            .I(N__8438));
    Odrv4 I__1905 (
            .O(N__8452),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__1904 (
            .O(N__8447),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1903 (
            .O(N__8438),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    InMux I__1902 (
            .O(N__8431),
            .I(N__8424));
    InMux I__1901 (
            .O(N__8430),
            .I(N__8424));
    CascadeMux I__1900 (
            .O(N__8429),
            .I(N__8412));
    LocalMux I__1899 (
            .O(N__8424),
            .I(N__8409));
    InMux I__1898 (
            .O(N__8423),
            .I(N__8406));
    CascadeMux I__1897 (
            .O(N__8422),
            .I(N__8403));
    InMux I__1896 (
            .O(N__8421),
            .I(N__8397));
    InMux I__1895 (
            .O(N__8420),
            .I(N__8391));
    CascadeMux I__1894 (
            .O(N__8419),
            .I(N__8384));
    InMux I__1893 (
            .O(N__8418),
            .I(N__8381));
    InMux I__1892 (
            .O(N__8417),
            .I(N__8378));
    InMux I__1891 (
            .O(N__8416),
            .I(N__8371));
    InMux I__1890 (
            .O(N__8415),
            .I(N__8371));
    InMux I__1889 (
            .O(N__8412),
            .I(N__8371));
    Span4Mux_v I__1888 (
            .O(N__8409),
            .I(N__8366));
    LocalMux I__1887 (
            .O(N__8406),
            .I(N__8366));
    InMux I__1886 (
            .O(N__8403),
            .I(N__8359));
    InMux I__1885 (
            .O(N__8402),
            .I(N__8359));
    InMux I__1884 (
            .O(N__8401),
            .I(N__8359));
    InMux I__1883 (
            .O(N__8400),
            .I(N__8356));
    LocalMux I__1882 (
            .O(N__8397),
            .I(N__8353));
    InMux I__1881 (
            .O(N__8396),
            .I(N__8346));
    InMux I__1880 (
            .O(N__8395),
            .I(N__8346));
    InMux I__1879 (
            .O(N__8394),
            .I(N__8346));
    LocalMux I__1878 (
            .O(N__8391),
            .I(N__8343));
    InMux I__1877 (
            .O(N__8390),
            .I(N__8336));
    InMux I__1876 (
            .O(N__8389),
            .I(N__8336));
    InMux I__1875 (
            .O(N__8388),
            .I(N__8336));
    InMux I__1874 (
            .O(N__8387),
            .I(N__8331));
    InMux I__1873 (
            .O(N__8384),
            .I(N__8331));
    LocalMux I__1872 (
            .O(N__8381),
            .I(N__8327));
    LocalMux I__1871 (
            .O(N__8378),
            .I(N__8318));
    LocalMux I__1870 (
            .O(N__8371),
            .I(N__8318));
    Span4Mux_h I__1869 (
            .O(N__8366),
            .I(N__8318));
    LocalMux I__1868 (
            .O(N__8359),
            .I(N__8318));
    LocalMux I__1867 (
            .O(N__8356),
            .I(N__8311));
    Span4Mux_v I__1866 (
            .O(N__8353),
            .I(N__8311));
    LocalMux I__1865 (
            .O(N__8346),
            .I(N__8311));
    Span4Mux_v I__1864 (
            .O(N__8343),
            .I(N__8304));
    LocalMux I__1863 (
            .O(N__8336),
            .I(N__8304));
    LocalMux I__1862 (
            .O(N__8331),
            .I(N__8304));
    InMux I__1861 (
            .O(N__8330),
            .I(N__8301));
    Span4Mux_v I__1860 (
            .O(N__8327),
            .I(N__8296));
    Span4Mux_v I__1859 (
            .O(N__8318),
            .I(N__8296));
    Span4Mux_h I__1858 (
            .O(N__8311),
            .I(N__8293));
    Odrv4 I__1857 (
            .O(N__8304),
            .I(CPU_CYCLEm));
    LocalMux I__1856 (
            .O(N__8301),
            .I(CPU_CYCLEm));
    Odrv4 I__1855 (
            .O(N__8296),
            .I(CPU_CYCLEm));
    Odrv4 I__1854 (
            .O(N__8293),
            .I(CPU_CYCLEm));
    CascadeMux I__1853 (
            .O(N__8284),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ));
    InMux I__1852 (
            .O(N__8281),
            .I(N__8278));
    LocalMux I__1851 (
            .O(N__8278),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    InMux I__1850 (
            .O(N__8275),
            .I(N__8272));
    LocalMux I__1849 (
            .O(N__8272),
            .I(N__8269));
    Span4Mux_v I__1848 (
            .O(N__8269),
            .I(N__8265));
    InMux I__1847 (
            .O(N__8268),
            .I(N__8262));
    Sp12to4 I__1846 (
            .O(N__8265),
            .I(N__8259));
    LocalMux I__1845 (
            .O(N__8262),
            .I(N__8256));
    Span12Mux_h I__1844 (
            .O(N__8259),
            .I(N__8253));
    Span12Mux_v I__1843 (
            .O(N__8256),
            .I(N__8250));
    Span12Mux_v I__1842 (
            .O(N__8253),
            .I(N__8245));
    Span12Mux_h I__1841 (
            .O(N__8250),
            .I(N__8245));
    Odrv12 I__1840 (
            .O(N__8245),
            .I(DRA_c_0));
    CascadeMux I__1839 (
            .O(N__8242),
            .I(N__8239));
    InMux I__1838 (
            .O(N__8239),
            .I(N__8236));
    LocalMux I__1837 (
            .O(N__8236),
            .I(N__8233));
    Span4Mux_h I__1836 (
            .O(N__8233),
            .I(N__8230));
    Odrv4 I__1835 (
            .O(N__8230),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__1834 (
            .O(N__8227),
            .I(N__8223));
    InMux I__1833 (
            .O(N__8226),
            .I(N__8220));
    LocalMux I__1832 (
            .O(N__8223),
            .I(N__8215));
    LocalMux I__1831 (
            .O(N__8220),
            .I(N__8215));
    Span4Mux_v I__1830 (
            .O(N__8215),
            .I(N__8212));
    Span4Mux_v I__1829 (
            .O(N__8212),
            .I(N__8209));
    Sp12to4 I__1828 (
            .O(N__8209),
            .I(N__8206));
    Span12Mux_h I__1827 (
            .O(N__8206),
            .I(N__8203));
    Odrv12 I__1826 (
            .O(N__8203),
            .I(DRA_c_3));
    InMux I__1825 (
            .O(N__8200),
            .I(N__8197));
    LocalMux I__1824 (
            .O(N__8197),
            .I(N__8194));
    Span4Mux_v I__1823 (
            .O(N__8194),
            .I(N__8191));
    Odrv4 I__1822 (
            .O(N__8191),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1821 (
            .O(N__8188),
            .I(N__8185));
    LocalMux I__1820 (
            .O(N__8185),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__1819 (
            .O(N__8182),
            .I(N__8179));
    LocalMux I__1818 (
            .O(N__8179),
            .I(N__8175));
    InMux I__1817 (
            .O(N__8178),
            .I(N__8172));
    Span4Mux_h I__1816 (
            .O(N__8175),
            .I(N__8167));
    LocalMux I__1815 (
            .O(N__8172),
            .I(N__8167));
    Sp12to4 I__1814 (
            .O(N__8167),
            .I(N__8164));
    Span12Mux_v I__1813 (
            .O(N__8164),
            .I(N__8161));
    Span12Mux_h I__1812 (
            .O(N__8161),
            .I(N__8158));
    Odrv12 I__1811 (
            .O(N__8158),
            .I(DRA_c_1));
    InMux I__1810 (
            .O(N__8155),
            .I(N__8149));
    InMux I__1809 (
            .O(N__8154),
            .I(N__8149));
    LocalMux I__1808 (
            .O(N__8149),
            .I(N__8146));
    Odrv4 I__1807 (
            .O(N__8146),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    CascadeMux I__1806 (
            .O(N__8143),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0_cascade_ ));
    InMux I__1805 (
            .O(N__8140),
            .I(N__8137));
    LocalMux I__1804 (
            .O(N__8137),
            .I(N__8131));
    InMux I__1803 (
            .O(N__8136),
            .I(N__8128));
    InMux I__1802 (
            .O(N__8135),
            .I(N__8125));
    InMux I__1801 (
            .O(N__8134),
            .I(N__8122));
    Span4Mux_h I__1800 (
            .O(N__8131),
            .I(N__8117));
    LocalMux I__1799 (
            .O(N__8128),
            .I(N__8117));
    LocalMux I__1798 (
            .O(N__8125),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__1797 (
            .O(N__8122),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    Odrv4 I__1796 (
            .O(N__8117),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    InMux I__1795 (
            .O(N__8110),
            .I(N__8107));
    LocalMux I__1794 (
            .O(N__8107),
            .I(N__8104));
    Span4Mux_v I__1793 (
            .O(N__8104),
            .I(N__8100));
    InMux I__1792 (
            .O(N__8103),
            .I(N__8096));
    Span4Mux_h I__1791 (
            .O(N__8100),
            .I(N__8093));
    InMux I__1790 (
            .O(N__8099),
            .I(N__8090));
    LocalMux I__1789 (
            .O(N__8096),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    Odrv4 I__1788 (
            .O(N__8093),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__1787 (
            .O(N__8090),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__1786 (
            .O(N__8083),
            .I(N__8077));
    InMux I__1785 (
            .O(N__8082),
            .I(N__8077));
    LocalMux I__1784 (
            .O(N__8077),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__1783 (
            .O(N__8074),
            .I(N__8071));
    LocalMux I__1782 (
            .O(N__8071),
            .I(N__8068));
    Span4Mux_v I__1781 (
            .O(N__8068),
            .I(N__8065));
    Span4Mux_v I__1780 (
            .O(N__8065),
            .I(N__8059));
    InMux I__1779 (
            .O(N__8064),
            .I(N__8054));
    InMux I__1778 (
            .O(N__8063),
            .I(N__8054));
    InMux I__1777 (
            .O(N__8062),
            .I(N__8051));
    Sp12to4 I__1776 (
            .O(N__8059),
            .I(N__8048));
    LocalMux I__1775 (
            .O(N__8054),
            .I(N__8043));
    LocalMux I__1774 (
            .O(N__8051),
            .I(N__8043));
    Span12Mux_h I__1773 (
            .O(N__8048),
            .I(N__8038));
    Span12Mux_v I__1772 (
            .O(N__8043),
            .I(N__8038));
    Odrv12 I__1771 (
            .O(N__8038),
            .I(CLK40_OUT_i));
    CascadeMux I__1770 (
            .O(N__8035),
            .I(N__8032));
    InMux I__1769 (
            .O(N__8032),
            .I(N__8026));
    InMux I__1768 (
            .O(N__8031),
            .I(N__8019));
    InMux I__1767 (
            .O(N__8030),
            .I(N__8019));
    InMux I__1766 (
            .O(N__8029),
            .I(N__8019));
    LocalMux I__1765 (
            .O(N__8026),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1764 (
            .O(N__8019),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    IoInMux I__1763 (
            .O(N__8014),
            .I(N__8011));
    LocalMux I__1762 (
            .O(N__8011),
            .I(N__8008));
    Span4Mux_s3_h I__1761 (
            .O(N__8008),
            .I(N__8005));
    Span4Mux_v I__1760 (
            .O(N__8005),
            .I(N__8002));
    Span4Mux_v I__1759 (
            .O(N__8002),
            .I(N__7999));
    Sp12to4 I__1758 (
            .O(N__7999),
            .I(N__7995));
    CascadeMux I__1757 (
            .O(N__7998),
            .I(N__7992));
    Span12Mux_h I__1756 (
            .O(N__7995),
            .I(N__7989));
    InMux I__1755 (
            .O(N__7992),
            .I(N__7986));
    Odrv12 I__1754 (
            .O(N__7989),
            .I(TACK_OUTn));
    LocalMux I__1753 (
            .O(N__7986),
            .I(TACK_OUTn));
    CascadeMux I__1752 (
            .O(N__7981),
            .I(N__7974));
    InMux I__1751 (
            .O(N__7980),
            .I(N__7971));
    InMux I__1750 (
            .O(N__7979),
            .I(N__7966));
    InMux I__1749 (
            .O(N__7978),
            .I(N__7966));
    CascadeMux I__1748 (
            .O(N__7977),
            .I(N__7962));
    InMux I__1747 (
            .O(N__7974),
            .I(N__7955));
    LocalMux I__1746 (
            .O(N__7971),
            .I(N__7952));
    LocalMux I__1745 (
            .O(N__7966),
            .I(N__7949));
    InMux I__1744 (
            .O(N__7965),
            .I(N__7946));
    InMux I__1743 (
            .O(N__7962),
            .I(N__7943));
    InMux I__1742 (
            .O(N__7961),
            .I(N__7938));
    InMux I__1741 (
            .O(N__7960),
            .I(N__7938));
    InMux I__1740 (
            .O(N__7959),
            .I(N__7934));
    InMux I__1739 (
            .O(N__7958),
            .I(N__7931));
    LocalMux I__1738 (
            .O(N__7955),
            .I(N__7928));
    Span4Mux_h I__1737 (
            .O(N__7952),
            .I(N__7925));
    Span4Mux_h I__1736 (
            .O(N__7949),
            .I(N__7920));
    LocalMux I__1735 (
            .O(N__7946),
            .I(N__7920));
    LocalMux I__1734 (
            .O(N__7943),
            .I(N__7915));
    LocalMux I__1733 (
            .O(N__7938),
            .I(N__7915));
    InMux I__1732 (
            .O(N__7937),
            .I(N__7912));
    LocalMux I__1731 (
            .O(N__7934),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1730 (
            .O(N__7931),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1729 (
            .O(N__7928),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1728 (
            .O(N__7925),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1727 (
            .O(N__7920),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv12 I__1726 (
            .O(N__7915),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1725 (
            .O(N__7912),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__1724 (
            .O(N__7897),
            .I(N__7893));
    InMux I__1723 (
            .O(N__7896),
            .I(N__7889));
    InMux I__1722 (
            .O(N__7893),
            .I(N__7886));
    InMux I__1721 (
            .O(N__7892),
            .I(N__7880));
    LocalMux I__1720 (
            .O(N__7889),
            .I(N__7875));
    LocalMux I__1719 (
            .O(N__7886),
            .I(N__7875));
    InMux I__1718 (
            .O(N__7885),
            .I(N__7872));
    InMux I__1717 (
            .O(N__7884),
            .I(N__7867));
    InMux I__1716 (
            .O(N__7883),
            .I(N__7867));
    LocalMux I__1715 (
            .O(N__7880),
            .I(\U712_CHIP_RAM.N_312 ));
    Odrv4 I__1714 (
            .O(N__7875),
            .I(\U712_CHIP_RAM.N_312 ));
    LocalMux I__1713 (
            .O(N__7872),
            .I(\U712_CHIP_RAM.N_312 ));
    LocalMux I__1712 (
            .O(N__7867),
            .I(\U712_CHIP_RAM.N_312 ));
    InMux I__1711 (
            .O(N__7858),
            .I(N__7855));
    LocalMux I__1710 (
            .O(N__7855),
            .I(N__7852));
    Odrv4 I__1709 (
            .O(N__7852),
            .I(\U712_CHIP_RAM.N_243 ));
    CascadeMux I__1708 (
            .O(N__7849),
            .I(N__7846));
    InMux I__1707 (
            .O(N__7846),
            .I(N__7838));
    InMux I__1706 (
            .O(N__7845),
            .I(N__7835));
    InMux I__1705 (
            .O(N__7844),
            .I(N__7832));
    InMux I__1704 (
            .O(N__7843),
            .I(N__7825));
    InMux I__1703 (
            .O(N__7842),
            .I(N__7825));
    InMux I__1702 (
            .O(N__7841),
            .I(N__7825));
    LocalMux I__1701 (
            .O(N__7838),
            .I(N__7812));
    LocalMux I__1700 (
            .O(N__7835),
            .I(N__7812));
    LocalMux I__1699 (
            .O(N__7832),
            .I(N__7812));
    LocalMux I__1698 (
            .O(N__7825),
            .I(N__7812));
    InMux I__1697 (
            .O(N__7824),
            .I(N__7809));
    InMux I__1696 (
            .O(N__7823),
            .I(N__7806));
    InMux I__1695 (
            .O(N__7822),
            .I(N__7803));
    InMux I__1694 (
            .O(N__7821),
            .I(N__7800));
    Span4Mux_v I__1693 (
            .O(N__7812),
            .I(N__7797));
    LocalMux I__1692 (
            .O(N__7809),
            .I(N__7788));
    LocalMux I__1691 (
            .O(N__7806),
            .I(N__7788));
    LocalMux I__1690 (
            .O(N__7803),
            .I(N__7788));
    LocalMux I__1689 (
            .O(N__7800),
            .I(N__7788));
    Sp12to4 I__1688 (
            .O(N__7797),
            .I(N__7785));
    Span12Mux_v I__1687 (
            .O(N__7788),
            .I(N__7782));
    Span12Mux_h I__1686 (
            .O(N__7785),
            .I(N__7779));
    Span12Mux_h I__1685 (
            .O(N__7782),
            .I(N__7776));
    Odrv12 I__1684 (
            .O(N__7779),
            .I(RESETn_c));
    Odrv12 I__1683 (
            .O(N__7776),
            .I(RESETn_c));
    IoInMux I__1682 (
            .O(N__7771),
            .I(N__7768));
    LocalMux I__1681 (
            .O(N__7768),
            .I(N__7765));
    Span12Mux_s1_v I__1680 (
            .O(N__7765),
            .I(N__7762));
    Odrv12 I__1679 (
            .O(N__7762),
            .I(RESETn_c_i));
    IoInMux I__1678 (
            .O(N__7759),
            .I(N__7756));
    LocalMux I__1677 (
            .O(N__7756),
            .I(N__7753));
    IoSpan4Mux I__1676 (
            .O(N__7753),
            .I(N__7750));
    IoSpan4Mux I__1675 (
            .O(N__7750),
            .I(N__7747));
    Span4Mux_s2_v I__1674 (
            .O(N__7747),
            .I(N__7743));
    InMux I__1673 (
            .O(N__7746),
            .I(N__7740));
    Span4Mux_v I__1672 (
            .O(N__7743),
            .I(N__7734));
    LocalMux I__1671 (
            .O(N__7740),
            .I(N__7734));
    CascadeMux I__1670 (
            .O(N__7739),
            .I(N__7729));
    Span4Mux_h I__1669 (
            .O(N__7734),
            .I(N__7725));
    InMux I__1668 (
            .O(N__7733),
            .I(N__7722));
    InMux I__1667 (
            .O(N__7732),
            .I(N__7719));
    InMux I__1666 (
            .O(N__7729),
            .I(N__7716));
    InMux I__1665 (
            .O(N__7728),
            .I(N__7713));
    Span4Mux_v I__1664 (
            .O(N__7725),
            .I(N__7710));
    LocalMux I__1663 (
            .O(N__7722),
            .I(N__7705));
    LocalMux I__1662 (
            .O(N__7719),
            .I(N__7705));
    LocalMux I__1661 (
            .O(N__7716),
            .I(N__7702));
    LocalMux I__1660 (
            .O(N__7713),
            .I(N__7699));
    Span4Mux_v I__1659 (
            .O(N__7710),
            .I(N__7692));
    Span4Mux_h I__1658 (
            .O(N__7705),
            .I(N__7692));
    Span4Mux_h I__1657 (
            .O(N__7702),
            .I(N__7692));
    Odrv12 I__1656 (
            .O(N__7699),
            .I(RAMENn_c));
    Odrv4 I__1655 (
            .O(N__7692),
            .I(RAMENn_c));
    InMux I__1654 (
            .O(N__7687),
            .I(N__7684));
    LocalMux I__1653 (
            .O(N__7684),
            .I(N__7680));
    InMux I__1652 (
            .O(N__7683),
            .I(N__7677));
    Span4Mux_v I__1651 (
            .O(N__7680),
            .I(N__7674));
    LocalMux I__1650 (
            .O(N__7677),
            .I(N__7671));
    Span4Mux_v I__1649 (
            .O(N__7674),
            .I(N__7667));
    Span4Mux_h I__1648 (
            .O(N__7671),
            .I(N__7664));
    InMux I__1647 (
            .O(N__7670),
            .I(N__7661));
    Odrv4 I__1646 (
            .O(N__7667),
            .I(REG_CYCLEm));
    Odrv4 I__1645 (
            .O(N__7664),
            .I(REG_CYCLEm));
    LocalMux I__1644 (
            .O(N__7661),
            .I(REG_CYCLEm));
    IoInMux I__1643 (
            .O(N__7654),
            .I(N__7651));
    LocalMux I__1642 (
            .O(N__7651),
            .I(N__7648));
    IoSpan4Mux I__1641 (
            .O(N__7648),
            .I(N__7645));
    Sp12to4 I__1640 (
            .O(N__7645),
            .I(N__7642));
    Span12Mux_s6_v I__1639 (
            .O(N__7642),
            .I(N__7639));
    Span12Mux_h I__1638 (
            .O(N__7639),
            .I(N__7636));
    Odrv12 I__1637 (
            .O(N__7636),
            .I(DRDENn_c));
    InMux I__1636 (
            .O(N__7633),
            .I(N__7630));
    LocalMux I__1635 (
            .O(N__7630),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__1634 (
            .O(N__7627),
            .I(N__7624));
    LocalMux I__1633 (
            .O(N__7624),
            .I(N__7621));
    Span12Mux_s0_v I__1632 (
            .O(N__7621),
            .I(N__7618));
    Span12Mux_v I__1631 (
            .O(N__7618),
            .I(N__7615));
    Odrv12 I__1630 (
            .O(N__7615),
            .I(CMA_c_0));
    CascadeMux I__1629 (
            .O(N__7612),
            .I(N__7609));
    InMux I__1628 (
            .O(N__7609),
            .I(N__7606));
    LocalMux I__1627 (
            .O(N__7606),
            .I(N__7603));
    Odrv12 I__1626 (
            .O(N__7603),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__1625 (
            .O(N__7600),
            .I(N__7597));
    LocalMux I__1624 (
            .O(N__7597),
            .I(N__7594));
    Odrv4 I__1623 (
            .O(N__7594),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__1622 (
            .O(N__7591),
            .I(N__7587));
    InMux I__1621 (
            .O(N__7590),
            .I(N__7584));
    LocalMux I__1620 (
            .O(N__7587),
            .I(N__7579));
    LocalMux I__1619 (
            .O(N__7584),
            .I(N__7579));
    Sp12to4 I__1618 (
            .O(N__7579),
            .I(N__7576));
    Span12Mux_v I__1617 (
            .O(N__7576),
            .I(N__7573));
    Span12Mux_h I__1616 (
            .O(N__7573),
            .I(N__7570));
    Odrv12 I__1615 (
            .O(N__7570),
            .I(DRA_c_2));
    InMux I__1614 (
            .O(N__7567),
            .I(N__7564));
    LocalMux I__1613 (
            .O(N__7564),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    CascadeMux I__1612 (
            .O(N__7561),
            .I(N__7558));
    InMux I__1611 (
            .O(N__7558),
            .I(N__7555));
    LocalMux I__1610 (
            .O(N__7555),
            .I(N__7552));
    Odrv4 I__1609 (
            .O(N__7552),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1608 (
            .O(N__7549),
            .I(N__7546));
    LocalMux I__1607 (
            .O(N__7546),
            .I(N__7543));
    Span4Mux_h I__1606 (
            .O(N__7543),
            .I(N__7540));
    Odrv4 I__1605 (
            .O(N__7540),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1604 (
            .O(N__7537),
            .I(N__7531));
    InMux I__1603 (
            .O(N__7536),
            .I(N__7528));
    InMux I__1602 (
            .O(N__7535),
            .I(N__7517));
    InMux I__1601 (
            .O(N__7534),
            .I(N__7517));
    LocalMux I__1600 (
            .O(N__7531),
            .I(N__7513));
    LocalMux I__1599 (
            .O(N__7528),
            .I(N__7510));
    InMux I__1598 (
            .O(N__7527),
            .I(N__7506));
    InMux I__1597 (
            .O(N__7526),
            .I(N__7500));
    InMux I__1596 (
            .O(N__7525),
            .I(N__7493));
    InMux I__1595 (
            .O(N__7524),
            .I(N__7493));
    InMux I__1594 (
            .O(N__7523),
            .I(N__7493));
    InMux I__1593 (
            .O(N__7522),
            .I(N__7490));
    LocalMux I__1592 (
            .O(N__7517),
            .I(N__7487));
    InMux I__1591 (
            .O(N__7516),
            .I(N__7484));
    Span4Mux_v I__1590 (
            .O(N__7513),
            .I(N__7479));
    Span4Mux_h I__1589 (
            .O(N__7510),
            .I(N__7479));
    InMux I__1588 (
            .O(N__7509),
            .I(N__7476));
    LocalMux I__1587 (
            .O(N__7506),
            .I(N__7473));
    InMux I__1586 (
            .O(N__7505),
            .I(N__7468));
    InMux I__1585 (
            .O(N__7504),
            .I(N__7468));
    InMux I__1584 (
            .O(N__7503),
            .I(N__7465));
    LocalMux I__1583 (
            .O(N__7500),
            .I(N__7460));
    LocalMux I__1582 (
            .O(N__7493),
            .I(N__7460));
    LocalMux I__1581 (
            .O(N__7490),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1580 (
            .O(N__7487),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1579 (
            .O(N__7484),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1578 (
            .O(N__7479),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1577 (
            .O(N__7476),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1576 (
            .O(N__7473),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1575 (
            .O(N__7468),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1574 (
            .O(N__7465),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1573 (
            .O(N__7460),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1572 (
            .O(N__7441),
            .I(N__7437));
    InMux I__1571 (
            .O(N__7440),
            .I(N__7434));
    LocalMux I__1570 (
            .O(N__7437),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1Z0Z_1 ));
    LocalMux I__1569 (
            .O(N__7434),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1Z0Z_1 ));
    InMux I__1568 (
            .O(N__7429),
            .I(N__7426));
    LocalMux I__1567 (
            .O(N__7426),
            .I(N__7423));
    Odrv12 I__1566 (
            .O(N__7423),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_0 ));
    InMux I__1565 (
            .O(N__7420),
            .I(N__7416));
    InMux I__1564 (
            .O(N__7419),
            .I(N__7413));
    LocalMux I__1563 (
            .O(N__7416),
            .I(CPU_TACKm));
    LocalMux I__1562 (
            .O(N__7413),
            .I(CPU_TACKm));
    InMux I__1561 (
            .O(N__7408),
            .I(N__7404));
    CascadeMux I__1560 (
            .O(N__7407),
            .I(N__7400));
    LocalMux I__1559 (
            .O(N__7404),
            .I(N__7397));
    InMux I__1558 (
            .O(N__7403),
            .I(N__7394));
    InMux I__1557 (
            .O(N__7400),
            .I(N__7391));
    Span4Mux_v I__1556 (
            .O(N__7397),
            .I(N__7388));
    LocalMux I__1555 (
            .O(N__7394),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1554 (
            .O(N__7391),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    Odrv4 I__1553 (
            .O(N__7388),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    CascadeMux I__1552 (
            .O(N__7381),
            .I(N__7378));
    InMux I__1551 (
            .O(N__7378),
            .I(N__7375));
    LocalMux I__1550 (
            .O(N__7375),
            .I(N__7370));
    InMux I__1549 (
            .O(N__7374),
            .I(N__7366));
    InMux I__1548 (
            .O(N__7373),
            .I(N__7363));
    Span4Mux_h I__1547 (
            .O(N__7370),
            .I(N__7360));
    InMux I__1546 (
            .O(N__7369),
            .I(N__7357));
    LocalMux I__1545 (
            .O(N__7366),
            .I(\U712_REG_SM.N_187 ));
    LocalMux I__1544 (
            .O(N__7363),
            .I(\U712_REG_SM.N_187 ));
    Odrv4 I__1543 (
            .O(N__7360),
            .I(\U712_REG_SM.N_187 ));
    LocalMux I__1542 (
            .O(N__7357),
            .I(\U712_REG_SM.N_187 ));
    CascadeMux I__1541 (
            .O(N__7348),
            .I(N__7345));
    InMux I__1540 (
            .O(N__7345),
            .I(N__7341));
    InMux I__1539 (
            .O(N__7344),
            .I(N__7338));
    LocalMux I__1538 (
            .O(N__7341),
            .I(N__7333));
    LocalMux I__1537 (
            .O(N__7338),
            .I(N__7330));
    InMux I__1536 (
            .O(N__7337),
            .I(N__7325));
    InMux I__1535 (
            .O(N__7336),
            .I(N__7325));
    Span4Mux_h I__1534 (
            .O(N__7333),
            .I(N__7322));
    Span4Mux_v I__1533 (
            .O(N__7330),
            .I(N__7319));
    LocalMux I__1532 (
            .O(N__7325),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    Odrv4 I__1531 (
            .O(N__7322),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    Odrv4 I__1530 (
            .O(N__7319),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    InMux I__1529 (
            .O(N__7312),
            .I(N__7306));
    InMux I__1528 (
            .O(N__7311),
            .I(N__7306));
    LocalMux I__1527 (
            .O(N__7306),
            .I(REG_TACK));
    InMux I__1526 (
            .O(N__7303),
            .I(N__7300));
    LocalMux I__1525 (
            .O(N__7300),
            .I(N__7297));
    Odrv4 I__1524 (
            .O(N__7297),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_0_a3_0 ));
    InMux I__1523 (
            .O(N__7294),
            .I(N__7291));
    LocalMux I__1522 (
            .O(N__7291),
            .I(N__7288));
    Span4Mux_v I__1521 (
            .O(N__7288),
            .I(N__7285));
    Odrv4 I__1520 (
            .O(N__7285),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    InMux I__1519 (
            .O(N__7282),
            .I(N__7279));
    LocalMux I__1518 (
            .O(N__7279),
            .I(N__7276));
    Odrv4 I__1517 (
            .O(N__7276),
            .I(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a3_0_a3_0 ));
    InMux I__1516 (
            .O(N__7273),
            .I(N__7259));
    InMux I__1515 (
            .O(N__7272),
            .I(N__7259));
    InMux I__1514 (
            .O(N__7271),
            .I(N__7259));
    InMux I__1513 (
            .O(N__7270),
            .I(N__7254));
    InMux I__1512 (
            .O(N__7269),
            .I(N__7254));
    InMux I__1511 (
            .O(N__7268),
            .I(N__7247));
    InMux I__1510 (
            .O(N__7267),
            .I(N__7247));
    InMux I__1509 (
            .O(N__7266),
            .I(N__7247));
    LocalMux I__1508 (
            .O(N__7259),
            .I(\U712_CHIP_RAM.N_96 ));
    LocalMux I__1507 (
            .O(N__7254),
            .I(\U712_CHIP_RAM.N_96 ));
    LocalMux I__1506 (
            .O(N__7247),
            .I(\U712_CHIP_RAM.N_96 ));
    CascadeMux I__1505 (
            .O(N__7240),
            .I(N__7235));
    CascadeMux I__1504 (
            .O(N__7239),
            .I(N__7232));
    InMux I__1503 (
            .O(N__7238),
            .I(N__7229));
    InMux I__1502 (
            .O(N__7235),
            .I(N__7224));
    InMux I__1501 (
            .O(N__7232),
            .I(N__7224));
    LocalMux I__1500 (
            .O(N__7229),
            .I(N__7221));
    LocalMux I__1499 (
            .O(N__7224),
            .I(N__7213));
    Span4Mux_v I__1498 (
            .O(N__7221),
            .I(N__7213));
    InMux I__1497 (
            .O(N__7220),
            .I(N__7210));
    InMux I__1496 (
            .O(N__7219),
            .I(N__7207));
    InMux I__1495 (
            .O(N__7218),
            .I(N__7204));
    Odrv4 I__1494 (
            .O(N__7213),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER16 ));
    LocalMux I__1493 (
            .O(N__7210),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER16 ));
    LocalMux I__1492 (
            .O(N__7207),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER16 ));
    LocalMux I__1491 (
            .O(N__7204),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER16 ));
    InMux I__1490 (
            .O(N__7195),
            .I(N__7192));
    LocalMux I__1489 (
            .O(N__7192),
            .I(N__7189));
    Span4Mux_h I__1488 (
            .O(N__7189),
            .I(N__7186));
    Odrv4 I__1487 (
            .O(N__7186),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    CEMux I__1486 (
            .O(N__7183),
            .I(N__7179));
    CEMux I__1485 (
            .O(N__7182),
            .I(N__7176));
    LocalMux I__1484 (
            .O(N__7179),
            .I(N__7173));
    LocalMux I__1483 (
            .O(N__7176),
            .I(N__7170));
    Span4Mux_h I__1482 (
            .O(N__7173),
            .I(N__7167));
    Odrv12 I__1481 (
            .O(N__7170),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv4 I__1480 (
            .O(N__7167),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    CascadeMux I__1479 (
            .O(N__7162),
            .I(N__7158));
    CascadeMux I__1478 (
            .O(N__7161),
            .I(N__7152));
    InMux I__1477 (
            .O(N__7158),
            .I(N__7146));
    InMux I__1476 (
            .O(N__7157),
            .I(N__7146));
    InMux I__1475 (
            .O(N__7156),
            .I(N__7141));
    InMux I__1474 (
            .O(N__7155),
            .I(N__7141));
    InMux I__1473 (
            .O(N__7152),
            .I(N__7125));
    InMux I__1472 (
            .O(N__7151),
            .I(N__7125));
    LocalMux I__1471 (
            .O(N__7146),
            .I(N__7122));
    LocalMux I__1470 (
            .O(N__7141),
            .I(N__7119));
    InMux I__1469 (
            .O(N__7140),
            .I(N__7110));
    InMux I__1468 (
            .O(N__7139),
            .I(N__7110));
    InMux I__1467 (
            .O(N__7138),
            .I(N__7110));
    InMux I__1466 (
            .O(N__7137),
            .I(N__7110));
    InMux I__1465 (
            .O(N__7136),
            .I(N__7107));
    InMux I__1464 (
            .O(N__7135),
            .I(N__7104));
    InMux I__1463 (
            .O(N__7134),
            .I(N__7099));
    InMux I__1462 (
            .O(N__7133),
            .I(N__7099));
    InMux I__1461 (
            .O(N__7132),
            .I(N__7096));
    InMux I__1460 (
            .O(N__7131),
            .I(N__7091));
    InMux I__1459 (
            .O(N__7130),
            .I(N__7091));
    LocalMux I__1458 (
            .O(N__7125),
            .I(N__7086));
    Span4Mux_h I__1457 (
            .O(N__7122),
            .I(N__7086));
    Span4Mux_h I__1456 (
            .O(N__7119),
            .I(N__7083));
    LocalMux I__1455 (
            .O(N__7110),
            .I(N__7080));
    LocalMux I__1454 (
            .O(N__7107),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1453 (
            .O(N__7104),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1452 (
            .O(N__7099),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1451 (
            .O(N__7096),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1450 (
            .O(N__7091),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1449 (
            .O(N__7086),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1448 (
            .O(N__7083),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv12 I__1447 (
            .O(N__7080),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__1446 (
            .O(N__7063),
            .I(N__7060));
    LocalMux I__1445 (
            .O(N__7060),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_0_a3_0 ));
    InMux I__1444 (
            .O(N__7057),
            .I(N__7054));
    LocalMux I__1443 (
            .O(N__7054),
            .I(\U712_CYCLE_TERM.N_214_i_0_en ));
    InMux I__1442 (
            .O(N__7051),
            .I(N__7034));
    InMux I__1441 (
            .O(N__7050),
            .I(N__7034));
    InMux I__1440 (
            .O(N__7049),
            .I(N__7031));
    InMux I__1439 (
            .O(N__7048),
            .I(N__7025));
    InMux I__1438 (
            .O(N__7047),
            .I(N__7022));
    InMux I__1437 (
            .O(N__7046),
            .I(N__7013));
    InMux I__1436 (
            .O(N__7045),
            .I(N__7013));
    InMux I__1435 (
            .O(N__7044),
            .I(N__7013));
    InMux I__1434 (
            .O(N__7043),
            .I(N__7013));
    InMux I__1433 (
            .O(N__7042),
            .I(N__7008));
    InMux I__1432 (
            .O(N__7041),
            .I(N__7008));
    CascadeMux I__1431 (
            .O(N__7040),
            .I(N__7004));
    CascadeMux I__1430 (
            .O(N__7039),
            .I(N__6995));
    LocalMux I__1429 (
            .O(N__7034),
            .I(N__6988));
    LocalMux I__1428 (
            .O(N__7031),
            .I(N__6985));
    InMux I__1427 (
            .O(N__7030),
            .I(N__6978));
    InMux I__1426 (
            .O(N__7029),
            .I(N__6978));
    InMux I__1425 (
            .O(N__7028),
            .I(N__6978));
    LocalMux I__1424 (
            .O(N__7025),
            .I(N__6975));
    LocalMux I__1423 (
            .O(N__7022),
            .I(N__6968));
    LocalMux I__1422 (
            .O(N__7013),
            .I(N__6968));
    LocalMux I__1421 (
            .O(N__7008),
            .I(N__6968));
    InMux I__1420 (
            .O(N__7007),
            .I(N__6965));
    InMux I__1419 (
            .O(N__7004),
            .I(N__6962));
    InMux I__1418 (
            .O(N__7003),
            .I(N__6959));
    InMux I__1417 (
            .O(N__7002),
            .I(N__6954));
    InMux I__1416 (
            .O(N__7001),
            .I(N__6954));
    InMux I__1415 (
            .O(N__7000),
            .I(N__6949));
    InMux I__1414 (
            .O(N__6999),
            .I(N__6949));
    InMux I__1413 (
            .O(N__6998),
            .I(N__6944));
    InMux I__1412 (
            .O(N__6995),
            .I(N__6944));
    InMux I__1411 (
            .O(N__6994),
            .I(N__6941));
    InMux I__1410 (
            .O(N__6993),
            .I(N__6934));
    InMux I__1409 (
            .O(N__6992),
            .I(N__6934));
    InMux I__1408 (
            .O(N__6991),
            .I(N__6934));
    Span4Mux_v I__1407 (
            .O(N__6988),
            .I(N__6927));
    Span4Mux_v I__1406 (
            .O(N__6985),
            .I(N__6927));
    LocalMux I__1405 (
            .O(N__6978),
            .I(N__6927));
    Span4Mux_h I__1404 (
            .O(N__6975),
            .I(N__6922));
    Span4Mux_h I__1403 (
            .O(N__6968),
            .I(N__6922));
    LocalMux I__1402 (
            .O(N__6965),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1401 (
            .O(N__6962),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1400 (
            .O(N__6959),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1399 (
            .O(N__6954),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1398 (
            .O(N__6949),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1397 (
            .O(N__6944),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1396 (
            .O(N__6941),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1395 (
            .O(N__6934),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1394 (
            .O(N__6927),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1393 (
            .O(N__6922),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    CascadeMux I__1392 (
            .O(N__6901),
            .I(N__6894));
    CascadeMux I__1391 (
            .O(N__6900),
            .I(N__6890));
    CascadeMux I__1390 (
            .O(N__6899),
            .I(N__6886));
    CascadeMux I__1389 (
            .O(N__6898),
            .I(N__6882));
    CascadeMux I__1388 (
            .O(N__6897),
            .I(N__6876));
    InMux I__1387 (
            .O(N__6894),
            .I(N__6873));
    InMux I__1386 (
            .O(N__6893),
            .I(N__6870));
    InMux I__1385 (
            .O(N__6890),
            .I(N__6866));
    InMux I__1384 (
            .O(N__6889),
            .I(N__6861));
    InMux I__1383 (
            .O(N__6886),
            .I(N__6861));
    InMux I__1382 (
            .O(N__6885),
            .I(N__6856));
    InMux I__1381 (
            .O(N__6882),
            .I(N__6856));
    InMux I__1380 (
            .O(N__6881),
            .I(N__6849));
    InMux I__1379 (
            .O(N__6880),
            .I(N__6849));
    InMux I__1378 (
            .O(N__6879),
            .I(N__6849));
    InMux I__1377 (
            .O(N__6876),
            .I(N__6846));
    LocalMux I__1376 (
            .O(N__6873),
            .I(N__6839));
    LocalMux I__1375 (
            .O(N__6870),
            .I(N__6839));
    InMux I__1374 (
            .O(N__6869),
            .I(N__6836));
    LocalMux I__1373 (
            .O(N__6866),
            .I(N__6829));
    LocalMux I__1372 (
            .O(N__6861),
            .I(N__6829));
    LocalMux I__1371 (
            .O(N__6856),
            .I(N__6829));
    LocalMux I__1370 (
            .O(N__6849),
            .I(N__6823));
    LocalMux I__1369 (
            .O(N__6846),
            .I(N__6823));
    InMux I__1368 (
            .O(N__6845),
            .I(N__6820));
    InMux I__1367 (
            .O(N__6844),
            .I(N__6817));
    Span4Mux_v I__1366 (
            .O(N__6839),
            .I(N__6810));
    LocalMux I__1365 (
            .O(N__6836),
            .I(N__6810));
    Span4Mux_v I__1364 (
            .O(N__6829),
            .I(N__6810));
    InMux I__1363 (
            .O(N__6828),
            .I(N__6807));
    Odrv4 I__1362 (
            .O(N__6823),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1361 (
            .O(N__6820),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1360 (
            .O(N__6817),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1359 (
            .O(N__6810),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1358 (
            .O(N__6807),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    IoInMux I__1357 (
            .O(N__6796),
            .I(N__6793));
    LocalMux I__1356 (
            .O(N__6793),
            .I(N__6790));
    Span4Mux_s3_h I__1355 (
            .O(N__6790),
            .I(N__6787));
    Sp12to4 I__1354 (
            .O(N__6787),
            .I(N__6784));
    Span12Mux_v I__1353 (
            .O(N__6784),
            .I(N__6781));
    Span12Mux_h I__1352 (
            .O(N__6781),
            .I(N__6778));
    Odrv12 I__1351 (
            .O(N__6778),
            .I(CMA_c_5));
    InMux I__1350 (
            .O(N__6775),
            .I(N__6772));
    LocalMux I__1349 (
            .O(N__6772),
            .I(N__6769));
    Span4Mux_v I__1348 (
            .O(N__6769),
            .I(N__6766));
    Sp12to4 I__1347 (
            .O(N__6766),
            .I(N__6763));
    Span12Mux_h I__1346 (
            .O(N__6763),
            .I(N__6760));
    Odrv12 I__1345 (
            .O(N__6760),
            .I(A_c_7));
    CascadeMux I__1344 (
            .O(N__6757),
            .I(\U712_CHIP_RAM.N_316_cascade_ ));
    InMux I__1343 (
            .O(N__6754),
            .I(N__6751));
    LocalMux I__1342 (
            .O(N__6751),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    InMux I__1341 (
            .O(N__6748),
            .I(N__6745));
    LocalMux I__1340 (
            .O(N__6745),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    InMux I__1339 (
            .O(N__6742),
            .I(N__6736));
    InMux I__1338 (
            .O(N__6741),
            .I(N__6736));
    LocalMux I__1337 (
            .O(N__6736),
            .I(N__6733));
    Span4Mux_h I__1336 (
            .O(N__6733),
            .I(N__6728));
    InMux I__1335 (
            .O(N__6732),
            .I(N__6723));
    InMux I__1334 (
            .O(N__6731),
            .I(N__6723));
    Odrv4 I__1333 (
            .O(N__6728),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1332 (
            .O(N__6723),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    CascadeMux I__1331 (
            .O(N__6718),
            .I(N__6715));
    InMux I__1330 (
            .O(N__6715),
            .I(N__6709));
    InMux I__1329 (
            .O(N__6714),
            .I(N__6709));
    LocalMux I__1328 (
            .O(N__6709),
            .I(N__6706));
    Span4Mux_h I__1327 (
            .O(N__6706),
            .I(N__6703));
    Sp12to4 I__1326 (
            .O(N__6703),
            .I(N__6700));
    Span12Mux_v I__1325 (
            .O(N__6700),
            .I(N__6697));
    Span12Mux_h I__1324 (
            .O(N__6697),
            .I(N__6694));
    Odrv12 I__1323 (
            .O(N__6694),
            .I(A_c_14));
    InMux I__1322 (
            .O(N__6691),
            .I(N__6688));
    LocalMux I__1321 (
            .O(N__6688),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__1320 (
            .O(N__6685),
            .I(N__6682));
    LocalMux I__1319 (
            .O(N__6682),
            .I(N__6679));
    Span4Mux_h I__1318 (
            .O(N__6679),
            .I(N__6670));
    InMux I__1317 (
            .O(N__6678),
            .I(N__6667));
    InMux I__1316 (
            .O(N__6677),
            .I(N__6662));
    InMux I__1315 (
            .O(N__6676),
            .I(N__6662));
    InMux I__1314 (
            .O(N__6675),
            .I(N__6659));
    InMux I__1313 (
            .O(N__6674),
            .I(N__6656));
    InMux I__1312 (
            .O(N__6673),
            .I(N__6653));
    Odrv4 I__1311 (
            .O(N__6670),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1310 (
            .O(N__6667),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1309 (
            .O(N__6662),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1308 (
            .O(N__6659),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1307 (
            .O(N__6656),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1306 (
            .O(N__6653),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    CEMux I__1305 (
            .O(N__6640),
            .I(N__6637));
    LocalMux I__1304 (
            .O(N__6637),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_3_0_0 ));
    InMux I__1303 (
            .O(N__6634),
            .I(N__6631));
    LocalMux I__1302 (
            .O(N__6631),
            .I(N__6627));
    InMux I__1301 (
            .O(N__6630),
            .I(N__6623));
    Span4Mux_v I__1300 (
            .O(N__6627),
            .I(N__6618));
    InMux I__1299 (
            .O(N__6626),
            .I(N__6615));
    LocalMux I__1298 (
            .O(N__6623),
            .I(N__6612));
    InMux I__1297 (
            .O(N__6622),
            .I(N__6609));
    InMux I__1296 (
            .O(N__6621),
            .I(N__6606));
    Odrv4 I__1295 (
            .O(N__6618),
            .I(\U712_CHIP_RAM.N_180 ));
    LocalMux I__1294 (
            .O(N__6615),
            .I(\U712_CHIP_RAM.N_180 ));
    Odrv4 I__1293 (
            .O(N__6612),
            .I(\U712_CHIP_RAM.N_180 ));
    LocalMux I__1292 (
            .O(N__6609),
            .I(\U712_CHIP_RAM.N_180 ));
    LocalMux I__1291 (
            .O(N__6606),
            .I(\U712_CHIP_RAM.N_180 ));
    InMux I__1290 (
            .O(N__6595),
            .I(N__6592));
    LocalMux I__1289 (
            .O(N__6592),
            .I(N__6589));
    Span4Mux_v I__1288 (
            .O(N__6589),
            .I(N__6586));
    Odrv4 I__1287 (
            .O(N__6586),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a3_2_1_0 ));
    InMux I__1286 (
            .O(N__6583),
            .I(N__6578));
    CascadeMux I__1285 (
            .O(N__6582),
            .I(N__6575));
    InMux I__1284 (
            .O(N__6581),
            .I(N__6572));
    LocalMux I__1283 (
            .O(N__6578),
            .I(N__6569));
    InMux I__1282 (
            .O(N__6575),
            .I(N__6566));
    LocalMux I__1281 (
            .O(N__6572),
            .I(\U712_CHIP_RAM.N_254_2 ));
    Odrv4 I__1280 (
            .O(N__6569),
            .I(\U712_CHIP_RAM.N_254_2 ));
    LocalMux I__1279 (
            .O(N__6566),
            .I(\U712_CHIP_RAM.N_254_2 ));
    InMux I__1278 (
            .O(N__6559),
            .I(N__6556));
    LocalMux I__1277 (
            .O(N__6556),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__1276 (
            .O(N__6553),
            .I(N__6550));
    LocalMux I__1275 (
            .O(N__6550),
            .I(N__6547));
    IoSpan4Mux I__1274 (
            .O(N__6547),
            .I(N__6544));
    Span4Mux_s2_h I__1273 (
            .O(N__6544),
            .I(N__6541));
    Sp12to4 I__1272 (
            .O(N__6541),
            .I(N__6538));
    Span12Mux_h I__1271 (
            .O(N__6538),
            .I(N__6535));
    Odrv12 I__1270 (
            .O(N__6535),
            .I(CMA_c_7));
    InMux I__1269 (
            .O(N__6532),
            .I(N__6529));
    LocalMux I__1268 (
            .O(N__6529),
            .I(N__6526));
    Span12Mux_v I__1267 (
            .O(N__6526),
            .I(N__6523));
    Span12Mux_h I__1266 (
            .O(N__6523),
            .I(N__6520));
    Odrv12 I__1265 (
            .O(N__6520),
            .I(A_c_15));
    InMux I__1264 (
            .O(N__6517),
            .I(N__6514));
    LocalMux I__1263 (
            .O(N__6514),
            .I(N__6511));
    Span4Mux_v I__1262 (
            .O(N__6511),
            .I(N__6508));
    Sp12to4 I__1261 (
            .O(N__6508),
            .I(N__6505));
    Span12Mux_h I__1260 (
            .O(N__6505),
            .I(N__6502));
    Odrv12 I__1259 (
            .O(N__6502),
            .I(A_c_8));
    CascadeMux I__1258 (
            .O(N__6499),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ));
    InMux I__1257 (
            .O(N__6496),
            .I(N__6493));
    LocalMux I__1256 (
            .O(N__6493),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    InMux I__1255 (
            .O(N__6490),
            .I(N__6487));
    LocalMux I__1254 (
            .O(N__6487),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    InMux I__1253 (
            .O(N__6484),
            .I(N__6481));
    LocalMux I__1252 (
            .O(N__6481),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ));
    InMux I__1251 (
            .O(N__6478),
            .I(N__6475));
    LocalMux I__1250 (
            .O(N__6475),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    CascadeMux I__1249 (
            .O(N__6472),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ));
    InMux I__1248 (
            .O(N__6469),
            .I(N__6466));
    LocalMux I__1247 (
            .O(N__6466),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    IoInMux I__1246 (
            .O(N__6463),
            .I(N__6460));
    LocalMux I__1245 (
            .O(N__6460),
            .I(N__6457));
    Span12Mux_s7_v I__1244 (
            .O(N__6457),
            .I(N__6454));
    Odrv12 I__1243 (
            .O(N__6454),
            .I(CMA_c_1));
    CEMux I__1242 (
            .O(N__6451),
            .I(N__6448));
    LocalMux I__1241 (
            .O(N__6448),
            .I(N__6445));
    Odrv4 I__1240 (
            .O(N__6445),
            .I(\U712_CYCLE_TERM.N_214_i_0_en_0 ));
    InMux I__1239 (
            .O(N__6442),
            .I(N__6439));
    LocalMux I__1238 (
            .O(N__6439),
            .I(N__6436));
    Odrv4 I__1237 (
            .O(N__6436),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_1 ));
    InMux I__1236 (
            .O(N__6433),
            .I(N__6430));
    LocalMux I__1235 (
            .O(N__6430),
            .I(N__6427));
    Odrv4 I__1234 (
            .O(N__6427),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_3 ));
    IoInMux I__1233 (
            .O(N__6424),
            .I(N__6421));
    LocalMux I__1232 (
            .O(N__6421),
            .I(N__6418));
    Span4Mux_s2_v I__1231 (
            .O(N__6418),
            .I(N__6415));
    Span4Mux_v I__1230 (
            .O(N__6415),
            .I(N__6412));
    Odrv4 I__1229 (
            .O(N__6412),
            .I(CONSTANT_ONE_NET));
    IoInMux I__1228 (
            .O(N__6409),
            .I(N__6406));
    LocalMux I__1227 (
            .O(N__6406),
            .I(N__6403));
    Span4Mux_s2_v I__1226 (
            .O(N__6403),
            .I(N__6400));
    Span4Mux_v I__1225 (
            .O(N__6400),
            .I(N__6397));
    Span4Mux_v I__1224 (
            .O(N__6397),
            .I(N__6394));
    Span4Mux_h I__1223 (
            .O(N__6394),
            .I(N__6391));
    Odrv4 I__1222 (
            .O(N__6391),
            .I(CRCSn_c));
    IoInMux I__1221 (
            .O(N__6388),
            .I(N__6385));
    LocalMux I__1220 (
            .O(N__6385),
            .I(N__6382));
    Span4Mux_s0_h I__1219 (
            .O(N__6382),
            .I(N__6379));
    Span4Mux_h I__1218 (
            .O(N__6379),
            .I(N__6376));
    Sp12to4 I__1217 (
            .O(N__6376),
            .I(N__6373));
    Span12Mux_s9_v I__1216 (
            .O(N__6373),
            .I(N__6370));
    Span12Mux_h I__1215 (
            .O(N__6370),
            .I(N__6367));
    Odrv12 I__1214 (
            .O(N__6367),
            .I(WEn_c));
    InMux I__1213 (
            .O(N__6364),
            .I(N__6361));
    LocalMux I__1212 (
            .O(N__6361),
            .I(N__6358));
    Span12Mux_v I__1211 (
            .O(N__6358),
            .I(N__6355));
    Span12Mux_h I__1210 (
            .O(N__6355),
            .I(N__6352));
    Odrv12 I__1209 (
            .O(N__6352),
            .I(A_c_19));
    CascadeMux I__1208 (
            .O(N__6349),
            .I(N__6346));
    InMux I__1207 (
            .O(N__6346),
            .I(N__6343));
    LocalMux I__1206 (
            .O(N__6343),
            .I(N__6340));
    Span12Mux_v I__1205 (
            .O(N__6340),
            .I(N__6337));
    Span12Mux_h I__1204 (
            .O(N__6337),
            .I(N__6334));
    Odrv12 I__1203 (
            .O(N__6334),
            .I(RAS0n_c));
    IoInMux I__1202 (
            .O(N__6331),
            .I(N__6328));
    LocalMux I__1201 (
            .O(N__6328),
            .I(N__6325));
    IoSpan4Mux I__1200 (
            .O(N__6325),
            .I(N__6322));
    Span4Mux_s2_h I__1199 (
            .O(N__6322),
            .I(N__6319));
    Sp12to4 I__1198 (
            .O(N__6319),
            .I(N__6316));
    Span12Mux_h I__1197 (
            .O(N__6316),
            .I(N__6313));
    Odrv12 I__1196 (
            .O(N__6313),
            .I(CMA_c_9));
    InMux I__1195 (
            .O(N__6310),
            .I(N__6307));
    LocalMux I__1194 (
            .O(N__6307),
            .I(N__6304));
    Span12Mux_v I__1193 (
            .O(N__6304),
            .I(N__6301));
    Span12Mux_h I__1192 (
            .O(N__6301),
            .I(N__6298));
    Odrv12 I__1191 (
            .O(N__6298),
            .I(A_c_17));
    IoInMux I__1190 (
            .O(N__6295),
            .I(N__6292));
    LocalMux I__1189 (
            .O(N__6292),
            .I(N__6289));
    IoSpan4Mux I__1188 (
            .O(N__6289),
            .I(N__6286));
    Span4Mux_s3_h I__1187 (
            .O(N__6286),
            .I(N__6283));
    Span4Mux_v I__1186 (
            .O(N__6283),
            .I(N__6280));
    Span4Mux_h I__1185 (
            .O(N__6280),
            .I(N__6277));
    Sp12to4 I__1184 (
            .O(N__6277),
            .I(N__6274));
    Odrv12 I__1183 (
            .O(N__6274),
            .I(CMA_c_8));
    IoInMux I__1182 (
            .O(N__6271),
            .I(N__6268));
    LocalMux I__1181 (
            .O(N__6268),
            .I(N__6265));
    IoSpan4Mux I__1180 (
            .O(N__6265),
            .I(N__6262));
    Span4Mux_s3_h I__1179 (
            .O(N__6262),
            .I(N__6259));
    Sp12to4 I__1178 (
            .O(N__6259),
            .I(N__6256));
    Span12Mux_s8_h I__1177 (
            .O(N__6256),
            .I(N__6253));
    Span12Mux_v I__1176 (
            .O(N__6253),
            .I(N__6250));
    Odrv12 I__1175 (
            .O(N__6250),
            .I(CMA_c_6));
    InMux I__1174 (
            .O(N__6247),
            .I(N__6242));
    InMux I__1173 (
            .O(N__6246),
            .I(N__6239));
    CascadeMux I__1172 (
            .O(N__6245),
            .I(N__6236));
    LocalMux I__1171 (
            .O(N__6242),
            .I(N__6230));
    LocalMux I__1170 (
            .O(N__6239),
            .I(N__6230));
    InMux I__1169 (
            .O(N__6236),
            .I(N__6227));
    InMux I__1168 (
            .O(N__6235),
            .I(N__6224));
    Span4Mux_v I__1167 (
            .O(N__6230),
            .I(N__6221));
    LocalMux I__1166 (
            .O(N__6227),
            .I(N__6216));
    LocalMux I__1165 (
            .O(N__6224),
            .I(N__6216));
    Odrv4 I__1164 (
            .O(N__6221),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1163 (
            .O(N__6216),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    InMux I__1162 (
            .O(N__6211),
            .I(N__6207));
    InMux I__1161 (
            .O(N__6210),
            .I(N__6204));
    LocalMux I__1160 (
            .O(N__6207),
            .I(N__6200));
    LocalMux I__1159 (
            .O(N__6204),
            .I(N__6197));
    CascadeMux I__1158 (
            .O(N__6203),
            .I(N__6193));
    Span4Mux_v I__1157 (
            .O(N__6200),
            .I(N__6187));
    Span4Mux_h I__1156 (
            .O(N__6197),
            .I(N__6187));
    InMux I__1155 (
            .O(N__6196),
            .I(N__6182));
    InMux I__1154 (
            .O(N__6193),
            .I(N__6179));
    InMux I__1153 (
            .O(N__6192),
            .I(N__6176));
    Span4Mux_v I__1152 (
            .O(N__6187),
            .I(N__6173));
    InMux I__1151 (
            .O(N__6186),
            .I(N__6168));
    InMux I__1150 (
            .O(N__6185),
            .I(N__6168));
    LocalMux I__1149 (
            .O(N__6182),
            .I(N__6165));
    LocalMux I__1148 (
            .O(N__6179),
            .I(N__6162));
    LocalMux I__1147 (
            .O(N__6176),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1146 (
            .O(N__6173),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1145 (
            .O(N__6168),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1144 (
            .O(N__6165),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1143 (
            .O(N__6162),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1142 (
            .O(N__6151),
            .I(N__6148));
    LocalMux I__1141 (
            .O(N__6148),
            .I(N__6145));
    Span4Mux_s1_v I__1140 (
            .O(N__6145),
            .I(N__6142));
    Sp12to4 I__1139 (
            .O(N__6142),
            .I(N__6139));
    Span12Mux_h I__1138 (
            .O(N__6139),
            .I(N__6136));
    Odrv12 I__1137 (
            .O(N__6136),
            .I(CMA_c_10));
    CascadeMux I__1136 (
            .O(N__6133),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_2_cascade_ ));
    InMux I__1135 (
            .O(N__6130),
            .I(N__6126));
    InMux I__1134 (
            .O(N__6129),
            .I(N__6123));
    LocalMux I__1133 (
            .O(N__6126),
            .I(\U712_CHIP_RAM.N_221 ));
    LocalMux I__1132 (
            .O(N__6123),
            .I(\U712_CHIP_RAM.N_221 ));
    CEMux I__1131 (
            .O(N__6118),
            .I(N__6114));
    CEMux I__1130 (
            .O(N__6117),
            .I(N__6111));
    LocalMux I__1129 (
            .O(N__6114),
            .I(N__6106));
    LocalMux I__1128 (
            .O(N__6111),
            .I(N__6106));
    Span4Mux_v I__1127 (
            .O(N__6106),
            .I(N__6103));
    Span4Mux_h I__1126 (
            .O(N__6103),
            .I(N__6100));
    Odrv4 I__1125 (
            .O(N__6100),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ));
    InMux I__1124 (
            .O(N__6097),
            .I(N__6094));
    LocalMux I__1123 (
            .O(N__6094),
            .I(N__6088));
    InMux I__1122 (
            .O(N__6093),
            .I(N__6085));
    InMux I__1121 (
            .O(N__6092),
            .I(N__6080));
    InMux I__1120 (
            .O(N__6091),
            .I(N__6080));
    Odrv12 I__1119 (
            .O(N__6088),
            .I(\U712_CHIP_RAM.N_305 ));
    LocalMux I__1118 (
            .O(N__6085),
            .I(\U712_CHIP_RAM.N_305 ));
    LocalMux I__1117 (
            .O(N__6080),
            .I(\U712_CHIP_RAM.N_305 ));
    CascadeMux I__1116 (
            .O(N__6073),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_cascade_ ));
    InMux I__1115 (
            .O(N__6070),
            .I(N__6067));
    LocalMux I__1114 (
            .O(N__6067),
            .I(N__6063));
    InMux I__1113 (
            .O(N__6066),
            .I(N__6059));
    Span4Mux_v I__1112 (
            .O(N__6063),
            .I(N__6056));
    InMux I__1111 (
            .O(N__6062),
            .I(N__6053));
    LocalMux I__1110 (
            .O(N__6059),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__1109 (
            .O(N__6056),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__1108 (
            .O(N__6053),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    IoInMux I__1107 (
            .O(N__6046),
            .I(N__6043));
    LocalMux I__1106 (
            .O(N__6043),
            .I(N__6040));
    IoSpan4Mux I__1105 (
            .O(N__6040),
            .I(N__6037));
    Span4Mux_s3_h I__1104 (
            .O(N__6037),
            .I(N__6034));
    Sp12to4 I__1103 (
            .O(N__6034),
            .I(N__6031));
    Span12Mux_h I__1102 (
            .O(N__6031),
            .I(N__6027));
    InMux I__1101 (
            .O(N__6030),
            .I(N__6024));
    Odrv12 I__1100 (
            .O(N__6027),
            .I(CLK_EN_c));
    LocalMux I__1099 (
            .O(N__6024),
            .I(CLK_EN_c));
    CascadeMux I__1098 (
            .O(N__6019),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ));
    CascadeMux I__1097 (
            .O(N__6016),
            .I(N__6013));
    InMux I__1096 (
            .O(N__6013),
            .I(N__6009));
    CascadeMux I__1095 (
            .O(N__6012),
            .I(N__6006));
    LocalMux I__1094 (
            .O(N__6009),
            .I(N__5998));
    InMux I__1093 (
            .O(N__6006),
            .I(N__5995));
    CascadeMux I__1092 (
            .O(N__6005),
            .I(N__5992));
    InMux I__1091 (
            .O(N__6004),
            .I(N__5980));
    InMux I__1090 (
            .O(N__6003),
            .I(N__5980));
    InMux I__1089 (
            .O(N__6002),
            .I(N__5980));
    InMux I__1088 (
            .O(N__6001),
            .I(N__5980));
    Span4Mux_h I__1087 (
            .O(N__5998),
            .I(N__5976));
    LocalMux I__1086 (
            .O(N__5995),
            .I(N__5973));
    InMux I__1085 (
            .O(N__5992),
            .I(N__5970));
    InMux I__1084 (
            .O(N__5991),
            .I(N__5967));
    InMux I__1083 (
            .O(N__5990),
            .I(N__5964));
    InMux I__1082 (
            .O(N__5989),
            .I(N__5961));
    LocalMux I__1081 (
            .O(N__5980),
            .I(N__5958));
    InMux I__1080 (
            .O(N__5979),
            .I(N__5955));
    Odrv4 I__1079 (
            .O(N__5976),
            .I(\U712_CHIP_RAM.N_10 ));
    Odrv4 I__1078 (
            .O(N__5973),
            .I(\U712_CHIP_RAM.N_10 ));
    LocalMux I__1077 (
            .O(N__5970),
            .I(\U712_CHIP_RAM.N_10 ));
    LocalMux I__1076 (
            .O(N__5967),
            .I(\U712_CHIP_RAM.N_10 ));
    LocalMux I__1075 (
            .O(N__5964),
            .I(\U712_CHIP_RAM.N_10 ));
    LocalMux I__1074 (
            .O(N__5961),
            .I(\U712_CHIP_RAM.N_10 ));
    Odrv4 I__1073 (
            .O(N__5958),
            .I(\U712_CHIP_RAM.N_10 ));
    LocalMux I__1072 (
            .O(N__5955),
            .I(\U712_CHIP_RAM.N_10 ));
    CascadeMux I__1071 (
            .O(N__5938),
            .I(N__5935));
    InMux I__1070 (
            .O(N__5935),
            .I(N__5932));
    LocalMux I__1069 (
            .O(N__5932),
            .I(\U712_CHIP_RAM.N_260 ));
    CascadeMux I__1068 (
            .O(N__5929),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_66_0_i_1_cascade_ ));
    InMux I__1067 (
            .O(N__5926),
            .I(N__5920));
    InMux I__1066 (
            .O(N__5925),
            .I(N__5920));
    LocalMux I__1065 (
            .O(N__5920),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI9MVM2Z0Z_1 ));
    InMux I__1064 (
            .O(N__5917),
            .I(N__5914));
    LocalMux I__1063 (
            .O(N__5914),
            .I(\U712_CHIP_RAM.N_222 ));
    CascadeMux I__1062 (
            .O(N__5911),
            .I(N__5907));
    InMux I__1061 (
            .O(N__5910),
            .I(N__5904));
    InMux I__1060 (
            .O(N__5907),
            .I(N__5901));
    LocalMux I__1059 (
            .O(N__5904),
            .I(N__5898));
    LocalMux I__1058 (
            .O(N__5901),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa ));
    Odrv12 I__1057 (
            .O(N__5898),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa ));
    CascadeMux I__1056 (
            .O(N__5893),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_9_0_cascade_ ));
    IoInMux I__1055 (
            .O(N__5890),
            .I(N__5887));
    LocalMux I__1054 (
            .O(N__5887),
            .I(N__5884));
    Span4Mux_s1_v I__1053 (
            .O(N__5884),
            .I(N__5881));
    Span4Mux_v I__1052 (
            .O(N__5881),
            .I(N__5878));
    Span4Mux_v I__1051 (
            .O(N__5878),
            .I(N__5875));
    Span4Mux_v I__1050 (
            .O(N__5875),
            .I(N__5870));
    InMux I__1049 (
            .O(N__5874),
            .I(N__5867));
    InMux I__1048 (
            .O(N__5873),
            .I(N__5864));
    Span4Mux_h I__1047 (
            .O(N__5870),
            .I(N__5857));
    LocalMux I__1046 (
            .O(N__5867),
            .I(N__5857));
    LocalMux I__1045 (
            .O(N__5864),
            .I(N__5857));
    Span4Mux_h I__1044 (
            .O(N__5857),
            .I(N__5853));
    InMux I__1043 (
            .O(N__5856),
            .I(N__5850));
    Odrv4 I__1042 (
            .O(N__5853),
            .I(DBENn_c));
    LocalMux I__1041 (
            .O(N__5850),
            .I(DBENn_c));
    InMux I__1040 (
            .O(N__5845),
            .I(N__5842));
    LocalMux I__1039 (
            .O(N__5842),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_3_0 ));
    CascadeMux I__1038 (
            .O(N__5839),
            .I(\U712_CHIP_RAM.N_305_cascade_ ));
    CascadeMux I__1037 (
            .O(N__5836),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_0_cascade_ ));
    CascadeMux I__1036 (
            .O(N__5833),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ));
    InMux I__1035 (
            .O(N__5830),
            .I(N__5827));
    LocalMux I__1034 (
            .O(N__5827),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    InMux I__1033 (
            .O(N__5824),
            .I(N__5821));
    LocalMux I__1032 (
            .O(N__5821),
            .I(N__5818));
    Span4Mux_v I__1031 (
            .O(N__5818),
            .I(N__5815));
    Sp12to4 I__1030 (
            .O(N__5815),
            .I(N__5812));
    Span12Mux_h I__1029 (
            .O(N__5812),
            .I(N__5809));
    Span12Mux_v I__1028 (
            .O(N__5809),
            .I(N__5806));
    Odrv12 I__1027 (
            .O(N__5806),
            .I(A_c_3));
    InMux I__1026 (
            .O(N__5803),
            .I(N__5800));
    LocalMux I__1025 (
            .O(N__5800),
            .I(N__5797));
    Span4Mux_v I__1024 (
            .O(N__5797),
            .I(N__5794));
    Sp12to4 I__1023 (
            .O(N__5794),
            .I(N__5791));
    Span12Mux_h I__1022 (
            .O(N__5791),
            .I(N__5788));
    Odrv12 I__1021 (
            .O(N__5788),
            .I(A_c_10));
    InMux I__1020 (
            .O(N__5785),
            .I(N__5782));
    LocalMux I__1019 (
            .O(N__5782),
            .I(N__5779));
    Span4Mux_v I__1018 (
            .O(N__5779),
            .I(N__5776));
    Sp12to4 I__1017 (
            .O(N__5776),
            .I(N__5773));
    Span12Mux_h I__1016 (
            .O(N__5773),
            .I(N__5770));
    Odrv12 I__1015 (
            .O(N__5770),
            .I(A_c_9));
    InMux I__1014 (
            .O(N__5767),
            .I(N__5764));
    LocalMux I__1013 (
            .O(N__5764),
            .I(N__5761));
    Span12Mux_h I__1012 (
            .O(N__5761),
            .I(N__5758));
    Span12Mux_v I__1011 (
            .O(N__5758),
            .I(N__5755));
    Odrv12 I__1010 (
            .O(N__5755),
            .I(A_c_2));
    InMux I__1009 (
            .O(N__5752),
            .I(N__5749));
    LocalMux I__1008 (
            .O(N__5749),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_0 ));
    CascadeMux I__1007 (
            .O(N__5746),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_1_cascade_ ));
    CascadeMux I__1006 (
            .O(N__5743),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_2_cascade_ ));
    InMux I__1005 (
            .O(N__5740),
            .I(N__5736));
    InMux I__1004 (
            .O(N__5739),
            .I(N__5733));
    LocalMux I__1003 (
            .O(N__5736),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__1002 (
            .O(N__5733),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__1001 (
            .O(N__5728),
            .I(N__5725));
    LocalMux I__1000 (
            .O(N__5725),
            .I(N__5722));
    Span4Mux_v I__999 (
            .O(N__5722),
            .I(N__5719));
    Odrv4 I__998 (
            .O(N__5719),
            .I(TACK_EN_i_ess));
    InMux I__997 (
            .O(N__5716),
            .I(N__5713));
    LocalMux I__996 (
            .O(N__5713),
            .I(N__5710));
    Span4Mux_v I__995 (
            .O(N__5710),
            .I(N__5707));
    Span4Mux_v I__994 (
            .O(N__5707),
            .I(N__5704));
    Sp12to4 I__993 (
            .O(N__5704),
            .I(N__5701));
    Span12Mux_h I__992 (
            .O(N__5701),
            .I(N__5698));
    Odrv12 I__991 (
            .O(N__5698),
            .I(A_c_18));
    InMux I__990 (
            .O(N__5695),
            .I(N__5692));
    LocalMux I__989 (
            .O(N__5692),
            .I(N__5689));
    Span4Mux_v I__988 (
            .O(N__5689),
            .I(N__5686));
    Span4Mux_v I__987 (
            .O(N__5686),
            .I(N__5683));
    Sp12to4 I__986 (
            .O(N__5683),
            .I(N__5680));
    Span12Mux_h I__985 (
            .O(N__5680),
            .I(N__5677));
    Odrv12 I__984 (
            .O(N__5677),
            .I(A_c_16));
    CascadeMux I__983 (
            .O(N__5674),
            .I(N__5671));
    InMux I__982 (
            .O(N__5671),
            .I(N__5668));
    LocalMux I__981 (
            .O(N__5668),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__980 (
            .O(N__5665),
            .I(N__5662));
    LocalMux I__979 (
            .O(N__5662),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__978 (
            .O(N__5659),
            .I(N__5656));
    LocalMux I__977 (
            .O(N__5656),
            .I(N__5653));
    Span12Mux_s5_v I__976 (
            .O(N__5653),
            .I(N__5650));
    Odrv12 I__975 (
            .O(N__5650),
            .I(CMA_c_2));
    IoInMux I__974 (
            .O(N__5647),
            .I(N__5644));
    LocalMux I__973 (
            .O(N__5644),
            .I(N__5641));
    Span12Mux_s8_h I__972 (
            .O(N__5641),
            .I(N__5638));
    Span12Mux_v I__971 (
            .O(N__5638),
            .I(N__5635));
    Odrv12 I__970 (
            .O(N__5635),
            .I(CMA_c_3));
    CascadeMux I__969 (
            .O(N__5632),
            .I(\U712_CHIP_RAM.un1_CMA30_0_i_cascade_ ));
    InMux I__968 (
            .O(N__5629),
            .I(N__5626));
    LocalMux I__967 (
            .O(N__5626),
            .I(N__5623));
    Sp12to4 I__966 (
            .O(N__5623),
            .I(N__5620));
    Span12Mux_v I__965 (
            .O(N__5620),
            .I(N__5617));
    Span12Mux_h I__964 (
            .O(N__5617),
            .I(N__5614));
    Odrv12 I__963 (
            .O(N__5614),
            .I(A_c_5));
    InMux I__962 (
            .O(N__5611),
            .I(N__5608));
    LocalMux I__961 (
            .O(N__5608),
            .I(N__5605));
    Span4Mux_v I__960 (
            .O(N__5605),
            .I(N__5602));
    Sp12to4 I__959 (
            .O(N__5602),
            .I(N__5599));
    Span12Mux_h I__958 (
            .O(N__5599),
            .I(N__5596));
    Odrv12 I__957 (
            .O(N__5596),
            .I(A_c_12));
    CascadeMux I__956 (
            .O(N__5593),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_cascade_ ));
    InMux I__955 (
            .O(N__5590),
            .I(bfn_10_14_0_));
    InMux I__954 (
            .O(N__5587),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__953 (
            .O(N__5584),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__952 (
            .O(N__5581),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    CascadeMux I__951 (
            .O(N__5578),
            .I(N__5575));
    InMux I__950 (
            .O(N__5575),
            .I(N__5571));
    InMux I__949 (
            .O(N__5574),
            .I(N__5568));
    LocalMux I__948 (
            .O(N__5571),
            .I(N__5565));
    LocalMux I__947 (
            .O(N__5568),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    Odrv4 I__946 (
            .O(N__5565),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__945 (
            .O(N__5560),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__944 (
            .O(N__5557),
            .I(N__5553));
    InMux I__943 (
            .O(N__5556),
            .I(N__5550));
    LocalMux I__942 (
            .O(N__5553),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__941 (
            .O(N__5550),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__940 (
            .O(N__5545),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__939 (
            .O(N__5542),
            .I(N__5538));
    InMux I__938 (
            .O(N__5541),
            .I(N__5535));
    LocalMux I__937 (
            .O(N__5538),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__936 (
            .O(N__5535),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__935 (
            .O(N__5530),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__934 (
            .O(N__5527),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    InMux I__933 (
            .O(N__5524),
            .I(N__5521));
    LocalMux I__932 (
            .O(N__5521),
            .I(\U712_CHIP_RAM.N_323 ));
    InMux I__931 (
            .O(N__5518),
            .I(N__5515));
    LocalMux I__930 (
            .O(N__5515),
            .I(\U712_CHIP_RAM.N_240 ));
    CascadeMux I__929 (
            .O(N__5512),
            .I(\U712_CHIP_RAM.N_10_cascade_ ));
    CascadeMux I__928 (
            .O(N__5509),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER16_cascade_ ));
    InMux I__927 (
            .O(N__5506),
            .I(N__5503));
    LocalMux I__926 (
            .O(N__5503),
            .I(N__5500));
    Odrv4 I__925 (
            .O(N__5500),
            .I(\U712_CHIP_RAM.N_328 ));
    InMux I__924 (
            .O(N__5497),
            .I(N__5494));
    LocalMux I__923 (
            .O(N__5494),
            .I(\U712_CHIP_RAM.N_307 ));
    CascadeMux I__922 (
            .O(N__5491),
            .I(\U712_CHIP_RAM.N_328_cascade_ ));
    InMux I__921 (
            .O(N__5488),
            .I(N__5484));
    InMux I__920 (
            .O(N__5487),
            .I(N__5481));
    LocalMux I__919 (
            .O(N__5484),
            .I(\U712_CHIP_RAM.N_177 ));
    LocalMux I__918 (
            .O(N__5481),
            .I(\U712_CHIP_RAM.N_177 ));
    CascadeMux I__917 (
            .O(N__5476),
            .I(\U712_CHIP_RAM.N_251_cascade_ ));
    InMux I__916 (
            .O(N__5473),
            .I(N__5470));
    LocalMux I__915 (
            .O(N__5470),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0 ));
    CascadeMux I__914 (
            .O(N__5467),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a3_3_2_0_cascade_ ));
    CascadeMux I__913 (
            .O(N__5464),
            .I(\U712_CHIP_RAM.N_242_cascade_ ));
    CascadeMux I__912 (
            .O(N__5461),
            .I(\U712_CHIP_RAM.N_188_cascade_ ));
    CEMux I__911 (
            .O(N__5458),
            .I(N__5455));
    LocalMux I__910 (
            .O(N__5455),
            .I(N__5452));
    Sp12to4 I__909 (
            .O(N__5452),
            .I(N__5449));
    Odrv12 I__908 (
            .O(N__5449),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0_0 ));
    InMux I__907 (
            .O(N__5446),
            .I(N__5438));
    InMux I__906 (
            .O(N__5445),
            .I(N__5438));
    InMux I__905 (
            .O(N__5444),
            .I(N__5433));
    InMux I__904 (
            .O(N__5443),
            .I(N__5433));
    LocalMux I__903 (
            .O(N__5438),
            .I(\U712_CHIP_RAM.N_306 ));
    LocalMux I__902 (
            .O(N__5433),
            .I(\U712_CHIP_RAM.N_306 ));
    InMux I__901 (
            .O(N__5428),
            .I(N__5423));
    InMux I__900 (
            .O(N__5427),
            .I(N__5420));
    InMux I__899 (
            .O(N__5426),
            .I(N__5417));
    LocalMux I__898 (
            .O(N__5423),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__897 (
            .O(N__5420),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__896 (
            .O(N__5417),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__895 (
            .O(N__5410),
            .I(N__5407));
    LocalMux I__894 (
            .O(N__5407),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0 ));
    InMux I__893 (
            .O(N__5404),
            .I(N__5401));
    LocalMux I__892 (
            .O(N__5401),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0 ));
    InMux I__891 (
            .O(N__5398),
            .I(N__5394));
    InMux I__890 (
            .O(N__5397),
            .I(N__5391));
    LocalMux I__889 (
            .O(N__5394),
            .I(\U712_CHIP_RAM.N_238 ));
    LocalMux I__888 (
            .O(N__5391),
            .I(\U712_CHIP_RAM.N_238 ));
    CascadeMux I__887 (
            .O(N__5386),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_ ));
    InMux I__886 (
            .O(N__5383),
            .I(N__5379));
    InMux I__885 (
            .O(N__5382),
            .I(N__5376));
    LocalMux I__884 (
            .O(N__5379),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    LocalMux I__883 (
            .O(N__5376),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    InMux I__882 (
            .O(N__5371),
            .I(N__5368));
    LocalMux I__881 (
            .O(N__5368),
            .I(N__5365));
    Span4Mux_v I__880 (
            .O(N__5365),
            .I(N__5362));
    Odrv4 I__879 (
            .O(N__5362),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    InMux I__878 (
            .O(N__5359),
            .I(N__5356));
    LocalMux I__877 (
            .O(N__5356),
            .I(N__5353));
    Span12Mux_v I__876 (
            .O(N__5353),
            .I(N__5350));
    Span12Mux_h I__875 (
            .O(N__5350),
            .I(N__5347));
    Odrv12 I__874 (
            .O(N__5347),
            .I(A_c_4));
    InMux I__873 (
            .O(N__5344),
            .I(N__5341));
    LocalMux I__872 (
            .O(N__5341),
            .I(N__5338));
    Span4Mux_v I__871 (
            .O(N__5338),
            .I(N__5335));
    Sp12to4 I__870 (
            .O(N__5335),
            .I(N__5332));
    Span12Mux_h I__869 (
            .O(N__5332),
            .I(N__5329));
    Odrv12 I__868 (
            .O(N__5329),
            .I(A_c_11));
    CascadeMux I__867 (
            .O(N__5326),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ));
    SRMux I__866 (
            .O(N__5323),
            .I(N__5320));
    LocalMux I__865 (
            .O(N__5320),
            .I(N__5317));
    Odrv12 I__864 (
            .O(N__5317),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    CascadeMux I__863 (
            .O(N__5314),
            .I(N__5311));
    InMux I__862 (
            .O(N__5311),
            .I(N__5304));
    InMux I__861 (
            .O(N__5310),
            .I(N__5304));
    InMux I__860 (
            .O(N__5309),
            .I(N__5301));
    LocalMux I__859 (
            .O(N__5304),
            .I(N__5296));
    LocalMux I__858 (
            .O(N__5301),
            .I(N__5296));
    Odrv4 I__857 (
            .O(N__5296),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    InMux I__856 (
            .O(N__5293),
            .I(N__5286));
    InMux I__855 (
            .O(N__5292),
            .I(N__5286));
    InMux I__854 (
            .O(N__5291),
            .I(N__5283));
    LocalMux I__853 (
            .O(N__5286),
            .I(\U712_REG_SM.N_209 ));
    LocalMux I__852 (
            .O(N__5283),
            .I(\U712_REG_SM.N_209 ));
    InMux I__851 (
            .O(N__5278),
            .I(N__5275));
    LocalMux I__850 (
            .O(N__5275),
            .I(N__5272));
    Span4Mux_v I__849 (
            .O(N__5272),
            .I(N__5269));
    Span4Mux_v I__848 (
            .O(N__5269),
            .I(N__5264));
    InMux I__847 (
            .O(N__5268),
            .I(N__5261));
    InMux I__846 (
            .O(N__5267),
            .I(N__5258));
    Span4Mux_v I__845 (
            .O(N__5264),
            .I(N__5253));
    LocalMux I__844 (
            .O(N__5261),
            .I(N__5253));
    LocalMux I__843 (
            .O(N__5258),
            .I(N__5250));
    Span4Mux_v I__842 (
            .O(N__5253),
            .I(N__5247));
    Span12Mux_h I__841 (
            .O(N__5250),
            .I(N__5244));
    IoSpan4Mux I__840 (
            .O(N__5247),
            .I(N__5241));
    Span12Mux_v I__839 (
            .O(N__5244),
            .I(N__5238));
    IoSpan4Mux I__838 (
            .O(N__5241),
            .I(N__5235));
    Odrv12 I__837 (
            .O(N__5238),
            .I(AWEn_c));
    Odrv4 I__836 (
            .O(N__5235),
            .I(AWEn_c));
    IoInMux I__835 (
            .O(N__5230),
            .I(N__5227));
    LocalMux I__834 (
            .O(N__5227),
            .I(N__5224));
    IoSpan4Mux I__833 (
            .O(N__5224),
            .I(N__5221));
    Span4Mux_s3_v I__832 (
            .O(N__5221),
            .I(N__5218));
    Sp12to4 I__831 (
            .O(N__5218),
            .I(N__5214));
    InMux I__830 (
            .O(N__5217),
            .I(N__5211));
    Odrv12 I__829 (
            .O(N__5214),
            .I(DBDIR_c));
    LocalMux I__828 (
            .O(N__5211),
            .I(DBDIR_c));
    CascadeMux I__827 (
            .O(N__5206),
            .I(\U712_CHIP_RAM.N_323_cascade_ ));
    InMux I__826 (
            .O(N__5203),
            .I(N__5200));
    LocalMux I__825 (
            .O(N__5200),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a2_0_0_0 ));
    InMux I__824 (
            .O(N__5197),
            .I(N__5193));
    InMux I__823 (
            .O(N__5196),
            .I(N__5190));
    LocalMux I__822 (
            .O(N__5193),
            .I(N__5187));
    LocalMux I__821 (
            .O(N__5190),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    Odrv12 I__820 (
            .O(N__5187),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__819 (
            .O(N__5182),
            .I(N__5178));
    InMux I__818 (
            .O(N__5181),
            .I(N__5175));
    LocalMux I__817 (
            .O(N__5178),
            .I(N__5172));
    LocalMux I__816 (
            .O(N__5175),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    Odrv12 I__815 (
            .O(N__5172),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__814 (
            .O(N__5167),
            .I(N__5164));
    LocalMux I__813 (
            .O(N__5164),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ));
    CascadeMux I__812 (
            .O(N__5161),
            .I(\U712_CHIP_RAM.N_307_cascade_ ));
    CascadeMux I__811 (
            .O(N__5158),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_cascade_ ));
    InMux I__810 (
            .O(N__5155),
            .I(N__5149));
    InMux I__809 (
            .O(N__5154),
            .I(N__5149));
    LocalMux I__808 (
            .O(N__5149),
            .I(N__5146));
    Span4Mux_v I__807 (
            .O(N__5146),
            .I(N__5142));
    InMux I__806 (
            .O(N__5145),
            .I(N__5139));
    Span4Mux_v I__805 (
            .O(N__5142),
            .I(N__5134));
    LocalMux I__804 (
            .O(N__5139),
            .I(N__5134));
    Span4Mux_h I__803 (
            .O(N__5134),
            .I(N__5131));
    Sp12to4 I__802 (
            .O(N__5131),
            .I(N__5128));
    Span12Mux_v I__801 (
            .O(N__5128),
            .I(N__5125));
    Span12Mux_h I__800 (
            .O(N__5125),
            .I(N__5122));
    Odrv12 I__799 (
            .O(N__5122),
            .I(CASUn_c));
    CascadeMux I__798 (
            .O(N__5119),
            .I(N__5116));
    InMux I__797 (
            .O(N__5116),
            .I(N__5110));
    InMux I__796 (
            .O(N__5115),
            .I(N__5110));
    LocalMux I__795 (
            .O(N__5110),
            .I(N__5106));
    InMux I__794 (
            .O(N__5109),
            .I(N__5103));
    Span4Mux_v I__793 (
            .O(N__5106),
            .I(N__5100));
    LocalMux I__792 (
            .O(N__5103),
            .I(N__5097));
    Sp12to4 I__791 (
            .O(N__5100),
            .I(N__5094));
    Sp12to4 I__790 (
            .O(N__5097),
            .I(N__5091));
    Span12Mux_h I__789 (
            .O(N__5094),
            .I(N__5088));
    Span12Mux_v I__788 (
            .O(N__5091),
            .I(N__5085));
    Span12Mux_v I__787 (
            .O(N__5088),
            .I(N__5082));
    Span12Mux_h I__786 (
            .O(N__5085),
            .I(N__5079));
    Odrv12 I__785 (
            .O(N__5082),
            .I(CASLn_c));
    Odrv12 I__784 (
            .O(N__5079),
            .I(CASLn_c));
    InMux I__783 (
            .O(N__5074),
            .I(N__5068));
    InMux I__782 (
            .O(N__5073),
            .I(N__5068));
    LocalMux I__781 (
            .O(N__5068),
            .I(N__5065));
    Odrv4 I__780 (
            .O(N__5065),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__779 (
            .O(N__5062),
            .I(N__5058));
    InMux I__778 (
            .O(N__5061),
            .I(N__5055));
    LocalMux I__777 (
            .O(N__5058),
            .I(N__5052));
    LocalMux I__776 (
            .O(N__5055),
            .I(U712_REG_SM_DBR_SYNC_0));
    Odrv12 I__775 (
            .O(N__5052),
            .I(U712_REG_SM_DBR_SYNC_0));
    InMux I__774 (
            .O(N__5047),
            .I(N__5043));
    InMux I__773 (
            .O(N__5046),
            .I(N__5040));
    LocalMux I__772 (
            .O(N__5043),
            .I(N__5036));
    LocalMux I__771 (
            .O(N__5040),
            .I(N__5033));
    InMux I__770 (
            .O(N__5039),
            .I(N__5030));
    Odrv4 I__769 (
            .O(N__5036),
            .I(\U712_REG_SM.DS_ENZ0 ));
    Odrv4 I__768 (
            .O(N__5033),
            .I(\U712_REG_SM.DS_ENZ0 ));
    LocalMux I__767 (
            .O(N__5030),
            .I(\U712_REG_SM.DS_ENZ0 ));
    InMux I__766 (
            .O(N__5023),
            .I(N__5020));
    LocalMux I__765 (
            .O(N__5020),
            .I(N__5016));
    CascadeMux I__764 (
            .O(N__5019),
            .I(N__5013));
    Span4Mux_v I__763 (
            .O(N__5016),
            .I(N__5010));
    InMux I__762 (
            .O(N__5013),
            .I(N__5007));
    Odrv4 I__761 (
            .O(N__5010),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    LocalMux I__760 (
            .O(N__5007),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    IoInMux I__759 (
            .O(N__5002),
            .I(N__4999));
    LocalMux I__758 (
            .O(N__4999),
            .I(N__4996));
    Span12Mux_s11_v I__757 (
            .O(N__4996),
            .I(N__4993));
    Span12Mux_h I__756 (
            .O(N__4993),
            .I(N__4990));
    Odrv12 I__755 (
            .O(N__4990),
            .I(U712_REG_SM_un1_UDSn_i));
    InMux I__754 (
            .O(N__4987),
            .I(N__4980));
    InMux I__753 (
            .O(N__4986),
            .I(N__4980));
    InMux I__752 (
            .O(N__4985),
            .I(N__4977));
    LocalMux I__751 (
            .O(N__4980),
            .I(N__4973));
    LocalMux I__750 (
            .O(N__4977),
            .I(N__4970));
    InMux I__749 (
            .O(N__4976),
            .I(N__4966));
    Span4Mux_v I__748 (
            .O(N__4973),
            .I(N__4963));
    Span4Mux_v I__747 (
            .O(N__4970),
            .I(N__4960));
    InMux I__746 (
            .O(N__4969),
            .I(N__4957));
    LocalMux I__745 (
            .O(N__4966),
            .I(N__4954));
    Sp12to4 I__744 (
            .O(N__4963),
            .I(N__4947));
    Sp12to4 I__743 (
            .O(N__4960),
            .I(N__4947));
    LocalMux I__742 (
            .O(N__4957),
            .I(N__4947));
    Span4Mux_v I__741 (
            .O(N__4954),
            .I(N__4944));
    Span12Mux_h I__740 (
            .O(N__4947),
            .I(N__4941));
    Sp12to4 I__739 (
            .O(N__4944),
            .I(N__4938));
    Span12Mux_v I__738 (
            .O(N__4941),
            .I(N__4935));
    Span12Mux_h I__737 (
            .O(N__4938),
            .I(N__4932));
    Odrv12 I__736 (
            .O(N__4935),
            .I(RnW_c));
    Odrv12 I__735 (
            .O(N__4932),
            .I(RnW_c));
    IoInMux I__734 (
            .O(N__4927),
            .I(N__4924));
    LocalMux I__733 (
            .O(N__4924),
            .I(N__4921));
    Span4Mux_s2_h I__732 (
            .O(N__4921),
            .I(N__4918));
    Sp12to4 I__731 (
            .O(N__4918),
            .I(N__4915));
    Span12Mux_s6_v I__730 (
            .O(N__4915),
            .I(N__4912));
    Span12Mux_h I__729 (
            .O(N__4912),
            .I(N__4909));
    Odrv12 I__728 (
            .O(N__4909),
            .I(DRDDIR_i_m4_i_m2));
    InMux I__727 (
            .O(N__4906),
            .I(N__4902));
    InMux I__726 (
            .O(N__4905),
            .I(N__4899));
    LocalMux I__725 (
            .O(N__4902),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    LocalMux I__724 (
            .O(N__4899),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__723 (
            .O(N__4894),
            .I(N__4890));
    InMux I__722 (
            .O(N__4893),
            .I(N__4887));
    LocalMux I__721 (
            .O(N__4890),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    LocalMux I__720 (
            .O(N__4887),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    CascadeMux I__719 (
            .O(N__4882),
            .I(N__4878));
    InMux I__718 (
            .O(N__4881),
            .I(N__4875));
    InMux I__717 (
            .O(N__4878),
            .I(N__4872));
    LocalMux I__716 (
            .O(N__4875),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__715 (
            .O(N__4872),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    CascadeMux I__714 (
            .O(N__4867),
            .I(N__4864));
    InMux I__713 (
            .O(N__4864),
            .I(N__4861));
    LocalMux I__712 (
            .O(N__4861),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_RNOZ0Z_0 ));
    CascadeMux I__711 (
            .O(N__4858),
            .I(N__4850));
    InMux I__710 (
            .O(N__4857),
            .I(N__4847));
    InMux I__709 (
            .O(N__4856),
            .I(N__4844));
    CascadeMux I__708 (
            .O(N__4855),
            .I(N__4841));
    CascadeMux I__707 (
            .O(N__4854),
            .I(N__4838));
    CascadeMux I__706 (
            .O(N__4853),
            .I(N__4835));
    InMux I__705 (
            .O(N__4850),
            .I(N__4832));
    LocalMux I__704 (
            .O(N__4847),
            .I(N__4825));
    LocalMux I__703 (
            .O(N__4844),
            .I(N__4825));
    InMux I__702 (
            .O(N__4841),
            .I(N__4820));
    InMux I__701 (
            .O(N__4838),
            .I(N__4820));
    InMux I__700 (
            .O(N__4835),
            .I(N__4817));
    LocalMux I__699 (
            .O(N__4832),
            .I(N__4814));
    InMux I__698 (
            .O(N__4831),
            .I(N__4809));
    InMux I__697 (
            .O(N__4830),
            .I(N__4809));
    Odrv4 I__696 (
            .O(N__4825),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__695 (
            .O(N__4820),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__694 (
            .O(N__4817),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    Odrv4 I__693 (
            .O(N__4814),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__692 (
            .O(N__4809),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__691 (
            .O(N__4798),
            .I(N__4795));
    LocalMux I__690 (
            .O(N__4795),
            .I(\U712_REG_SM.N_265 ));
    InMux I__689 (
            .O(N__4792),
            .I(N__4788));
    InMux I__688 (
            .O(N__4791),
            .I(N__4785));
    LocalMux I__687 (
            .O(N__4788),
            .I(\U712_REG_SM.N_183 ));
    LocalMux I__686 (
            .O(N__4785),
            .I(\U712_REG_SM.N_183 ));
    InMux I__685 (
            .O(N__4780),
            .I(N__4777));
    LocalMux I__684 (
            .O(N__4777),
            .I(N__4772));
    InMux I__683 (
            .O(N__4776),
            .I(N__4769));
    InMux I__682 (
            .O(N__4775),
            .I(N__4766));
    Odrv4 I__681 (
            .O(N__4772),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__680 (
            .O(N__4769),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__679 (
            .O(N__4766),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    InMux I__678 (
            .O(N__4759),
            .I(N__4753));
    InMux I__677 (
            .O(N__4758),
            .I(N__4750));
    InMux I__676 (
            .O(N__4757),
            .I(N__4747));
    InMux I__675 (
            .O(N__4756),
            .I(N__4744));
    LocalMux I__674 (
            .O(N__4753),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__673 (
            .O(N__4750),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__672 (
            .O(N__4747),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__671 (
            .O(N__4744),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__670 (
            .O(N__4735),
            .I(N__4731));
    InMux I__669 (
            .O(N__4734),
            .I(N__4728));
    LocalMux I__668 (
            .O(N__4731),
            .I(N__4725));
    LocalMux I__667 (
            .O(N__4728),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    Odrv12 I__666 (
            .O(N__4725),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    CascadeMux I__665 (
            .O(N__4720),
            .I(N__4717));
    InMux I__664 (
            .O(N__4717),
            .I(N__4713));
    InMux I__663 (
            .O(N__4716),
            .I(N__4710));
    LocalMux I__662 (
            .O(N__4713),
            .I(N__4707));
    LocalMux I__661 (
            .O(N__4710),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv4 I__660 (
            .O(N__4707),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__659 (
            .O(N__4702),
            .I(N__4699));
    LocalMux I__658 (
            .O(N__4699),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__657 (
            .O(N__4696),
            .I(N__4693));
    LocalMux I__656 (
            .O(N__4693),
            .I(N__4689));
    InMux I__655 (
            .O(N__4692),
            .I(N__4685));
    Span4Mux_h I__654 (
            .O(N__4689),
            .I(N__4682));
    InMux I__653 (
            .O(N__4688),
            .I(N__4679));
    LocalMux I__652 (
            .O(N__4685),
            .I(U712_REG_SM_DBR_SYNC_1));
    Odrv4 I__651 (
            .O(N__4682),
            .I(U712_REG_SM_DBR_SYNC_1));
    LocalMux I__650 (
            .O(N__4679),
            .I(U712_REG_SM_DBR_SYNC_1));
    InMux I__649 (
            .O(N__4672),
            .I(N__4669));
    LocalMux I__648 (
            .O(N__4669),
            .I(\U712_CHIP_RAM.DBR_SYNCZ0Z_2 ));
    InMux I__647 (
            .O(N__4666),
            .I(N__4662));
    InMux I__646 (
            .O(N__4665),
            .I(N__4659));
    LocalMux I__645 (
            .O(N__4662),
            .I(N__4656));
    LocalMux I__644 (
            .O(N__4659),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv4 I__643 (
            .O(N__4656),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__642 (
            .O(N__4651),
            .I(\U712_CHIP_RAM.N_177_cascade_ ));
    InMux I__641 (
            .O(N__4648),
            .I(N__4645));
    LocalMux I__640 (
            .O(N__4645),
            .I(N__4641));
    InMux I__639 (
            .O(N__4644),
            .I(N__4638));
    Odrv4 I__638 (
            .O(N__4641),
            .I(\U712_CHIP_RAM.N_197 ));
    LocalMux I__637 (
            .O(N__4638),
            .I(\U712_CHIP_RAM.N_197 ));
    InMux I__636 (
            .O(N__4633),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__635 (
            .O(N__4630),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__634 (
            .O(N__4627),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__633 (
            .O(N__4624),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    InMux I__632 (
            .O(N__4621),
            .I(N__4617));
    InMux I__631 (
            .O(N__4620),
            .I(N__4614));
    LocalMux I__630 (
            .O(N__4617),
            .I(N__4611));
    LocalMux I__629 (
            .O(N__4614),
            .I(N__4608));
    Span4Mux_v I__628 (
            .O(N__4611),
            .I(N__4605));
    Span4Mux_v I__627 (
            .O(N__4608),
            .I(N__4602));
    Sp12to4 I__626 (
            .O(N__4605),
            .I(N__4599));
    Span4Mux_h I__625 (
            .O(N__4602),
            .I(N__4596));
    Span12Mux_h I__624 (
            .O(N__4599),
            .I(N__4591));
    Sp12to4 I__623 (
            .O(N__4596),
            .I(N__4591));
    Span12Mux_v I__622 (
            .O(N__4591),
            .I(N__4588));
    Odrv12 I__621 (
            .O(N__4588),
            .I(TSn_c));
    CascadeMux I__620 (
            .O(N__4585),
            .I(N__4582));
    InMux I__619 (
            .O(N__4582),
            .I(N__4579));
    LocalMux I__618 (
            .O(N__4579),
            .I(N__4576));
    Span4Mux_v I__617 (
            .O(N__4576),
            .I(N__4573));
    Sp12to4 I__616 (
            .O(N__4573),
            .I(N__4570));
    Span12Mux_h I__615 (
            .O(N__4570),
            .I(N__4567));
    Span12Mux_v I__614 (
            .O(N__4567),
            .I(N__4564));
    Odrv12 I__613 (
            .O(N__4564),
            .I(RAMSPACEn_c));
    InMux I__612 (
            .O(N__4561),
            .I(N__4557));
    InMux I__611 (
            .O(N__4560),
            .I(N__4552));
    LocalMux I__610 (
            .O(N__4557),
            .I(N__4549));
    InMux I__609 (
            .O(N__4556),
            .I(N__4546));
    InMux I__608 (
            .O(N__4555),
            .I(N__4543));
    LocalMux I__607 (
            .O(N__4552),
            .I(N__4540));
    Odrv4 I__606 (
            .O(N__4549),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__605 (
            .O(N__4546),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__604 (
            .O(N__4543),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    Odrv12 I__603 (
            .O(N__4540),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__602 (
            .O(N__4531),
            .I(N__4527));
    InMux I__601 (
            .O(N__4530),
            .I(N__4524));
    LocalMux I__600 (
            .O(N__4527),
            .I(N__4519));
    LocalMux I__599 (
            .O(N__4524),
            .I(N__4519));
    Odrv4 I__598 (
            .O(N__4519),
            .I(\U712_REG_SM.N_325 ));
    InMux I__597 (
            .O(N__4516),
            .I(N__4512));
    CascadeMux I__596 (
            .O(N__4515),
            .I(N__4509));
    LocalMux I__595 (
            .O(N__4512),
            .I(N__4505));
    InMux I__594 (
            .O(N__4509),
            .I(N__4502));
    InMux I__593 (
            .O(N__4508),
            .I(N__4496));
    Span4Mux_h I__592 (
            .O(N__4505),
            .I(N__4493));
    LocalMux I__591 (
            .O(N__4502),
            .I(N__4490));
    InMux I__590 (
            .O(N__4501),
            .I(N__4487));
    InMux I__589 (
            .O(N__4500),
            .I(N__4482));
    InMux I__588 (
            .O(N__4499),
            .I(N__4482));
    LocalMux I__587 (
            .O(N__4496),
            .I(\U712_REG_SM.N_201 ));
    Odrv4 I__586 (
            .O(N__4493),
            .I(\U712_REG_SM.N_201 ));
    Odrv4 I__585 (
            .O(N__4490),
            .I(\U712_REG_SM.N_201 ));
    LocalMux I__584 (
            .O(N__4487),
            .I(\U712_REG_SM.N_201 ));
    LocalMux I__583 (
            .O(N__4482),
            .I(\U712_REG_SM.N_201 ));
    CascadeMux I__582 (
            .O(N__4471),
            .I(N__4468));
    InMux I__581 (
            .O(N__4468),
            .I(N__4463));
    InMux I__580 (
            .O(N__4467),
            .I(N__4460));
    CascadeMux I__579 (
            .O(N__4466),
            .I(N__4457));
    LocalMux I__578 (
            .O(N__4463),
            .I(N__4452));
    LocalMux I__577 (
            .O(N__4460),
            .I(N__4452));
    InMux I__576 (
            .O(N__4457),
            .I(N__4449));
    Span4Mux_v I__575 (
            .O(N__4452),
            .I(N__4446));
    LocalMux I__574 (
            .O(N__4449),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    Odrv4 I__573 (
            .O(N__4446),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    InMux I__572 (
            .O(N__4441),
            .I(N__4437));
    IoInMux I__571 (
            .O(N__4440),
            .I(N__4434));
    LocalMux I__570 (
            .O(N__4437),
            .I(N__4431));
    LocalMux I__569 (
            .O(N__4434),
            .I(N__4428));
    Span4Mux_v I__568 (
            .O(N__4431),
            .I(N__4425));
    IoSpan4Mux I__567 (
            .O(N__4428),
            .I(N__4422));
    Sp12to4 I__566 (
            .O(N__4425),
            .I(N__4419));
    IoSpan4Mux I__565 (
            .O(N__4422),
            .I(N__4416));
    Span12Mux_h I__564 (
            .O(N__4419),
            .I(N__4413));
    IoSpan4Mux I__563 (
            .O(N__4416),
            .I(N__4410));
    Odrv12 I__562 (
            .O(N__4413),
            .I(C3_c));
    Odrv4 I__561 (
            .O(N__4410),
            .I(C3_c));
    InMux I__560 (
            .O(N__4405),
            .I(N__4400));
    InMux I__559 (
            .O(N__4404),
            .I(N__4394));
    InMux I__558 (
            .O(N__4403),
            .I(N__4394));
    LocalMux I__557 (
            .O(N__4400),
            .I(N__4391));
    InMux I__556 (
            .O(N__4399),
            .I(N__4388));
    LocalMux I__555 (
            .O(N__4394),
            .I(N__4385));
    Odrv12 I__554 (
            .O(N__4391),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__553 (
            .O(N__4388),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    Odrv4 I__552 (
            .O(N__4385),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    CascadeMux I__551 (
            .O(N__4378),
            .I(N__4374));
    InMux I__550 (
            .O(N__4377),
            .I(N__4371));
    InMux I__549 (
            .O(N__4374),
            .I(N__4368));
    LocalMux I__548 (
            .O(N__4371),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    LocalMux I__547 (
            .O(N__4368),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    IoInMux I__546 (
            .O(N__4363),
            .I(N__4360));
    LocalMux I__545 (
            .O(N__4360),
            .I(N__4357));
    IoSpan4Mux I__544 (
            .O(N__4357),
            .I(N__4354));
    IoSpan4Mux I__543 (
            .O(N__4354),
            .I(N__4351));
    Span4Mux_s0_v I__542 (
            .O(N__4351),
            .I(N__4348));
    Sp12to4 I__541 (
            .O(N__4348),
            .I(N__4345));
    Span12Mux_v I__540 (
            .O(N__4345),
            .I(N__4342));
    Odrv12 I__539 (
            .O(N__4342),
            .I(U712_REG_SM_un1_LDSn_i));
    InMux I__538 (
            .O(N__4339),
            .I(N__4333));
    InMux I__537 (
            .O(N__4338),
            .I(N__4333));
    LocalMux I__536 (
            .O(N__4333),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0 ));
    InMux I__535 (
            .O(N__4330),
            .I(bfn_9_9_0_));
    InMux I__534 (
            .O(N__4327),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__533 (
            .O(N__4324),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__532 (
            .O(N__4321),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    CascadeMux I__531 (
            .O(N__4318),
            .I(\U712_REG_SM.N_215_cascade_ ));
    CascadeMux I__530 (
            .O(N__4315),
            .I(\U712_REG_SM.N_200_cascade_ ));
    InMux I__529 (
            .O(N__4312),
            .I(N__4308));
    InMux I__528 (
            .O(N__4311),
            .I(N__4305));
    LocalMux I__527 (
            .O(N__4308),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    LocalMux I__526 (
            .O(N__4305),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    InMux I__525 (
            .O(N__4300),
            .I(N__4296));
    InMux I__524 (
            .O(N__4299),
            .I(N__4293));
    LocalMux I__523 (
            .O(N__4296),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    LocalMux I__522 (
            .O(N__4293),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    InMux I__521 (
            .O(N__4288),
            .I(N__4281));
    InMux I__520 (
            .O(N__4287),
            .I(N__4281));
    InMux I__519 (
            .O(N__4286),
            .I(N__4278));
    LocalMux I__518 (
            .O(N__4281),
            .I(\U712_REG_SM.N_200 ));
    LocalMux I__517 (
            .O(N__4278),
            .I(\U712_REG_SM.N_200 ));
    InMux I__516 (
            .O(N__4273),
            .I(N__4269));
    InMux I__515 (
            .O(N__4272),
            .I(N__4266));
    LocalMux I__514 (
            .O(N__4269),
            .I(\U712_REG_SM.N_219 ));
    LocalMux I__513 (
            .O(N__4266),
            .I(\U712_REG_SM.N_219 ));
    CascadeMux I__512 (
            .O(N__4261),
            .I(\U712_REG_SM.N_325_cascade_ ));
    CascadeMux I__511 (
            .O(N__4258),
            .I(N__4249));
    InMux I__510 (
            .O(N__4257),
            .I(N__4246));
    InMux I__509 (
            .O(N__4256),
            .I(N__4241));
    InMux I__508 (
            .O(N__4255),
            .I(N__4241));
    InMux I__507 (
            .O(N__4254),
            .I(N__4238));
    InMux I__506 (
            .O(N__4253),
            .I(N__4231));
    InMux I__505 (
            .O(N__4252),
            .I(N__4231));
    InMux I__504 (
            .O(N__4249),
            .I(N__4231));
    LocalMux I__503 (
            .O(N__4246),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__502 (
            .O(N__4241),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__501 (
            .O(N__4238),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__500 (
            .O(N__4231),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    InMux I__499 (
            .O(N__4222),
            .I(N__4219));
    LocalMux I__498 (
            .O(N__4219),
            .I(N__4216));
    Odrv4 I__497 (
            .O(N__4216),
            .I(\U712_REG_SM.N_198 ));
    InMux I__496 (
            .O(N__4213),
            .I(N__4210));
    LocalMux I__495 (
            .O(N__4210),
            .I(N__4205));
    InMux I__494 (
            .O(N__4209),
            .I(N__4202));
    InMux I__493 (
            .O(N__4208),
            .I(N__4199));
    Odrv4 I__492 (
            .O(N__4205),
            .I(\U712_REG_SM.N_212 ));
    LocalMux I__491 (
            .O(N__4202),
            .I(\U712_REG_SM.N_212 ));
    LocalMux I__490 (
            .O(N__4199),
            .I(\U712_REG_SM.N_212 ));
    InMux I__489 (
            .O(N__4192),
            .I(N__4187));
    InMux I__488 (
            .O(N__4191),
            .I(N__4184));
    InMux I__487 (
            .O(N__4190),
            .I(N__4181));
    LocalMux I__486 (
            .O(N__4187),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__485 (
            .O(N__4184),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__484 (
            .O(N__4181),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    CascadeMux I__483 (
            .O(N__4174),
            .I(\U712_REG_SM.N_198_cascade_ ));
    CascadeMux I__482 (
            .O(N__4171),
            .I(\U712_REG_SM.DS_EN_RNOZ0Z_0_cascade_ ));
    CascadeMux I__481 (
            .O(N__4168),
            .I(\U712_BYTE_ENABLE.N_271_cascade_ ));
    IoInMux I__480 (
            .O(N__4165),
            .I(N__4162));
    LocalMux I__479 (
            .O(N__4162),
            .I(N__4159));
    Span4Mux_s3_h I__478 (
            .O(N__4159),
            .I(N__4156));
    Span4Mux_v I__477 (
            .O(N__4156),
            .I(N__4153));
    Sp12to4 I__476 (
            .O(N__4153),
            .I(N__4150));
    Span12Mux_s11_h I__475 (
            .O(N__4150),
            .I(N__4147));
    Odrv12 I__474 (
            .O(N__4147),
            .I(N_44_i));
    InMux I__473 (
            .O(N__4144),
            .I(N__4135));
    InMux I__472 (
            .O(N__4143),
            .I(N__4135));
    InMux I__471 (
            .O(N__4142),
            .I(N__4135));
    LocalMux I__470 (
            .O(N__4135),
            .I(N__4131));
    InMux I__469 (
            .O(N__4134),
            .I(N__4128));
    Span4Mux_h I__468 (
            .O(N__4131),
            .I(N__4121));
    LocalMux I__467 (
            .O(N__4128),
            .I(N__4121));
    InMux I__466 (
            .O(N__4127),
            .I(N__4118));
    InMux I__465 (
            .O(N__4126),
            .I(N__4115));
    Span4Mux_v I__464 (
            .O(N__4121),
            .I(N__4110));
    LocalMux I__463 (
            .O(N__4118),
            .I(N__4110));
    LocalMux I__462 (
            .O(N__4115),
            .I(N__4107));
    Span4Mux_v I__461 (
            .O(N__4110),
            .I(N__4104));
    Span12Mux_v I__460 (
            .O(N__4107),
            .I(N__4099));
    Sp12to4 I__459 (
            .O(N__4104),
            .I(N__4099));
    Odrv12 I__458 (
            .O(N__4099),
            .I(A_c_0));
    InMux I__457 (
            .O(N__4096),
            .I(N__4086));
    InMux I__456 (
            .O(N__4095),
            .I(N__4086));
    InMux I__455 (
            .O(N__4094),
            .I(N__4086));
    InMux I__454 (
            .O(N__4093),
            .I(N__4083));
    LocalMux I__453 (
            .O(N__4086),
            .I(N__4078));
    LocalMux I__452 (
            .O(N__4083),
            .I(N__4078));
    Span12Mux_v I__451 (
            .O(N__4078),
            .I(N__4075));
    Odrv12 I__450 (
            .O(N__4075),
            .I(A_c_1));
    InMux I__449 (
            .O(N__4072),
            .I(N__4069));
    LocalMux I__448 (
            .O(N__4069),
            .I(\U712_BYTE_ENABLE.N_277 ));
    CascadeMux I__447 (
            .O(N__4066),
            .I(N__4063));
    InMux I__446 (
            .O(N__4063),
            .I(N__4059));
    CascadeMux I__445 (
            .O(N__4062),
            .I(N__4056));
    LocalMux I__444 (
            .O(N__4059),
            .I(N__4052));
    InMux I__443 (
            .O(N__4056),
            .I(N__4047));
    InMux I__442 (
            .O(N__4055),
            .I(N__4047));
    Span4Mux_h I__441 (
            .O(N__4052),
            .I(N__4042));
    LocalMux I__440 (
            .O(N__4047),
            .I(N__4042));
    Span4Mux_v I__439 (
            .O(N__4042),
            .I(N__4039));
    Sp12to4 I__438 (
            .O(N__4039),
            .I(N__4036));
    Span12Mux_h I__437 (
            .O(N__4036),
            .I(N__4033));
    Span12Mux_v I__436 (
            .O(N__4033),
            .I(N__4030));
    Odrv12 I__435 (
            .O(N__4030),
            .I(SIZ_c_1));
    InMux I__434 (
            .O(N__4027),
            .I(N__4024));
    LocalMux I__433 (
            .O(N__4024),
            .I(N__4019));
    InMux I__432 (
            .O(N__4023),
            .I(N__4016));
    InMux I__431 (
            .O(N__4022),
            .I(N__4013));
    Span4Mux_v I__430 (
            .O(N__4019),
            .I(N__4006));
    LocalMux I__429 (
            .O(N__4016),
            .I(N__4006));
    LocalMux I__428 (
            .O(N__4013),
            .I(N__4006));
    Sp12to4 I__427 (
            .O(N__4006),
            .I(N__4003));
    Span12Mux_v I__426 (
            .O(N__4003),
            .I(N__4000));
    Odrv12 I__425 (
            .O(N__4000),
            .I(SIZ_c_0));
    InMux I__424 (
            .O(N__3997),
            .I(N__3985));
    InMux I__423 (
            .O(N__3996),
            .I(N__3985));
    InMux I__422 (
            .O(N__3995),
            .I(N__3985));
    InMux I__421 (
            .O(N__3994),
            .I(N__3985));
    LocalMux I__420 (
            .O(N__3985),
            .I(\U712_BYTE_ENABLE.N_270 ));
    IoInMux I__419 (
            .O(N__3982),
            .I(N__3979));
    LocalMux I__418 (
            .O(N__3979),
            .I(N__3975));
    IoInMux I__417 (
            .O(N__3978),
            .I(N__3972));
    Span4Mux_s0_v I__416 (
            .O(N__3975),
            .I(N__3969));
    LocalMux I__415 (
            .O(N__3972),
            .I(N__3966));
    Span4Mux_h I__414 (
            .O(N__3969),
            .I(N__3963));
    Span4Mux_s0_v I__413 (
            .O(N__3966),
            .I(N__3960));
    Sp12to4 I__412 (
            .O(N__3963),
            .I(N__3957));
    Sp12to4 I__411 (
            .O(N__3960),
            .I(N__3954));
    Span12Mux_h I__410 (
            .O(N__3957),
            .I(N__3949));
    Span12Mux_s11_h I__409 (
            .O(N__3954),
            .I(N__3949));
    Span12Mux_v I__408 (
            .O(N__3949),
            .I(N__3945));
    InMux I__407 (
            .O(N__3948),
            .I(N__3942));
    Odrv12 I__406 (
            .O(N__3945),
            .I(ASn_c));
    LocalMux I__405 (
            .O(N__3942),
            .I(ASn_c));
    CascadeMux I__404 (
            .O(N__3937),
            .I(\U712_REG_SM.N_266_cascade_ ));
    InMux I__403 (
            .O(N__3934),
            .I(N__3931));
    LocalMux I__402 (
            .O(N__3931),
            .I(\U712_REG_SM.N_215 ));
    IoInMux I__401 (
            .O(N__3928),
            .I(N__3925));
    LocalMux I__400 (
            .O(N__3925),
            .I(N__3922));
    IoSpan4Mux I__399 (
            .O(N__3922),
            .I(N__3919));
    Span4Mux_s2_h I__398 (
            .O(N__3919),
            .I(N__3916));
    Span4Mux_h I__397 (
            .O(N__3916),
            .I(N__3913));
    Span4Mux_h I__396 (
            .O(N__3913),
            .I(N__3910));
    Odrv4 I__395 (
            .O(N__3910),
            .I(N_944_i));
    IoInMux I__394 (
            .O(N__3907),
            .I(N__3904));
    LocalMux I__393 (
            .O(N__3904),
            .I(N__3901));
    Span12Mux_s5_v I__392 (
            .O(N__3901),
            .I(N__3898));
    Odrv12 I__391 (
            .O(N__3898),
            .I(VBENn_c));
    CascadeMux I__390 (
            .O(N__3895),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_cascade_ ));
    IoInMux I__389 (
            .O(N__3892),
            .I(N__3889));
    LocalMux I__388 (
            .O(N__3889),
            .I(N__3886));
    Span12Mux_s11_v I__387 (
            .O(N__3886),
            .I(N__3883));
    Odrv12 I__386 (
            .O(N__3883),
            .I(N_41_i));
    InMux I__385 (
            .O(N__3880),
            .I(N__3877));
    LocalMux I__384 (
            .O(N__3877),
            .I(N__3874));
    Odrv4 I__383 (
            .O(N__3874),
            .I(\U712_BYTE_ENABLE.N_273 ));
    IoInMux I__382 (
            .O(N__3871),
            .I(N__3868));
    LocalMux I__381 (
            .O(N__3868),
            .I(N__3865));
    Span12Mux_s8_h I__380 (
            .O(N__3865),
            .I(N__3862));
    Span12Mux_h I__379 (
            .O(N__3862),
            .I(N__3859));
    Span12Mux_v I__378 (
            .O(N__3859),
            .I(N__3856));
    Odrv12 I__377 (
            .O(N__3856),
            .I(N_43_i));
    InMux I__376 (
            .O(N__3853),
            .I(N__3850));
    LocalMux I__375 (
            .O(N__3850),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0 ));
    CascadeMux I__374 (
            .O(N__3847),
            .I(\U712_BYTE_ENABLE.N_275_cascade_ ));
    IoInMux I__373 (
            .O(N__3844),
            .I(N__3841));
    LocalMux I__372 (
            .O(N__3841),
            .I(N__3838));
    Span12Mux_s5_h I__371 (
            .O(N__3838),
            .I(N__3835));
    Span12Mux_h I__370 (
            .O(N__3835),
            .I(N__3832));
    Span12Mux_v I__369 (
            .O(N__3832),
            .I(N__3829));
    Odrv12 I__368 (
            .O(N__3829),
            .I(N_42_i));
    InMux I__367 (
            .O(N__3826),
            .I(N__3822));
    InMux I__366 (
            .O(N__3825),
            .I(N__3819));
    LocalMux I__365 (
            .O(N__3822),
            .I(\U712_REG_SM.REG_CYCLE_GOZ0 ));
    LocalMux I__364 (
            .O(N__3819),
            .I(\U712_REG_SM.REG_CYCLE_GOZ0 ));
    InMux I__363 (
            .O(N__3814),
            .I(N__3811));
    LocalMux I__362 (
            .O(N__3811),
            .I(\U712_REG_SM.UDS_OUT_2_0_a2_0_a3_0 ));
    InMux I__361 (
            .O(N__3808),
            .I(N__3805));
    LocalMux I__360 (
            .O(N__3805),
            .I(N__3801));
    IoInMux I__359 (
            .O(N__3804),
            .I(N__3798));
    Span4Mux_h I__358 (
            .O(N__3801),
            .I(N__3795));
    LocalMux I__357 (
            .O(N__3798),
            .I(N__3792));
    Span4Mux_h I__356 (
            .O(N__3795),
            .I(N__3787));
    Span4Mux_s3_h I__355 (
            .O(N__3792),
            .I(N__3787));
    Sp12to4 I__354 (
            .O(N__3787),
            .I(N__3784));
    Span12Mux_v I__353 (
            .O(N__3784),
            .I(N__3781));
    Odrv12 I__352 (
            .O(N__3781),
            .I(C1_c));
    CascadeMux I__351 (
            .O(N__3778),
            .I(\U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1_cascade_ ));
    InMux I__350 (
            .O(N__3775),
            .I(N__3769));
    InMux I__349 (
            .O(N__3774),
            .I(N__3769));
    LocalMux I__348 (
            .O(N__3769),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    InMux I__347 (
            .O(N__3766),
            .I(N__3763));
    LocalMux I__346 (
            .O(N__3763),
            .I(\U712_REG_SM.LDS_OUT_2_0_a2_0_a3_0 ));
    InMux I__345 (
            .O(N__3760),
            .I(N__3750));
    InMux I__344 (
            .O(N__3759),
            .I(N__3750));
    InMux I__343 (
            .O(N__3758),
            .I(N__3750));
    InMux I__342 (
            .O(N__3757),
            .I(N__3747));
    LocalMux I__341 (
            .O(N__3750),
            .I(N__3744));
    LocalMux I__340 (
            .O(N__3747),
            .I(\U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1 ));
    Odrv4 I__339 (
            .O(N__3744),
            .I(\U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1 ));
    IoInMux I__338 (
            .O(N__3739),
            .I(N__3736));
    LocalMux I__337 (
            .O(N__3736),
            .I(N__3733));
    Span4Mux_s2_v I__336 (
            .O(N__3733),
            .I(N__3730));
    Span4Mux_v I__335 (
            .O(N__3730),
            .I(N__3727));
    Odrv4 I__334 (
            .O(N__3727),
            .I(CLK80_OUT_i_i));
    IoInMux I__333 (
            .O(N__3724),
            .I(N__3721));
    LocalMux I__332 (
            .O(N__3721),
            .I(N__3718));
    Odrv12 I__331 (
            .O(N__3718),
            .I(CLK40_OUT_i_i));
    CascadeMux I__330 (
            .O(N__3715),
            .I(N__3712));
    InMux I__329 (
            .O(N__3712),
            .I(N__3709));
    LocalMux I__328 (
            .O(N__3709),
            .I(N__3706));
    Span4Mux_v I__327 (
            .O(N__3706),
            .I(N__3703));
    Span4Mux_h I__326 (
            .O(N__3703),
            .I(N__3700));
    Sp12to4 I__325 (
            .O(N__3700),
            .I(N__3697));
    Span12Mux_v I__324 (
            .O(N__3697),
            .I(N__3694));
    Odrv12 I__323 (
            .O(N__3694),
            .I(REGSPACEn_c));
    IoInMux I__322 (
            .O(N__3691),
            .I(N__3688));
    LocalMux I__321 (
            .O(N__3688),
            .I(N__3685));
    IoSpan4Mux I__320 (
            .O(N__3685),
            .I(N__3682));
    Span4Mux_s2_v I__319 (
            .O(N__3682),
            .I(N__3679));
    Sp12to4 I__318 (
            .O(N__3679),
            .I(N__3676));
    Span12Mux_v I__317 (
            .O(N__3676),
            .I(N__3673));
    Odrv12 I__316 (
            .O(N__3673),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__9309));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_8C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_8C_net ),
            .I(N__9307));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__9308));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__9304));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__9305));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__9306));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7771),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__3804),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__4440),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_3_1_2.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_3_1_2.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_3_1_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_3_1_2 (
            .in0(N__8788),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLK40C_obuf_RNO_LC_5_10_7.C_ON=1'b0;
    defparam CLK40C_obuf_RNO_LC_5_10_7.SEQ_MODE=4'b0000;
    defparam CLK40C_obuf_RNO_LC_5_10_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLK40C_obuf_RNO_LC_5_10_7 (
            .in0(N__8074),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDS_OUT_RNO_0_LC_6_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_RNO_0_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDS_OUT_RNO_0_LC_6_11_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_REG_SM.UDS_OUT_RNO_0_LC_6_11_4  (
            .in0(N__4985),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4134),
            .lcout(\U712_REG_SM.UDS_OUT_2_0_a2_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDS_OUT_RNO_0_LC_6_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_RNO_0_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_RNO_0_LC_6_13_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_REG_SM.LDS_OUT_RNO_0_LC_6_13_6  (
            .in0(N__4969),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4127),
            .lcout(\U712_REG_SM.LDS_OUT_2_0_a2_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_7_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_7_10_5 .LUT_INIT=16'b0000010111001101;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_7_10_5  (
            .in0(N__4620),
            .in1(N__4555),
            .in2(N__3715),
            .in3(N__3826),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8772),
            .ce(),
            .sr(N__9496));
    defparam \U712_REG_SM.C3_SYNC_2_LC_7_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_2_LC_7_11_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_2_LC_7_11_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C3_SYNC_2_LC_7_11_0  (
            .in0(N__4759),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8777),
            .ce(),
            .sr(N__9490));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_7_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_7_11_1 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_7_11_1  (
            .in0(N__3759),
            .in1(N__4191),
            .in2(_gnd_net_),
            .in3(N__4213),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8777),
            .ce(),
            .sr(N__9490));
    defparam \U712_REG_SM.C1_SYNC_2_LC_7_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_2_LC_7_11_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_2_LC_7_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_2_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4257),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8777),
            .ce(),
            .sr(N__9490));
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_7_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_7_11_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_GO_LC_7_11_3  (
            .in0(N__3758),
            .in1(N__4556),
            .in2(N__4471),
            .in3(N__3825),
            .lcout(\U712_REG_SM.REG_CYCLE_GOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8777),
            .ce(),
            .sr(N__9490));
    defparam \U712_REG_SM.UDS_OUT_LC_7_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.UDS_OUT_LC_7_11_4 .LUT_INIT=16'b1111000001110111;
    LogicCell40 \U712_REG_SM.UDS_OUT_LC_7_11_4  (
            .in0(N__4023),
            .in1(N__3814),
            .in2(N__5019),
            .in3(N__3760),
            .lcout(\U712_REG_SM.UDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8777),
            .ce(),
            .sr(N__9490));
    defparam \U712_REG_SM.C1_SYNC_1_LC_7_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_7_11_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_7_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4857),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8777),
            .ce(),
            .sr(N__9490));
    defparam \U712_REG_SM.C1_SYNC_0_LC_7_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_7_11_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_7_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3808),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8777),
            .ce(),
            .sr(N__9490));
    defparam \U712_REG_SM.C1_SYNC_RNITQLC2_1_LC_7_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNITQLC2_1_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNITQLC2_1_LC_7_12_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNITQLC2_1_LC_7_12_4  (
            .in0(N__4273),
            .in1(N__4254),
            .in2(N__4853),
            .in3(N__4501),
            .lcout(\U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1 ),
            .ltout(\U712_REG_SM.C1_SYNC_RNITQLC2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_7_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_7_12_5 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_7_12_5  (
            .in0(N__4467),
            .in1(N__4561),
            .in2(N__3778),
            .in3(N__3775),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8780),
            .ce(),
            .sr(N__9483));
    defparam \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_7_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_7_12_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_7_12_6  (
            .in0(N__3774),
            .in1(N__4776),
            .in2(_gnd_net_),
            .in3(N__4757),
            .lcout(\U712_REG_SM.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_7_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_7_12_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(N__4399),
            .in2(_gnd_net_),
            .in3(N__4312),
            .lcout(\U712_REG_SM.N_201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDS_OUT_LC_7_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.LDS_OUT_LC_7_13_5 .LUT_INIT=16'b1111000001110111;
    LogicCell40 \U712_REG_SM.LDS_OUT_LC_7_13_5  (
            .in0(N__3766),
            .in1(N__4022),
            .in2(N__4378),
            .in3(N__3757),
            .lcout(\U712_REG_SM.LDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8784),
            .ce(),
            .sr(N__9472));
    defparam TACKn_obuft_RNO_LC_7_16_1.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_7_16_1.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_7_16_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 TACKn_obuft_RNO_LC_7_16_1 (
            .in0(N__5728),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_944_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_0_a3_LC_8_6_6 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_0_a3_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_0_a3_LC_8_6_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_0_a3_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(N__8420),
            .in2(_gnd_net_),
            .in3(N__7683),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_LC_8_8_0 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_LC_8_8_0  (
            .in0(N__4095),
            .in1(N__4143),
            .in2(N__4066),
            .in3(N__8389),
            .lcout(\U712_BYTE_ENABLE.N_273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_0_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_0_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_0_LC_8_8_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_0_LC_8_8_1  (
            .in0(N__5874),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7733),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0 ),
            .ltout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_41_i_LC_8_8_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_41_i_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_41_i_LC_8_8_2 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_41_i_LC_8_8_2  (
            .in0(N__4072),
            .in1(N__3994),
            .in2(N__3895),
            .in3(N__5115),
            .lcout(N_41_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_43_i_LC_8_8_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_43_i_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_43_i_LC_8_8_3 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \U712_BYTE_ENABLE.N_43_i_LC_8_8_3  (
            .in0(N__3996),
            .in1(N__3880),
            .in2(N__5119),
            .in3(N__4338),
            .lcout(N_43_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_LC_8_8_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_LC_8_8_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a3_LC_8_8_4  (
            .in0(N__4094),
            .in1(N__4142),
            .in2(_gnd_net_),
            .in3(N__8388),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_275_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_42_i_LC_8_8_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_42_i_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_42_i_LC_8_8_5 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_42_i_LC_8_8_5  (
            .in0(N__3995),
            .in1(N__3853),
            .in2(N__3847),
            .in3(N__5154),
            .lcout(N_42_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_0_LC_8_8_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_0_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_0_LC_8_8_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_0_LC_8_8_6  (
            .in0(N__4096),
            .in1(N__4144),
            .in2(_gnd_net_),
            .in3(N__8390),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_271_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_44_i_LC_8_8_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_44_i_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_44_i_LC_8_8_7 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \U712_BYTE_ENABLE.N_44_i_LC_8_8_7  (
            .in0(N__3997),
            .in1(N__4339),
            .in2(N__4168),
            .in3(N__5155),
            .lcout(N_44_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_LC_8_9_0 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_LC_8_9_0  (
            .in0(N__4126),
            .in1(N__4093),
            .in2(N__8419),
            .in3(N__4055),
            .lcout(\U712_BYTE_ENABLE.N_277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_8_9_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_8_9_3 .LUT_INIT=16'b1100000000001100;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__8387),
            .in2(N__4062),
            .in3(N__4027),
            .lcout(\U712_BYTE_ENABLE.N_270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_8_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_8_10_2 .LUT_INIT=16'b1111001000000010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_8_10_2  (
            .in0(N__5310),
            .in1(N__5293),
            .in2(N__7407),
            .in3(N__7374),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8768),
            .ce(),
            .sr(N__9491));
    defparam \U712_REG_SM.REGENn_1_LC_8_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_1_LC_8_10_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_1_LC_8_10_4 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \U712_REG_SM.REGENn_1_LC_8_10_4  (
            .in0(N__4531),
            .in1(N__3948),
            .in2(N__4515),
            .in3(N__4222),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8768),
            .ce(),
            .sr(N__9491));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_8_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_8_10_6 .LUT_INIT=16'b0111001000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_8_10_6  (
            .in0(N__4192),
            .in1(N__4209),
            .in2(N__5314),
            .in3(N__5292),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8768),
            .ce(),
            .sr(N__9491));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_8_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_8_11_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_8_11_0  (
            .in0(N__4256),
            .in1(N__4500),
            .in2(N__4855),
            .in3(N__4288),
            .lcout(),
            .ltout(\U712_REG_SM.N_266_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_8_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_8_11_1 .LUT_INIT=16'b0000011100000010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_8_11_1  (
            .in0(N__7336),
            .in1(N__3934),
            .in2(N__3937),
            .in3(N__4300),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8773),
            .ce(),
            .sr(N__9484));
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_8_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_8_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_8_11_2  (
            .in0(N__4255),
            .in1(N__4499),
            .in2(N__4854),
            .in3(N__4287),
            .lcout(\U712_REG_SM.N_215 ),
            .ltout(\U712_REG_SM.N_215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_8_11_3 .LUT_INIT=16'b1010000011100000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_8_11_3  (
            .in0(N__7337),
            .in1(N__7403),
            .in2(N__4318),
            .in3(N__7373),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8773),
            .ce(),
            .sr(N__9484));
    defparam \U712_REG_SM.C3_SYNC_1_LC_8_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_8_11_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_8_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4405),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8773),
            .ce(),
            .sr(N__9484));
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_8_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_8_11_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__4775),
            .in2(_gnd_net_),
            .in3(N__4756),
            .lcout(\U712_REG_SM.N_200 ),
            .ltout(\U712_REG_SM.N_200_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_8_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_8_11_7 .LUT_INIT=16'b1111110011111100;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__4792),
            .in2(N__4315),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.N_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_8_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_8_12_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_8_12_0  (
            .in0(N__4311),
            .in1(N__4830),
            .in2(N__4258),
            .in3(N__4403),
            .lcout(\U712_REG_SM.N_183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_8_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_8_12_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_8_12_4  (
            .in0(N__4252),
            .in1(N__4299),
            .in2(N__4858),
            .in3(N__4286),
            .lcout(\U712_REG_SM.N_325 ),
            .ltout(\U712_REG_SM.N_325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIJS6A3_1_LC_8_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIJS6A3_1_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIJS6A3_1_LC_8_12_5 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIJS6A3_1_LC_8_12_5  (
            .in0(N__4831),
            .in1(N__4272),
            .in2(N__4261),
            .in3(N__4253),
            .lcout(\U712_REG_SM.N_198 ),
            .ltout(\U712_REG_SM.N_198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_8_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_8_12_6 .LUT_INIT=16'b0100010011110100;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_8_12_6  (
            .in0(N__4208),
            .in1(N__4190),
            .in2(N__4174),
            .in3(N__4508),
            .lcout(),
            .ltout(\U712_REG_SM.DS_EN_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_LC_8_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_8_12_7 .LUT_INIT=16'b1111110010101100;
    LogicCell40 \U712_REG_SM.DS_EN_LC_8_12_7  (
            .in0(N__4404),
            .in1(N__5039),
            .in2(N__4171),
            .in3(N__4798),
            .lcout(\U712_REG_SM.DS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8778),
            .ce(),
            .sr(N__9473));
    defparam \U712_CHIP_RAM.DBR_SYNC_2_LC_8_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_SYNC_2_LC_8_13_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBR_SYNC_2_LC_8_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DBR_SYNC_2_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4692),
            .lcout(\U712_CHIP_RAM.DBR_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8781),
            .ce(),
            .sr(N__9468));
    defparam \U712_REG_SM.DBR_SYNC_1_LC_8_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_8_13_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_8_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_1_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5061),
            .lcout(U712_REG_SM_DBR_SYNC_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8781),
            .ce(),
            .sr(N__9468));
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_13_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4441),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8781),
            .ce(),
            .sr(N__9468));
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_14_6 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_14_6  (
            .in0(N__5046),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4377),
            .lcout(U712_REG_SM_un1_LDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_0_LC_9_8_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_0_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_0_LC_9_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_0_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__7732),
            .in2(_gnd_net_),
            .in3(N__5873),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_9_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_9_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__4906),
            .in2(_gnd_net_),
            .in3(N__4330),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__9303),
            .ce(),
            .sr(N__5323));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_9_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_9_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__5383),
            .in2(_gnd_net_),
            .in3(N__4327),
            .lcout(\U712_CHIP_RAM.REFRESH5lto1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__9303),
            .ce(),
            .sr(N__5323));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_9_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__4894),
            .in2(_gnd_net_),
            .in3(N__4324),
            .lcout(\U712_CHIP_RAM.REFRESH5lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__9303),
            .ce(),
            .sr(N__5323));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_9_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_9_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__4734),
            .in2(_gnd_net_),
            .in3(N__4321),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__9303),
            .ce(),
            .sr(N__5323));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_9_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__4881),
            .in2(_gnd_net_),
            .in3(N__4633),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__9303),
            .ce(),
            .sr(N__5323));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_9_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_9_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__5181),
            .in2(_gnd_net_),
            .in3(N__4630),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__9303),
            .ce(),
            .sr(N__5323));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_9_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_9_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__5196),
            .in2(_gnd_net_),
            .in3(N__4627),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__9303),
            .ce(),
            .sr(N__5323));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_9_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__4716),
            .in2(_gnd_net_),
            .in3(N__4624),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9303),
            .ce(),
            .sr(N__5323));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_10_0 .LUT_INIT=16'b0101011100000011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_10_0  (
            .in0(N__8330),
            .in1(N__4621),
            .in2(N__4585),
            .in3(N__4665),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8764),
            .ce(),
            .sr(N__9485));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_10_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_9_10_2 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_9_10_2  (
            .in0(N__4560),
            .in1(N__4530),
            .in2(N__4466),
            .in3(N__4516),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8764),
            .ce(),
            .sr(N__9485));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_10_4 .LUT_INIT=16'b0100111011001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_9_10_4  (
            .in0(N__5506),
            .in1(N__6066),
            .in2(N__4867),
            .in3(N__4648),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8764),
            .ce(),
            .sr(N__9485));
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_10_5 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_10_5  (
            .in0(N__4696),
            .in1(N__7369),
            .in2(_gnd_net_),
            .in3(N__5062),
            .lcout(\U712_REG_SM.N_209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_11_0  (
            .in0(N__7537),
            .in1(N__7047),
            .in2(N__6016),
            .in3(N__6634),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8769),
            .ce(N__5458),
            .sr(N__9474));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_11_3  (
            .in0(N__4986),
            .in1(N__5267),
            .in2(_gnd_net_),
            .in3(N__6678),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_9_11_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_1_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__4987),
            .in2(_gnd_net_),
            .in3(N__4856),
            .lcout(\U712_REG_SM.N_265 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_9_11_7 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_9_11_7  (
            .in0(N__4791),
            .in1(N__4780),
            .in2(_gnd_net_),
            .in3(N__4758),
            .lcout(\U712_REG_SM.N_187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_9_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_9_12_0 .LUT_INIT=16'b1111001111111011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_9_12_0  (
            .in0(N__4735),
            .in1(N__5167),
            .in2(N__4720),
            .in3(N__5371),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8774),
            .ce(),
            .sr(N__9469));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_12_2 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_12_2  (
            .in0(N__6677),
            .in1(N__5073),
            .in2(N__7739),
            .in3(N__4702),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8774),
            .ce(),
            .sr(N__9469));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_3  (
            .in0(N__5074),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8774),
            .ce(),
            .sr(N__9469));
    defparam \U712_CHIP_RAM.DBR_SYNC_RNIMGL61_2_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_SYNC_RNIMGL61_2_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBR_SYNC_RNIMGL61_2_LC_9_12_4 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U712_CHIP_RAM.DBR_SYNC_RNIMGL61_2_LC_9_12_4  (
            .in0(N__4688),
            .in1(N__4672),
            .in2(_gnd_net_),
            .in3(N__4666),
            .lcout(\U712_CHIP_RAM.N_177 ),
            .ltout(\U712_CHIP_RAM.N_177_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIH3B52_LC_9_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIH3B52_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIH3B52_LC_9_12_5 .LUT_INIT=16'b1111111100000011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIH3B52_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__5427),
            .in2(N__4651),
            .in3(N__6676),
            .lcout(\U712_CHIP_RAM.N_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__5444),
            .in2(_gnd_net_),
            .in3(N__4644),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a3_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_13_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__5197),
            .in2(_gnd_net_),
            .in3(N__5182),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_9_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_9_13_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIRILU_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__5426),
            .in2(_gnd_net_),
            .in3(N__6673),
            .lcout(\U712_CHIP_RAM.N_307 ),
            .ltout(\U712_CHIP_RAM.N_307_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNI6A2O6_LC_9_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNI6A2O6_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNI6A2O6_LC_9_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNI6A2O6_LC_9_13_5  (
            .in0(N__5443),
            .in1(N__5488),
            .in2(N__5161),
            .in3(N__7218),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNI6A2O6_0_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNI6A2O6_0_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNI6A2O6_0_LC_9_13_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNI6A2O6_0_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5158),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_9_14_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_9_14_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_9_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__5145),
            .in2(_gnd_net_),
            .in3(N__5109),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8782),
            .ce(),
            .sr(N__9451));
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_9_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_9_14_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_9_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DBR_SYNC_0_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9275),
            .lcout(U712_REG_SM_DBR_SYNC_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8782),
            .ce(),
            .sr(N__9451));
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_9_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_9_15_6 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_REG_SM.UDS_OUT_RNIUP9B_LC_9_15_6  (
            .in0(N__5047),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5023),
            .lcout(U712_REG_SM_un1_UDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_i_m4_i_m2_LC_9_20_3 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_m4_i_m2_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_m4_i_m2_LC_9_20_3 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_m4_i_m2_LC_9_20_3  (
            .in0(N__4976),
            .in1(N__5268),
            .in2(_gnd_net_),
            .in3(N__7746),
            .lcout(DRDDIR_i_m4_i_m2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_8_2 .LUT_INIT=16'b0001111100111111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_8_2  (
            .in0(N__4905),
            .in1(N__4893),
            .in2(N__4882),
            .in3(N__5382),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_8_5  (
            .in0(N__5359),
            .in1(N__5344),
            .in2(_gnd_net_),
            .in3(N__8546),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_8_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_8_6  (
            .in0(N__8547),
            .in1(N__8400),
            .in2(N__5326),
            .in3(N__8200),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_9_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_9_7  (
            .in0(N__6235),
            .in1(N__9025),
            .in2(N__6203),
            .in3(N__8545),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_10_10_1 .LUT_INIT=16'b1010110010101110;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_10_10_1  (
            .in0(N__5309),
            .in1(N__7670),
            .in2(N__7348),
            .in3(N__5291),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8761),
            .ce(),
            .sr(N__9475));
    defparam \U712_CHIP_RAM.DBDIR_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_10_10_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_10_10_2 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_10_10_2  (
            .in0(N__5278),
            .in1(N__5217),
            .in2(_gnd_net_),
            .in3(N__5910),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8761),
            .ce(),
            .sr(N__9475));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7MG83_3_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7MG83_3_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7MG83_3_LC_10_11_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI7MG83_3_LC_10_11_0  (
            .in0(N__6885),
            .in1(N__7524),
            .in2(N__7977),
            .in3(N__6001),
            .lcout(\U712_CHIP_RAM.N_323 ),
            .ltout(\U712_CHIP_RAM.N_323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISS7R7_3_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISS7R7_3_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISS7R7_3_LC_10_11_1 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNISS7R7_3_LC_10_11_1  (
            .in0(N__6002),
            .in1(N__5203),
            .in2(N__5206),
            .in3(N__5446),
            .lcout(\U712_CHIP_RAM.N_238 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_10_11_2 .LUT_INIT=16'b1100000000001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_10_11_2  (
            .in0(N__7041),
            .in1(N__7523),
            .in2(N__6898),
            .in3(N__7960),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_4_0_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_4_0_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_4_0_LC_10_11_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_4_0_LC_10_11_3  (
            .in0(N__7961),
            .in1(N__7042),
            .in2(N__6900),
            .in3(N__6062),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a3_3_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_11_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_11_4  (
            .in0(N__5445),
            .in1(N__6003),
            .in2(N__5467),
            .in3(N__7525),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_11_5 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_11_5  (
            .in0(N__6004),
            .in1(N__6595),
            .in2(N__5464),
            .in3(N__5518),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_188_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_11_6 .LUT_INIT=16'b1110111100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_11_6  (
            .in0(N__5404),
            .in1(N__5398),
            .in2(N__5461),
            .in3(N__6192),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8765),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_12_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(N__9524),
            .in2(_gnd_net_),
            .in3(N__5473),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_12_1  (
            .in0(N__7842),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7137),
            .lcout(\U712_CHIP_RAM.N_306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIM32A1_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIM32A1_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIM32A1_LC_10_12_2 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIM32A1_LC_10_12_2  (
            .in0(N__7138),
            .in1(N__5428),
            .in2(_gnd_net_),
            .in3(N__6675),
            .lcout(\U712_CHIP_RAM.N_221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIRGPAB_LC_10_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIRGPAB_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIRGPAB_LC_10_12_3 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIRGPAB_LC_10_12_3  (
            .in0(N__7843),
            .in1(N__7139),
            .in2(N__6582),
            .in3(N__5410),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIND16J_LC_10_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIND16J_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIND16J_LC_10_12_4 .LUT_INIT=16'b0000001100000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIND16J_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(N__5397),
            .in2(N__5386),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_12_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_12_5  (
            .in0(_gnd_net_),
            .in1(N__5524),
            .in2(_gnd_net_),
            .in3(N__7140),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_12_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_12_6  (
            .in0(N__7051),
            .in1(N__7841),
            .in2(N__7897),
            .in3(N__6889),
            .lcout(\U712_CHIP_RAM.N_240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_12_7 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_10_12_7  (
            .in0(N__7526),
            .in1(N__7050),
            .in2(N__6899),
            .in3(N__5991),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_13_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_13_0  (
            .in0(N__7845),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6129),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_13_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_13_1  (
            .in0(N__5541),
            .in1(N__5556),
            .in2(N__5578),
            .in3(N__5739),
            .lcout(\U712_CHIP_RAM.N_10 ),
            .ltout(\U712_CHIP_RAM.N_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_1_LC_10_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_1_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_1_LC_10_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_1_LC_10_13_2  (
            .in0(N__7503),
            .in1(N__7028),
            .in2(N__5512),
            .in3(N__6621),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER16 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_13_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5509),
            .in3(N__7157),
            .lcout(\U712_CHIP_RAM.N_328 ),
            .ltout(\U712_CHIP_RAM.N_328_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_13_4 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(N__5497),
            .in2(N__5491),
            .in3(N__5487),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_251_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_13_5 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_13_5  (
            .in0(N__7029),
            .in1(N__6092),
            .in2(N__5476),
            .in3(N__7883),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_13_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_13_6  (
            .in0(N__6674),
            .in1(_gnd_net_),
            .in2(N__7162),
            .in3(N__7219),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_1_esr_RNO_0_LC_10_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_1_esr_RNO_0_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_1_esr_RNO_0_LC_10_13_7 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_1_esr_RNO_0_LC_10_13_7  (
            .in0(N__7030),
            .in1(N__6091),
            .in2(N__5593),
            .in3(N__7884),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_14_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__7049),
            .in2(_gnd_net_),
            .in3(N__5590),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_14_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_14_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_14_1  (
            .in0(N__7271),
            .in1(N__7516),
            .in2(_gnd_net_),
            .in3(N__5587),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__8779),
            .ce(N__7183),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_10_14_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_10_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__6893),
            .in2(_gnd_net_),
            .in3(N__5584),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_14_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_14_3  (
            .in0(N__7272),
            .in1(N__7959),
            .in2(_gnd_net_),
            .in3(N__5581),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__8779),
            .ce(N__7183),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_14_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_14_4  (
            .in0(N__7266),
            .in1(N__5574),
            .in2(_gnd_net_),
            .in3(N__5560),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__8779),
            .ce(N__7183),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_14_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_14_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_14_5  (
            .in0(N__7273),
            .in1(N__5557),
            .in2(_gnd_net_),
            .in3(N__5545),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__8779),
            .ce(N__7183),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_14_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_14_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_14_6  (
            .in0(N__7267),
            .in1(N__5542),
            .in2(_gnd_net_),
            .in3(N__5530),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__8779),
            .ce(N__7183),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_14_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_14_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_14_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_14_7  (
            .in0(N__5740),
            .in1(N__7268),
            .in2(_gnd_net_),
            .in3(N__5527),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8779),
            .ce(N__7183),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_10_15_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_10_15_7 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_10_15_7 .LUT_INIT=16'b1111111101011111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_10_15_7  (
            .in0(N__8110),
            .in1(_gnd_net_),
            .in2(N__7849),
            .in3(N__8140),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8783),
            .ce(N__6451),
            .sr(N__9445));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_6_7  (
            .in0(N__5716),
            .in1(N__5695),
            .in2(_gnd_net_),
            .in3(N__8528),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_7_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_7_2  (
            .in0(N__8423),
            .in1(N__8548),
            .in2(N__5674),
            .in3(N__9151),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_8_4 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_11_8_4  (
            .in0(N__8909),
            .in1(N__7600),
            .in2(N__8849),
            .in3(N__5665),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8754),
            .ce(N__8664),
            .sr(N__9486));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_11_8_7 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_11_8_7  (
            .in0(N__8910),
            .in1(N__8840),
            .in2(N__7612),
            .in3(N__5830),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8754),
            .ce(N__8664),
            .sr(N__9486));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_9_0 .LUT_INIT=16'b0000011000000111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_9_0  (
            .in0(N__8523),
            .in1(N__9026),
            .in2(N__6245),
            .in3(N__6196),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_CMA30_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_9_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5632),
            .in3(N__9526),
            .lcout(\U712_CHIP_RAM.un1_CMA30_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_9_3  (
            .in0(N__5629),
            .in1(N__5611),
            .in2(_gnd_net_),
            .in3(N__8526),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_9_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_9_4  (
            .in0(N__8527),
            .in1(N__8417),
            .in2(N__5833),
            .in3(N__9598),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_9_5  (
            .in0(N__5824),
            .in1(N__5803),
            .in2(_gnd_net_),
            .in3(N__8525),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_9_7  (
            .in0(N__5785),
            .in1(N__5767),
            .in2(_gnd_net_),
            .in3(N__8524),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_2_LC_11_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_2_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_2_LC_11_10_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_2_LC_11_10_1  (
            .in0(N__9020),
            .in1(N__8499),
            .in2(_gnd_net_),
            .in3(N__6185),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_2_LC_11_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_2_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_2_LC_11_10_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_2_LC_11_10_5  (
            .in0(N__9021),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6186),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9MVM2_1_LC_11_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9MVM2_1_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9MVM2_1_LC_11_11_0 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9MVM2_1_LC_11_11_0  (
            .in0(N__7135),
            .in1(N__7535),
            .in2(N__6897),
            .in3(N__7441),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_RNI9MVM2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_11_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_11_11_1 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_11_11_1  (
            .in0(N__5752),
            .in1(N__7044),
            .in2(N__7161),
            .in3(N__6630),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_11_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_11_11_2 .LUT_INIT=16'b1111100011110010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_11_11_2  (
            .in0(N__7045),
            .in1(N__7978),
            .in2(N__5746),
            .in3(N__6880),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_101_i_a2_0_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_11_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_11_11_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5743),
            .in3(N__5925),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8762),
            .ce(N__6118),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_11_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_11_11_4 .LUT_INIT=16'b1111010011110110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_11_11_4  (
            .in0(N__7046),
            .in1(N__7979),
            .in2(N__6012),
            .in3(N__6879),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_66_0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_11_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_11_5  (
            .in0(N__6881),
            .in1(N__5917),
            .in2(N__5929),
            .in3(N__5926),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8762),
            .ce(N__6118),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_11_6 .LUT_INIT=16'b1001100111011101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_11_6  (
            .in0(N__7043),
            .in1(N__7151),
            .in2(_gnd_net_),
            .in3(N__7534),
            .lcout(\U712_CHIP_RAM.N_222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_11_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_11_12_0 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_11_12_0  (
            .in0(N__7896),
            .in1(N__6992),
            .in2(N__5911),
            .in3(N__6093),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_11_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_11_12_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_11_12_1 .LUT_INIT=16'b1010110011111100;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_11_12_1  (
            .in0(N__6993),
            .in1(N__5856),
            .in2(N__5893),
            .in3(N__7549),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8766),
            .ce(),
            .sr(N__9452));
    defparam \U712_CHIP_RAM.DMA_CYCLE_1_esr_RNO_LC_11_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_1_esr_RNO_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_1_esr_RNO_LC_11_12_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_1_esr_RNO_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__9523),
            .in2(_gnd_net_),
            .in3(N__5845),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_3_LC_11_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_3_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_3_LC_11_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_0_3_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(N__7965),
            .in2(_gnd_net_),
            .in3(N__6844),
            .lcout(\U712_CHIP_RAM.N_305 ),
            .ltout(\U712_CHIP_RAM.N_305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_11_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_11_12_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_11_12_5  (
            .in0(N__6991),
            .in1(N__5989),
            .in2(N__5839),
            .in3(N__7527),
            .lcout(\U712_CHIP_RAM.N_254_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_13_0 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_13_0  (
            .in0(N__7440),
            .in1(N__7001),
            .in2(_gnd_net_),
            .in3(N__6622),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_13_1 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_13_1  (
            .in0(N__7002),
            .in1(N__7131),
            .in2(N__5836),
            .in3(N__7522),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_13_2 .LUT_INIT=16'b1111110011111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_13_2  (
            .in0(N__7007),
            .in1(N__6433),
            .in2(N__6133),
            .in3(N__6130),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8770),
            .ce(N__6117),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_11_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_11_13_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__7937),
            .in2(_gnd_net_),
            .in3(N__6828),
            .lcout(\U712_CHIP_RAM.N_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_11_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_11_13_4 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_11_13_4  (
            .in0(N__7130),
            .in1(N__5990),
            .in2(_gnd_net_),
            .in3(N__7509),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_11_14_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_11_14_0 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_11_14_0  (
            .in0(N__6097),
            .in1(N__7000),
            .in2(N__5938),
            .in3(N__7892),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_11_14_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_11_14_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_11_14_1 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_11_14_1  (
            .in0(N__6030),
            .in1(N__7003),
            .in2(N__6073),
            .in3(N__6070),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8775),
            .ce(),
            .sr(N__9446));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_11_14_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_11_14_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_0_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__7156),
            .in2(_gnd_net_),
            .in3(N__6583),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOF0DC_LC_11_14_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOF0DC_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOF0DC_LC_11_14_3 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOF0DC_LC_11_14_3  (
            .in0(N__7844),
            .in1(N__7858),
            .in2(N__6019),
            .in3(N__7220),
            .lcout(\U712_CHIP_RAM.N_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_11_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_11_14_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_11_14_5  (
            .in0(N__7155),
            .in1(N__5979),
            .in2(_gnd_net_),
            .in3(N__7504),
            .lcout(\U712_CHIP_RAM.N_312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_11_14_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_11_14_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_11_14_7  (
            .in0(N__6999),
            .in1(N__7505),
            .in2(N__6005),
            .in3(N__7063),
            .lcout(\U712_CHIP_RAM.N_260 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_15_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_15_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__7057),
            .in2(_gnd_net_),
            .in3(N__9521),
            .lcout(\U712_CYCLE_TERM.N_214_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_15_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_15_5 .LUT_INIT=16'b1111111111000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_15_5  (
            .in0(N__7048),
            .in1(N__7958),
            .in2(N__6901),
            .in3(N__6442),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_a2_2_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CRCSn_LC_12_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_12_5_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_12_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6246),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8747),
            .ce(),
            .sr(N__9495));
    defparam \U712_CHIP_RAM.WEn_LC_12_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_12_5_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_12_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6211),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8747),
            .ce(),
            .sr(N__9495));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_6_1 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_12_6_1  (
            .in0(N__8430),
            .in1(N__6364),
            .in2(N__6349),
            .in3(N__6742),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8749),
            .ce(N__8668),
            .sr(N__9489));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_6_4 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_12_6_4  (
            .in0(N__6741),
            .in1(N__6310),
            .in2(N__9337),
            .in3(N__8431),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8749),
            .ce(N__8668),
            .sr(N__9489));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_7_0 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_12_7_0  (
            .in0(N__8911),
            .in1(N__8844),
            .in2(N__8932),
            .in3(N__6496),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8750),
            .ce(N__8654),
            .sr(N__9482));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_7_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_12_7_1  (
            .in0(N__9033),
            .in1(N__6247),
            .in2(N__8572),
            .in3(N__6210),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8750),
            .ce(N__8654),
            .sr(N__9482));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_7_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_12_7_3  (
            .in0(N__8912),
            .in1(N__9226),
            .in2(N__8850),
            .in3(N__6559),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8750),
            .ce(N__8654),
            .sr(N__9482));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_3  (
            .in0(N__6532),
            .in1(N__6517),
            .in2(_gnd_net_),
            .in3(N__8562),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_8_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_8_4  (
            .in0(N__8395),
            .in1(N__8564),
            .in2(N__6499),
            .in3(N__9187),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_8_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(N__8394),
            .in2(_gnd_net_),
            .in3(N__8561),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_8_7 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_8_7  (
            .in0(N__6490),
            .in1(N__8563),
            .in2(N__7561),
            .in3(N__8396),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_9_0 .LUT_INIT=16'b0001101000001010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_9_0  (
            .in0(N__8889),
            .in1(N__8415),
            .in2(N__8570),
            .in3(N__8154),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_9_1 .LUT_INIT=16'b0011001111111011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_9_1  (
            .in0(N__8155),
            .in1(N__8554),
            .in2(N__8429),
            .in3(N__8890),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_9_4 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_9_4  (
            .in0(N__6484),
            .in1(N__8416),
            .in2(N__8571),
            .in3(N__7567),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_9_5 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(N__6478),
            .in2(N__6472),
            .in3(N__6469),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8753),
            .ce(N__8671),
            .sr(N__9467));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_12_9_7  (
            .in0(N__6691),
            .in1(N__6748),
            .in2(_gnd_net_),
            .in3(N__6754),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8753),
            .ce(N__8671),
            .sr(N__9467));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_10_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_10_0  (
            .in0(N__6775),
            .in1(N__8401),
            .in2(_gnd_net_),
            .in3(N__8188),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_316_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_10_1 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__8888),
            .in2(N__6757),
            .in3(N__8565),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_10_3 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_10_3  (
            .in0(N__6714),
            .in1(N__6731),
            .in2(N__8422),
            .in3(N__9114),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_10_7 .LUT_INIT=16'b1111011110110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_10_7  (
            .in0(N__8402),
            .in1(N__6732),
            .in2(N__6718),
            .in3(N__9115),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_1_esr_LC_12_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_1_esr_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_1_esr_LC_12_11_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_1_esr_LC_12_11_0  (
            .in0(N__7136),
            .in1(N__6685),
            .in2(_gnd_net_),
            .in3(N__7238),
            .lcout(RAMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8759),
            .ce(N__6640),
            .sr(N__9450));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_12_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_12_12_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_12_12_0  (
            .in0(N__7821),
            .in1(N__7133),
            .in2(N__7039),
            .in3(N__6626),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_0_a3_2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_12_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_12_1  (
            .in0(N__7134),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6581),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8760),
            .ce(),
            .sr(N__9448));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1_1_LC_12_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1_1_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1_1_LC_12_12_3 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1_1_LC_12_12_3  (
            .in0(N__7822),
            .in1(N__6998),
            .in2(_gnd_net_),
            .in3(N__7536),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_RNIHMND1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_12_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_12_12_5 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_12_12_5  (
            .in0(N__8418),
            .in1(N__7420),
            .in2(N__7040),
            .in3(N__7429),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8760),
            .ce(),
            .sr(N__9448));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_12_12_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_12_12_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__7311),
            .in2(_gnd_net_),
            .in3(N__7419),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_LC_12_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_12_12_7 .LUT_INIT=16'b1100110010101110;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_12_12_7  (
            .in0(N__7312),
            .in1(N__7408),
            .in2(N__7381),
            .in3(N__7344),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8760),
            .ce(),
            .sr(N__9448));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_13_0 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_13_0  (
            .in0(N__7303),
            .in1(N__7269),
            .in2(N__7239),
            .in3(N__7294),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8763),
            .ce(N__7182),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_12_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_12_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_12_13_2 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_12_13_2  (
            .in0(N__7282),
            .in1(N__7270),
            .in2(N__7240),
            .in3(N__7195),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8763),
            .ce(N__7182),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_12_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_12_13_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_2_LC_12_13_3  (
            .in0(N__7132),
            .in1(N__7980),
            .in2(_gnd_net_),
            .in3(N__6869),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_14_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_14_0 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_14_0  (
            .in0(N__7823),
            .in1(N__8099),
            .in2(N__9049),
            .in3(N__8136),
            .lcout(\U712_CYCLE_TERM.N_214_i_0_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_12_14_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_12_14_1 .LUT_INIT=16'b1000001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_12_14_1  (
            .in0(N__6994),
            .in1(N__6845),
            .in2(N__7981),
            .in3(N__7885),
            .lcout(\U712_CHIP_RAM.N_243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_0.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_0.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_17_0 (
            .in0(N__7824),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_12_17_3 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_12_17_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_12_17_3  (
            .in0(N__7728),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7687),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_7_3 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_13_7_3  (
            .in0(N__8919),
            .in1(N__8845),
            .in2(N__8242),
            .in3(N__7633),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8752),
            .ce(N__8669),
            .sr(N__9492));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8227),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9093),
            .ce(N__9692),
            .sr(N__9487));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_6  (
            .in0(N__7591),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9093),
            .ce(N__9692),
            .sr(N__9487));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7590),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__9588),
            .sr(N__9476));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_7  (
            .in0(N__8182),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__9588),
            .sr(N__9476));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8275),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__9585),
            .sr(N__9470));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8226),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__9585),
            .sr(N__9470));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_10_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_10_4  (
            .in0(N__8949),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__9585),
            .sr(N__9470));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8178),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9090),
            .ce(N__9667),
            .sr(N__9460));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_13_12_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_13_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_13_12_4 .LUT_INIT=16'b1110000011101100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_13_12_4  (
            .in0(N__8062),
            .in1(N__8103),
            .in2(N__8035),
            .in3(N__8135),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8767),
            .ce(),
            .sr(N__9453));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_13_13_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_13_13_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_13_13_0  (
            .in0(N__8030),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8064),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8771),
            .ce(),
            .sr(N__9449));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_13_13_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_13_13_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__9062),
            .in2(_gnd_net_),
            .in3(N__8082),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_13_13_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_13_13_2 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_13_13_2 .LUT_INIT=16'b0101010001000100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_13_13_2  (
            .in0(N__8029),
            .in1(N__9048),
            .in2(N__8143),
            .in3(N__8134),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8771),
            .ce(),
            .sr(N__9449));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_13_13_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_13_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8083),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8771),
            .ce(),
            .sr(N__9449));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_13_13_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_13_13_5 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_13_13_5 .LUT_INIT=16'b1111111110110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_13_13_5  (
            .in0(N__8063),
            .in1(N__8031),
            .in2(N__7998),
            .in3(N__9063),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8771),
            .ce(),
            .sr(N__9449));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_13_14_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_13_14_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_13_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9064),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8776),
            .ce(),
            .sr(N__9447));
    defparam \U712_CHIP_RAM.RASn_LC_14_3_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_14_3_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_14_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_14_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9034),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8748),
            .ce(),
            .sr(N__9502));
    defparam \U712_CHIP_RAM.CASn_LC_14_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_14_5_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_14_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_14_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8569),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8751),
            .ce(),
            .sr(N__9501));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8956),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9094),
            .ce(N__9691),
            .sr(N__9497));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_8_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_14_8_3  (
            .in0(N__8920),
            .in1(N__9217),
            .in2(N__8851),
            .in3(N__8281),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8758),
            .ce(N__8670),
            .sr(N__9493));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_9_4  (
            .in0(N__8608),
            .in1(N__8590),
            .in2(_gnd_net_),
            .in3(N__8552),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_9_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_9_5  (
            .in0(N__8553),
            .in1(N__8421),
            .in2(N__8284),
            .in3(N__9322),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8268),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9091),
            .ce(N__9678),
            .sr(N__9477));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9175),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9091),
            .ce(N__9678),
            .sr(N__9477));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9139),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__9578),
            .sr(N__9471));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_8_LC_14_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_8_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_8_LC_14_12_3 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_8_LC_14_12_3  (
            .in0(N__9525),
            .in1(N__9277),
            .in2(_gnd_net_),
            .in3(N__9313),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_ctle_8_LC_14_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_ctle_8_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_ctle_8_LC_14_13_2 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_ctle_8_LC_14_13_2  (
            .in0(N__9522),
            .in1(N__9276),
            .in2(_gnd_net_),
            .in3(N__9100),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9211),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9096),
            .ce(N__9694),
            .sr(N__9500));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9631),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9095),
            .ce(N__9693),
            .sr(N__9498));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9204),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__9587),
            .sr(N__9494));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_8_LC_15_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_8_LC_15_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_8_LC_15_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_8_LC_15_10_1  (
            .in0(N__9174),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_8C_net ),
            .ce(N__9586),
            .sr(N__9488));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_11_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_11_3  (
            .in0(N__9138),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9092),
            .ce(N__9668),
            .sr(N__9478));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_16_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_16_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_16_9_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_16_9_3  (
            .in0(N__9630),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__9589),
            .sr(N__9499));
endmodule // U712_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 18 2024 20:38:43

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RAMENn : out std_logic;
    RASn : out std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__10019\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_OUT_i_i\ : std_logic;
signal \N_882_i\ : std_logic;
signal \CLK40_OUT_i_i\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \CLK40_OUT_i\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \N_46_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_383\ : std_logic;
signal \U712_BYTE_ENABLE.N_379\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_0_cascade_\ : std_logic;
signal \N_48_i\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \U712_BYTE_ENABLE.N_381\ : std_logic;
signal \U712_BYTE_ENABLE.N_376_cascade_\ : std_logic;
signal \N_47_i\ : std_logic;
signal \A_c_1\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_376\ : std_logic;
signal \U712_BYTE_ENABLE.N_377_cascade_\ : std_logic;
signal \N_49_i\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_2_1_0\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0Z0Z_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_295\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.N_338\ : std_logic;
signal \U712_REG_SM.N_292\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_2_0\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_e_1_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_296\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_tz_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_1\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_139\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_1\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6\ : std_logic;
signal \U712_REG_SM.N_492\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c4\ : std_logic;
signal \U712_REG_SM.N_273_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_273\ : std_logic;
signal \U712_REG_SM.N_420\ : std_logic;
signal \U712_REG_SM.N_491\ : std_logic;
signal \U712_REG_SM.N_420_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \U712_REG_SM.N_281\ : std_logic;
signal \U712_REG_SM.N_281_cascade_\ : std_logic;
signal \U712_REG_SM.N_300\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_274\ : std_logic;
signal \U712_REG_SM.N_282\ : std_logic;
signal \U712_REG_SM.N_274_cascade_\ : std_logic;
signal \U712_REG_SM.N_297\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_308\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.N_310\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST_cascade_\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_340_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_278\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_1_0\ : std_logic;
signal \U712_CHIP_RAM.N_417_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_427\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.N_298_i_0_en_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_298_i_0_en_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_267_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_204_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_204_0_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.DS_EN_RNOZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_210\ : std_logic;
signal \U712_REG_SM.N_355\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_5\ : std_logic;
signal \U712_REG_SM.N_279\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_301\ : std_logic;
signal \U712_REG_SM.N_302_cascade_\ : std_logic;
signal \U712_REG_SM.LDS_OUT_2_0_a2_0_a2Z0Z_0\ : std_logic;
signal \A_c_0\ : std_logic;
signal \U712_REG_SM.N_302\ : std_logic;
signal \U712_REG_SM.LDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_LDSn_i\ : std_logic;
signal \U712_REG_SM.DS_ENZ0\ : std_logic;
signal \U712_REG_SM.UDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_UDSn_i\ : std_logic;
signal \RnW_c\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \N_208\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5_cascade_\ : std_logic;
signal \A_c_7\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.N_307\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.N_311\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.N_312\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0\ : std_logic;
signal \U712_CHIP_RAM.N_306\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_336\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_3_1\ : std_logic;
signal \U712_CHIP_RAM.N_369\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c2\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_START_RNIQU7BEZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_3\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_275_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_423_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_265\ : std_logic;
signal \U712_CHIP_RAM.N_303\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a3_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGURED_e_1\ : std_logic;
signal \U712_CHIP_RAM.N_276_i\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_428\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_275\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_0_a2_0_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_375_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_263\ : std_logic;
signal \U712_CHIP_RAM.N_267\ : std_logic;
signal \U712_CHIP_RAM.N_270\ : std_logic;
signal \U712_CHIP_RAM.N_289\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \RASn_c\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.N_313_cascade_\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.N_309\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i_0\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \A_c_20\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_7_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_148\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    CLK_EN <= \CLK_EN_wire\;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    LDSn <= \LDSn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_OUT_i\,
            REFERENCECLK => \N__3610\,
            RESETB => \N__5941\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_OUT\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10019\,
            DIN => \N__10018\,
            DOUT => \N__10017\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10019\,
            PADOUT => \N__10018\,
            PADIN => \N__10017\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8098\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10010\,
            DIN => \N__10009\,
            DOUT => \N__10008\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10010\,
            PADOUT => \N__10009\,
            PADIN => \N__10008\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10001\,
            DIN => \N__10000\,
            DOUT => \N__9999\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10001\,
            PADOUT => \N__10000\,
            PADIN => \N__9999\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8794\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9992\,
            DIN => \N__9991\,
            DOUT => \N__9990\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9992\,
            PADOUT => \N__9991\,
            PADIN => \N__9990\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5956\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9983\,
            DIN => \N__9982\,
            DOUT => \N__9981\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9983\,
            PADOUT => \N__9982\,
            PADIN => \N__9981\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9974\,
            DIN => \N__9973\,
            DOUT => \N__9972\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9974\,
            PADOUT => \N__9973\,
            PADIN => \N__9972\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9965\,
            DIN => \N__9964\,
            DOUT => \N__9963\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9965\,
            PADOUT => \N__9964\,
            PADIN => \N__9963\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9956\,
            DIN => \N__9955\,
            DOUT => \N__9954\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9956\,
            PADOUT => \N__9955\,
            PADIN => \N__9954\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9947\,
            DIN => \N__9946\,
            DOUT => \N__9945\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9947\,
            PADOUT => \N__9946\,
            PADIN => \N__9945\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9938\,
            DIN => \N__9937\,
            DOUT => \N__9936\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9938\,
            PADOUT => \N__9937\,
            PADIN => \N__9936\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9929\,
            DIN => \N__9928\,
            DOUT => \N__9927\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9929\,
            PADOUT => \N__9928\,
            PADIN => \N__9927\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7456\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9920\,
            DIN => \N__9919\,
            DOUT => \N__9918\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9920\,
            PADOUT => \N__9919\,
            PADIN => \N__9918\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4269\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9911\,
            DIN => \N__9910\,
            DOUT => \N__9909\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9911\,
            PADOUT => \N__9910\,
            PADIN => \N__9909\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9902\,
            DIN => \N__9901\,
            DOUT => \N__9900\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9902\,
            PADOUT => \N__9901\,
            PADIN => \N__9900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9893\,
            DIN => \N__9892\,
            DOUT => \N__9891\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9893\,
            PADOUT => \N__9892\,
            PADIN => \N__9891\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3622\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9884\,
            DIN => \N__9883\,
            DOUT => \N__9882\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9884\,
            PADOUT => \N__9883\,
            PADIN => \N__9882\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9875\,
            DIN => \N__9874\,
            DOUT => \N__9873\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9875\,
            PADOUT => \N__9874\,
            PADIN => \N__9873\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9866\,
            DIN => \N__9865\,
            DOUT => \N__9864\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9866\,
            PADOUT => \N__9865\,
            PADIN => \N__9864\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6241\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9857\,
            DIN => \N__9856\,
            DOUT => \N__9855\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9857\,
            PADOUT => \N__9856\,
            PADIN => \N__9855\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9848\,
            DIN => \N__9847\,
            DOUT => \N__9846\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9848\,
            PADOUT => \N__9847\,
            PADIN => \N__9846\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8740\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9839\,
            DIN => \N__9838\,
            DOUT => \N__9837\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9839\,
            PADOUT => \N__9838\,
            PADIN => \N__9837\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9830\,
            DIN => \N__9829\,
            DOUT => \N__9828\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9830\,
            PADOUT => \N__9829\,
            PADIN => \N__9828\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9821\,
            DIN => \N__9820\,
            DOUT => \N__9819\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9821\,
            PADOUT => \N__9820\,
            PADIN => \N__9819\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9812\,
            DIN => \N__9811\,
            DOUT => \N__9810\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9812\,
            PADOUT => \N__9811\,
            PADIN => \N__9810\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9803\,
            DIN => \N__9802\,
            DOUT => \N__9801\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9803\,
            PADOUT => \N__9802\,
            PADIN => \N__9801\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9794\,
            DIN => \N__9793\,
            DOUT => \N__9792\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9794\,
            PADOUT => \N__9793\,
            PADIN => \N__9792\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7825\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9785\,
            DIN => \N__9784\,
            DOUT => \N__9783\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9785\,
            PADOUT => \N__9784\,
            PADIN => \N__9783\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9776\,
            DIN => \N__9775\,
            DOUT => \N__9774\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9776\,
            PADOUT => \N__9775\,
            PADIN => \N__9774\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9767\,
            DIN => \N__9766\,
            DOUT => \N__9765\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9767\,
            PADOUT => \N__9766\,
            PADIN => \N__9765\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9758\,
            DIN => \N__9757\,
            DOUT => \N__9756\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9758\,
            PADOUT => \N__9757\,
            PADIN => \N__9756\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9749\,
            DIN => \N__9748\,
            DOUT => \N__9747\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9749\,
            PADOUT => \N__9748\,
            PADIN => \N__9747\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9740\,
            DIN => \N__9739\,
            DOUT => \N__9738\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9740\,
            PADOUT => \N__9739\,
            PADIN => \N__9738\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5824\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9731\,
            DIN => \N__9730\,
            DOUT => \N__9729\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9731\,
            PADOUT => \N__9730\,
            PADIN => \N__9729\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9722\,
            DIN => \N__9721\,
            DOUT => \N__9720\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9722\,
            PADOUT => \N__9721\,
            PADIN => \N__9720\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9713\,
            DIN => \N__9712\,
            DOUT => \N__9711\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9713\,
            PADOUT => \N__9712\,
            PADIN => \N__9711\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9704\,
            DIN => \N__9703\,
            DOUT => \N__9702\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9704\,
            PADOUT => \N__9703\,
            PADIN => \N__9702\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9695\,
            DIN => \N__9694\,
            DOUT => \N__9693\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9695\,
            PADOUT => \N__9694\,
            PADIN => \N__9693\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3721\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9686\,
            DIN => \N__9685\,
            DOUT => \N__9684\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9686\,
            PADOUT => \N__9685\,
            PADIN => \N__9684\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5503\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9677\,
            DIN => \N__9676\,
            DOUT => \N__9675\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9677\,
            PADOUT => \N__9676\,
            PADIN => \N__9675\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9668\,
            DIN => \N__9667\,
            DOUT => \N__9666\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9668\,
            PADOUT => \N__9667\,
            PADIN => \N__9666\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7516\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9659\,
            DIN => \N__9658\,
            DOUT => \N__9657\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9659\,
            PADOUT => \N__9658\,
            PADIN => \N__9657\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9650\,
            DIN => \N__9649\,
            DOUT => \N__9648\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9650\,
            PADOUT => \N__9649\,
            PADIN => \N__9648\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8200\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9641\,
            DIN => \N__9640\,
            DOUT => \N__9639\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9641\,
            PADOUT => \N__9640\,
            PADIN => \N__9639\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3757\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9632\,
            DIN => \N__9631\,
            DOUT => \N__9630\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9632\,
            PADOUT => \N__9631\,
            PADIN => \N__9630\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9623\,
            DIN => \N__9622\,
            DOUT => \N__9621\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9623\,
            PADOUT => \N__9622\,
            PADIN => \N__9621\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4231\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9614\,
            DIN => \N__9613\,
            DOUT => \N__9612\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9614\,
            PADOUT => \N__9613\,
            PADIN => \N__9612\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7246\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9605\,
            DIN => \N__9604\,
            DOUT => \N__9603\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9605\,
            PADOUT => \N__9604\,
            PADIN => \N__9603\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9596\,
            DIN => \N__9595\,
            DOUT => \N__9594\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9596\,
            PADOUT => \N__9595\,
            PADIN => \N__9594\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9587\,
            DIN => \N__9586\,
            DOUT => \N__9585\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9587\,
            PADOUT => \N__9586\,
            PADIN => \N__9585\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9578\,
            DIN => \N__9577\,
            DOUT => \N__9576\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9578\,
            PADOUT => \N__9577\,
            PADIN => \N__9576\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9569\,
            DIN => \N__9568\,
            DOUT => \N__9567\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9569\,
            PADOUT => \N__9568\,
            PADIN => \N__9567\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6283\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9560\,
            DIN => \N__9559\,
            DOUT => \N__9558\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9560\,
            PADOUT => \N__9559\,
            PADIN => \N__9558\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9551\,
            DIN => \N__9550\,
            DOUT => \N__9549\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9551\,
            PADOUT => \N__9550\,
            PADIN => \N__9549\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5095\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9542\,
            DIN => \N__9541\,
            DOUT => \N__9540\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9542\,
            PADOUT => \N__9541\,
            PADIN => \N__9540\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7612\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9533\,
            DIN => \N__9532\,
            DOUT => \N__9531\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9533\,
            PADOUT => \N__9532\,
            PADIN => \N__9531\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3844\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9524\,
            DIN => \N__9523\,
            DOUT => \N__9522\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9524\,
            PADOUT => \N__9523\,
            PADIN => \N__9522\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7360\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9515\,
            DIN => \N__9514\,
            DOUT => \N__9513\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9515\,
            PADOUT => \N__9514\,
            PADIN => \N__9513\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4227\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9506\,
            DIN => \N__9505\,
            DOUT => \N__9504\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9506\,
            PADOUT => \N__9505\,
            PADIN => \N__9504\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9497\,
            DIN => \N__9496\,
            DOUT => \N__9495\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9497\,
            PADOUT => \N__9496\,
            PADIN => \N__9495\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9488\,
            DIN => \N__9487\,
            DOUT => \N__9486\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9488\,
            PADOUT => \N__9487\,
            PADIN => \N__9486\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4093\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9479\,
            DIN => \N__9478\,
            DOUT => \N__9477\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9479\,
            PADOUT => \N__9478\,
            PADIN => \N__9477\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8437\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9470\,
            DIN => \N__9469\,
            DOUT => \N__9468\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9470\,
            PADOUT => \N__9469\,
            PADIN => \N__9468\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5992\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9461\,
            DIN => \N__9460\,
            DOUT => \N__9459\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9461\,
            PADOUT => \N__9460\,
            PADIN => \N__9459\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4168\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9452\,
            DIN => \N__9451\,
            DOUT => \N__9450\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9452\,
            PADOUT => \N__9451\,
            PADIN => \N__9450\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9443\,
            DIN => \N__9442\,
            DOUT => \N__9441\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9443\,
            PADOUT => \N__9442\,
            PADIN => \N__9441\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9434\,
            DIN => \N__9433\,
            DOUT => \N__9432\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9434\,
            PADOUT => \N__9433\,
            PADIN => \N__9432\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9425\,
            DIN => \N__9424\,
            DOUT => \N__9423\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9425\,
            PADOUT => \N__9424\,
            PADIN => \N__9423\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9416\,
            DIN => \N__9415\,
            DOUT => \N__9414\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9416\,
            PADOUT => \N__9415\,
            PADIN => \N__9414\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6292\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9407\,
            DIN => \N__9406\,
            DOUT => \N__9405\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9407\,
            PADOUT => \N__9406\,
            PADIN => \N__9405\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9398\,
            DIN => \N__9397\,
            DOUT => \N__9396\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9398\,
            PADOUT => \N__9397\,
            PADIN => \N__9396\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4009\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9389\,
            DIN => \N__9388\,
            DOUT => \N__9387\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9389\,
            PADOUT => \N__9388\,
            PADIN => \N__9387\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3742\,
            DIN0 => OPEN,
            DOUT0 => \N__3652\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9380\,
            DIN => \N__9379\,
            DOUT => \N__9378\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9380\,
            PADOUT => \N__9379\,
            PADIN => \N__9378\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5113\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9371\,
            DIN => \N__9370\,
            DOUT => \N__9369\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9371\,
            PADOUT => \N__9370\,
            PADIN => \N__9369\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9362\,
            DIN => \N__9361\,
            DOUT => \N__9360\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9362\,
            PADOUT => \N__9361\,
            PADIN => \N__9360\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9353\,
            DIN => \N__9352\,
            DOUT => \N__9351\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9353\,
            PADOUT => \N__9352\,
            PADIN => \N__9351\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7414\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9344\,
            DIN => \N__9343\,
            DOUT => \N__9342\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9344\,
            PADOUT => \N__9343\,
            PADIN => \N__9342\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9335\,
            DIN => \N__9334\,
            DOUT => \N__9333\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9335\,
            PADOUT => \N__9334\,
            PADIN => \N__9333\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9326\,
            DIN => \N__9325\,
            DOUT => \N__9324\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9326\,
            PADOUT => \N__9325\,
            PADIN => \N__9324\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9317\,
            DIN => \N__9316\,
            DOUT => \N__9315\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9317\,
            PADOUT => \N__9316\,
            PADIN => \N__9315\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9308\,
            DIN => \N__9307\,
            DOUT => \N__9306\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9308\,
            PADOUT => \N__9307\,
            PADIN => \N__9306\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6256\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9299\,
            DIN => \N__9298\,
            DOUT => \N__9297\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9299\,
            PADOUT => \N__9298\,
            PADIN => \N__9297\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6055\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2200\ : InMux
    port map (
            O => \N__9280\,
            I => \N__9277\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__9277\,
            I => \N__9273\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9276\,
            I => \N__9270\
        );

    \I__2197\ : Span4Mux_v
    port map (
            O => \N__9273\,
            I => \N__9267\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__9270\,
            I => \N__9264\
        );

    \I__2195\ : Sp12to4
    port map (
            O => \N__9267\,
            I => \N__9261\
        );

    \I__2194\ : Span12Mux_v
    port map (
            O => \N__9264\,
            I => \N__9258\
        );

    \I__2193\ : Span12Mux_h
    port map (
            O => \N__9261\,
            I => \N__9255\
        );

    \I__2192\ : Span12Mux_h
    port map (
            O => \N__9258\,
            I => \N__9252\
        );

    \I__2191\ : Odrv12
    port map (
            O => \N__9255\,
            I => \RAS0n_c\
        );

    \I__2190\ : Odrv12
    port map (
            O => \N__9252\,
            I => \RAS0n_c\
        );

    \I__2189\ : InMux
    port map (
            O => \N__9247\,
            I => \N__9243\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9246\,
            I => \N__9240\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__9243\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9240\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9232\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__9232\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9229\,
            I => \N__9226\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__9226\,
            I => \N__9207\
        );

    \I__2181\ : ClkMux
    port map (
            O => \N__9225\,
            I => \N__9097\
        );

    \I__2180\ : ClkMux
    port map (
            O => \N__9224\,
            I => \N__9097\
        );

    \I__2179\ : ClkMux
    port map (
            O => \N__9223\,
            I => \N__9097\
        );

    \I__2178\ : ClkMux
    port map (
            O => \N__9222\,
            I => \N__9097\
        );

    \I__2177\ : ClkMux
    port map (
            O => \N__9221\,
            I => \N__9097\
        );

    \I__2176\ : ClkMux
    port map (
            O => \N__9220\,
            I => \N__9097\
        );

    \I__2175\ : ClkMux
    port map (
            O => \N__9219\,
            I => \N__9097\
        );

    \I__2174\ : ClkMux
    port map (
            O => \N__9218\,
            I => \N__9097\
        );

    \I__2173\ : ClkMux
    port map (
            O => \N__9217\,
            I => \N__9097\
        );

    \I__2172\ : ClkMux
    port map (
            O => \N__9216\,
            I => \N__9097\
        );

    \I__2171\ : ClkMux
    port map (
            O => \N__9215\,
            I => \N__9097\
        );

    \I__2170\ : ClkMux
    port map (
            O => \N__9214\,
            I => \N__9097\
        );

    \I__2169\ : ClkMux
    port map (
            O => \N__9213\,
            I => \N__9097\
        );

    \I__2168\ : ClkMux
    port map (
            O => \N__9212\,
            I => \N__9097\
        );

    \I__2167\ : ClkMux
    port map (
            O => \N__9211\,
            I => \N__9097\
        );

    \I__2166\ : ClkMux
    port map (
            O => \N__9210\,
            I => \N__9097\
        );

    \I__2165\ : Glb2LocalMux
    port map (
            O => \N__9207\,
            I => \N__9097\
        );

    \I__2164\ : ClkMux
    port map (
            O => \N__9206\,
            I => \N__9097\
        );

    \I__2163\ : ClkMux
    port map (
            O => \N__9205\,
            I => \N__9097\
        );

    \I__2162\ : ClkMux
    port map (
            O => \N__9204\,
            I => \N__9097\
        );

    \I__2161\ : ClkMux
    port map (
            O => \N__9203\,
            I => \N__9097\
        );

    \I__2160\ : ClkMux
    port map (
            O => \N__9202\,
            I => \N__9097\
        );

    \I__2159\ : ClkMux
    port map (
            O => \N__9201\,
            I => \N__9097\
        );

    \I__2158\ : ClkMux
    port map (
            O => \N__9200\,
            I => \N__9097\
        );

    \I__2157\ : ClkMux
    port map (
            O => \N__9199\,
            I => \N__9097\
        );

    \I__2156\ : ClkMux
    port map (
            O => \N__9198\,
            I => \N__9097\
        );

    \I__2155\ : ClkMux
    port map (
            O => \N__9197\,
            I => \N__9097\
        );

    \I__2154\ : ClkMux
    port map (
            O => \N__9196\,
            I => \N__9097\
        );

    \I__2153\ : ClkMux
    port map (
            O => \N__9195\,
            I => \N__9097\
        );

    \I__2152\ : ClkMux
    port map (
            O => \N__9194\,
            I => \N__9097\
        );

    \I__2151\ : ClkMux
    port map (
            O => \N__9193\,
            I => \N__9097\
        );

    \I__2150\ : ClkMux
    port map (
            O => \N__9192\,
            I => \N__9097\
        );

    \I__2149\ : ClkMux
    port map (
            O => \N__9191\,
            I => \N__9097\
        );

    \I__2148\ : ClkMux
    port map (
            O => \N__9190\,
            I => \N__9097\
        );

    \I__2147\ : ClkMux
    port map (
            O => \N__9189\,
            I => \N__9097\
        );

    \I__2146\ : ClkMux
    port map (
            O => \N__9188\,
            I => \N__9097\
        );

    \I__2145\ : ClkMux
    port map (
            O => \N__9187\,
            I => \N__9097\
        );

    \I__2144\ : ClkMux
    port map (
            O => \N__9186\,
            I => \N__9097\
        );

    \I__2143\ : ClkMux
    port map (
            O => \N__9185\,
            I => \N__9097\
        );

    \I__2142\ : ClkMux
    port map (
            O => \N__9184\,
            I => \N__9097\
        );

    \I__2141\ : ClkMux
    port map (
            O => \N__9183\,
            I => \N__9097\
        );

    \I__2140\ : ClkMux
    port map (
            O => \N__9182\,
            I => \N__9097\
        );

    \I__2139\ : GlobalMux
    port map (
            O => \N__9097\,
            I => \CLK80_OUT\
        );

    \I__2138\ : CascadeMux
    port map (
            O => \N__9094\,
            I => \N__9086\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9078\
        );

    \I__2136\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9075\
        );

    \I__2135\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9072\
        );

    \I__2134\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9063\
        );

    \I__2133\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9063\
        );

    \I__2132\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9063\
        );

    \I__2131\ : InMux
    port map (
            O => \N__9085\,
            I => \N__9063\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9058\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9083\,
            I => \N__9058\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9082\,
            I => \N__9055\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9081\,
            I => \N__9052\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__9078\,
            I => \N__9039\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__9075\,
            I => \N__9027\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9072\,
            I => \N__9024\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__9063\,
            I => \N__9017\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9058\,
            I => \N__9012\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__9055\,
            I => \N__9007\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9052\,
            I => \N__8999\
        );

    \I__2119\ : SRMux
    port map (
            O => \N__9051\,
            I => \N__8911\
        );

    \I__2118\ : SRMux
    port map (
            O => \N__9050\,
            I => \N__8911\
        );

    \I__2117\ : SRMux
    port map (
            O => \N__9049\,
            I => \N__8911\
        );

    \I__2116\ : SRMux
    port map (
            O => \N__9048\,
            I => \N__8911\
        );

    \I__2115\ : SRMux
    port map (
            O => \N__9047\,
            I => \N__8911\
        );

    \I__2114\ : SRMux
    port map (
            O => \N__9046\,
            I => \N__8911\
        );

    \I__2113\ : SRMux
    port map (
            O => \N__9045\,
            I => \N__8911\
        );

    \I__2112\ : SRMux
    port map (
            O => \N__9044\,
            I => \N__8911\
        );

    \I__2111\ : SRMux
    port map (
            O => \N__9043\,
            I => \N__8911\
        );

    \I__2110\ : SRMux
    port map (
            O => \N__9042\,
            I => \N__8911\
        );

    \I__2109\ : Glb2LocalMux
    port map (
            O => \N__9039\,
            I => \N__8911\
        );

    \I__2108\ : SRMux
    port map (
            O => \N__9038\,
            I => \N__8911\
        );

    \I__2107\ : SRMux
    port map (
            O => \N__9037\,
            I => \N__8911\
        );

    \I__2106\ : SRMux
    port map (
            O => \N__9036\,
            I => \N__8911\
        );

    \I__2105\ : SRMux
    port map (
            O => \N__9035\,
            I => \N__8911\
        );

    \I__2104\ : SRMux
    port map (
            O => \N__9034\,
            I => \N__8911\
        );

    \I__2103\ : SRMux
    port map (
            O => \N__9033\,
            I => \N__8911\
        );

    \I__2102\ : SRMux
    port map (
            O => \N__9032\,
            I => \N__8911\
        );

    \I__2101\ : SRMux
    port map (
            O => \N__9031\,
            I => \N__8911\
        );

    \I__2100\ : SRMux
    port map (
            O => \N__9030\,
            I => \N__8911\
        );

    \I__2099\ : Glb2LocalMux
    port map (
            O => \N__9027\,
            I => \N__8911\
        );

    \I__2098\ : Glb2LocalMux
    port map (
            O => \N__9024\,
            I => \N__8911\
        );

    \I__2097\ : SRMux
    port map (
            O => \N__9023\,
            I => \N__8911\
        );

    \I__2096\ : SRMux
    port map (
            O => \N__9022\,
            I => \N__8911\
        );

    \I__2095\ : SRMux
    port map (
            O => \N__9021\,
            I => \N__8911\
        );

    \I__2094\ : SRMux
    port map (
            O => \N__9020\,
            I => \N__8911\
        );

    \I__2093\ : Glb2LocalMux
    port map (
            O => \N__9017\,
            I => \N__8911\
        );

    \I__2092\ : SRMux
    port map (
            O => \N__9016\,
            I => \N__8911\
        );

    \I__2091\ : SRMux
    port map (
            O => \N__9015\,
            I => \N__8911\
        );

    \I__2090\ : Glb2LocalMux
    port map (
            O => \N__9012\,
            I => \N__8911\
        );

    \I__2089\ : SRMux
    port map (
            O => \N__9011\,
            I => \N__8911\
        );

    \I__2088\ : SRMux
    port map (
            O => \N__9010\,
            I => \N__8911\
        );

    \I__2087\ : Glb2LocalMux
    port map (
            O => \N__9007\,
            I => \N__8911\
        );

    \I__2086\ : SRMux
    port map (
            O => \N__9006\,
            I => \N__8911\
        );

    \I__2085\ : SRMux
    port map (
            O => \N__9005\,
            I => \N__8911\
        );

    \I__2084\ : SRMux
    port map (
            O => \N__9004\,
            I => \N__8911\
        );

    \I__2083\ : SRMux
    port map (
            O => \N__9003\,
            I => \N__8911\
        );

    \I__2082\ : SRMux
    port map (
            O => \N__9002\,
            I => \N__8911\
        );

    \I__2081\ : Glb2LocalMux
    port map (
            O => \N__8999\,
            I => \N__8911\
        );

    \I__2080\ : SRMux
    port map (
            O => \N__8998\,
            I => \N__8911\
        );

    \I__2079\ : SRMux
    port map (
            O => \N__8997\,
            I => \N__8911\
        );

    \I__2078\ : SRMux
    port map (
            O => \N__8996\,
            I => \N__8911\
        );

    \I__2077\ : GlobalMux
    port map (
            O => \N__8911\,
            I => \N__8908\
        );

    \I__2076\ : gio2CtrlBuf
    port map (
            O => \N__8908\,
            I => \RESETn_c_i_g\
        );

    \I__2075\ : CascadeMux
    port map (
            O => \N__8905\,
            I => \N__8898\
        );

    \I__2074\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8893\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__8903\,
            I => \N__8890\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__8902\,
            I => \N__8887\
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__8901\,
            I => \N__8884\
        );

    \I__2070\ : InMux
    port map (
            O => \N__8898\,
            I => \N__8881\
        );

    \I__2069\ : InMux
    port map (
            O => \N__8897\,
            I => \N__8876\
        );

    \I__2068\ : InMux
    port map (
            O => \N__8896\,
            I => \N__8876\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__8893\,
            I => \N__8873\
        );

    \I__2066\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8870\
        );

    \I__2065\ : InMux
    port map (
            O => \N__8887\,
            I => \N__8863\
        );

    \I__2064\ : InMux
    port map (
            O => \N__8884\,
            I => \N__8863\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__8881\,
            I => \N__8853\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__8876\,
            I => \N__8853\
        );

    \I__2061\ : Span4Mux_v
    port map (
            O => \N__8873\,
            I => \N__8853\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__8870\,
            I => \N__8853\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__8869\,
            I => \N__8849\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__8868\,
            I => \N__8845\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__8863\,
            I => \N__8842\
        );

    \I__2056\ : CascadeMux
    port map (
            O => \N__8862\,
            I => \N__8838\
        );

    \I__2055\ : Span4Mux_h
    port map (
            O => \N__8853\,
            I => \N__8832\
        );

    \I__2054\ : InMux
    port map (
            O => \N__8852\,
            I => \N__8829\
        );

    \I__2053\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8826\
        );

    \I__2052\ : InMux
    port map (
            O => \N__8848\,
            I => \N__8821\
        );

    \I__2051\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8821\
        );

    \I__2050\ : Span4Mux_h
    port map (
            O => \N__8842\,
            I => \N__8818\
        );

    \I__2049\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8807\
        );

    \I__2048\ : InMux
    port map (
            O => \N__8838\,
            I => \N__8807\
        );

    \I__2047\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8807\
        );

    \I__2046\ : InMux
    port map (
            O => \N__8836\,
            I => \N__8807\
        );

    \I__2045\ : InMux
    port map (
            O => \N__8835\,
            I => \N__8807\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__8832\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__8829\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__8826\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__8821\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__8818\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__8807\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2038\ : IoInMux
    port map (
            O => \N__8794\,
            I => \N__8791\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__8791\,
            I => \N__8788\
        );

    \I__2036\ : IoSpan4Mux
    port map (
            O => \N__8788\,
            I => \N__8785\
        );

    \I__2035\ : Span4Mux_s0_v
    port map (
            O => \N__8785\,
            I => \N__8782\
        );

    \I__2034\ : Sp12to4
    port map (
            O => \N__8782\,
            I => \N__8779\
        );

    \I__2033\ : Span12Mux_h
    port map (
            O => \N__8779\,
            I => \N__8776\
        );

    \I__2032\ : Odrv12
    port map (
            O => \N__8776\,
            I => \CASn_c\
        );

    \I__2031\ : InMux
    port map (
            O => \N__8773\,
            I => \N__8769\
        );

    \I__2030\ : InMux
    port map (
            O => \N__8772\,
            I => \N__8766\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__8769\,
            I => \N__8763\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__8766\,
            I => \N__8760\
        );

    \I__2027\ : Span4Mux_h
    port map (
            O => \N__8763\,
            I => \N__8755\
        );

    \I__2026\ : Span4Mux_h
    port map (
            O => \N__8760\,
            I => \N__8752\
        );

    \I__2025\ : InMux
    port map (
            O => \N__8759\,
            I => \N__8747\
        );

    \I__2024\ : InMux
    port map (
            O => \N__8758\,
            I => \N__8747\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__8755\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2022\ : Odrv4
    port map (
            O => \N__8752\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__8747\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2020\ : IoInMux
    port map (
            O => \N__8740\,
            I => \N__8737\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__8737\,
            I => \N__8734\
        );

    \I__2018\ : Span4Mux_s2_v
    port map (
            O => \N__8734\,
            I => \N__8731\
        );

    \I__2017\ : Sp12to4
    port map (
            O => \N__8731\,
            I => \N__8728\
        );

    \I__2016\ : Span12Mux_h
    port map (
            O => \N__8728\,
            I => \N__8725\
        );

    \I__2015\ : Odrv12
    port map (
            O => \N__8725\,
            I => \CRCSn_c\
        );

    \I__2014\ : InMux
    port map (
            O => \N__8722\,
            I => \N__8719\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__8719\,
            I => \N__8715\
        );

    \I__2012\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8712\
        );

    \I__2011\ : Span4Mux_v
    port map (
            O => \N__8715\,
            I => \N__8709\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__8712\,
            I => \N__8706\
        );

    \I__2009\ : Sp12to4
    port map (
            O => \N__8709\,
            I => \N__8701\
        );

    \I__2008\ : Span12Mux_v
    port map (
            O => \N__8706\,
            I => \N__8701\
        );

    \I__2007\ : Span12Mux_h
    port map (
            O => \N__8701\,
            I => \N__8698\
        );

    \I__2006\ : Span12Mux_v
    port map (
            O => \N__8698\,
            I => \N__8695\
        );

    \I__2005\ : Odrv12
    port map (
            O => \N__8695\,
            I => \DRA_c_1\
        );

    \I__2004\ : InMux
    port map (
            O => \N__8692\,
            I => \N__8689\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__8689\,
            I => \N__8686\
        );

    \I__2002\ : Span4Mux_v
    port map (
            O => \N__8686\,
            I => \N__8683\
        );

    \I__2001\ : Odrv4
    port map (
            O => \N__8683\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2000\ : InMux
    port map (
            O => \N__8680\,
            I => \N__8676\
        );

    \I__1999\ : InMux
    port map (
            O => \N__8679\,
            I => \N__8673\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__8676\,
            I => \N__8670\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__8673\,
            I => \N__8667\
        );

    \I__1996\ : Span4Mux_h
    port map (
            O => \N__8670\,
            I => \N__8664\
        );

    \I__1995\ : Span4Mux_v
    port map (
            O => \N__8667\,
            I => \N__8661\
        );

    \I__1994\ : Span4Mux_v
    port map (
            O => \N__8664\,
            I => \N__8658\
        );

    \I__1993\ : Sp12to4
    port map (
            O => \N__8661\,
            I => \N__8655\
        );

    \I__1992\ : Span4Mux_h
    port map (
            O => \N__8658\,
            I => \N__8652\
        );

    \I__1991\ : Span12Mux_h
    port map (
            O => \N__8655\,
            I => \N__8649\
        );

    \I__1990\ : Span4Mux_h
    port map (
            O => \N__8652\,
            I => \N__8646\
        );

    \I__1989\ : Odrv12
    port map (
            O => \N__8649\,
            I => \DRA_c_7\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__8646\,
            I => \DRA_c_7\
        );

    \I__1987\ : InMux
    port map (
            O => \N__8641\,
            I => \N__8638\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__8638\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__8635\,
            I => \N__8632\
        );

    \I__1984\ : InMux
    port map (
            O => \N__8632\,
            I => \N__8629\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__8629\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8626\,
            I => \N__8622\
        );

    \I__1981\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8619\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__8622\,
            I => \N__8614\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__8619\,
            I => \N__8614\
        );

    \I__1978\ : Span4Mux_v
    port map (
            O => \N__8614\,
            I => \N__8611\
        );

    \I__1977\ : Sp12to4
    port map (
            O => \N__8611\,
            I => \N__8608\
        );

    \I__1976\ : Span12Mux_h
    port map (
            O => \N__8608\,
            I => \N__8605\
        );

    \I__1975\ : Odrv12
    port map (
            O => \N__8605\,
            I => \DRA_c_8\
        );

    \I__1974\ : InMux
    port map (
            O => \N__8602\,
            I => \N__8599\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__8599\,
            I => \N__8596\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__8596\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1971\ : CEMux
    port map (
            O => \N__8593\,
            I => \N__8589\
        );

    \I__1970\ : CEMux
    port map (
            O => \N__8592\,
            I => \N__8586\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__8589\,
            I => \N__8582\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__8586\,
            I => \N__8578\
        );

    \I__1967\ : CEMux
    port map (
            O => \N__8585\,
            I => \N__8575\
        );

    \I__1966\ : Span4Mux_h
    port map (
            O => \N__8582\,
            I => \N__8572\
        );

    \I__1965\ : CEMux
    port map (
            O => \N__8581\,
            I => \N__8569\
        );

    \I__1964\ : Span4Mux_h
    port map (
            O => \N__8578\,
            I => \N__8566\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__8575\,
            I => \N__8563\
        );

    \I__1962\ : Span4Mux_h
    port map (
            O => \N__8572\,
            I => \N__8558\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__8569\,
            I => \N__8558\
        );

    \I__1960\ : Odrv4
    port map (
            O => \N__8566\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__8563\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__8558\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1957\ : CEMux
    port map (
            O => \N__8551\,
            I => \N__8548\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__8548\,
            I => \N__8544\
        );

    \I__1955\ : CEMux
    port map (
            O => \N__8547\,
            I => \N__8541\
        );

    \I__1954\ : Span4Mux_v
    port map (
            O => \N__8544\,
            I => \N__8536\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__8541\,
            I => \N__8536\
        );

    \I__1952\ : Span4Mux_h
    port map (
            O => \N__8536\,
            I => \N__8533\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__8533\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8530\,
            I => \N__8524\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__8529\,
            I => \N__8518\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__8528\,
            I => \N__8515\
        );

    \I__1947\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8507\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__8524\,
            I => \N__8504\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8523\,
            I => \N__8501\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8490\
        );

    \I__1943\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8490\
        );

    \I__1942\ : InMux
    port map (
            O => \N__8518\,
            I => \N__8490\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8515\,
            I => \N__8490\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8514\,
            I => \N__8490\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8487\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__8512\,
            I => \N__8483\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8511\,
            I => \N__8478\
        );

    \I__1936\ : InMux
    port map (
            O => \N__8510\,
            I => \N__8478\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__8507\,
            I => \N__8475\
        );

    \I__1934\ : Span4Mux_v
    port map (
            O => \N__8504\,
            I => \N__8472\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__8501\,
            I => \N__8465\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__8490\,
            I => \N__8465\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__8487\,
            I => \N__8465\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__8486\,
            I => \N__8462\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8459\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__8478\,
            I => \N__8456\
        );

    \I__1927\ : Span4Mux_v
    port map (
            O => \N__8475\,
            I => \N__8449\
        );

    \I__1926\ : Span4Mux_h
    port map (
            O => \N__8472\,
            I => \N__8449\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__8465\,
            I => \N__8449\
        );

    \I__1924\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8446\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__8459\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__8456\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__8449\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__8446\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1919\ : IoInMux
    port map (
            O => \N__8437\,
            I => \N__8434\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__8434\,
            I => \N__8431\
        );

    \I__1917\ : Span4Mux_s0_h
    port map (
            O => \N__8431\,
            I => \N__8428\
        );

    \I__1916\ : Sp12to4
    port map (
            O => \N__8428\,
            I => \N__8425\
        );

    \I__1915\ : Span12Mux_s7_v
    port map (
            O => \N__8425\,
            I => \N__8422\
        );

    \I__1914\ : Span12Mux_h
    port map (
            O => \N__8422\,
            I => \N__8419\
        );

    \I__1913\ : Odrv12
    port map (
            O => \N__8419\,
            I => \WEn_c\
        );

    \I__1912\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8413\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__8413\,
            I => \N__8410\
        );

    \I__1910\ : Span12Mux_h
    port map (
            O => \N__8410\,
            I => \N__8407\
        );

    \I__1909\ : Odrv12
    port map (
            O => \N__8407\,
            I => \RAS1n_c\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__8404\,
            I => \N__8392\
        );

    \I__1907\ : InMux
    port map (
            O => \N__8403\,
            I => \N__8377\
        );

    \I__1906\ : InMux
    port map (
            O => \N__8402\,
            I => \N__8374\
        );

    \I__1905\ : InMux
    port map (
            O => \N__8401\,
            I => \N__8368\
        );

    \I__1904\ : InMux
    port map (
            O => \N__8400\,
            I => \N__8365\
        );

    \I__1903\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8362\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8398\,
            I => \N__8357\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8397\,
            I => \N__8357\
        );

    \I__1900\ : InMux
    port map (
            O => \N__8396\,
            I => \N__8354\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__8395\,
            I => \N__8350\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8392\,
            I => \N__8347\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8391\,
            I => \N__8342\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8342\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8337\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8388\,
            I => \N__8337\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8334\
        );

    \I__1892\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8331\
        );

    \I__1891\ : InMux
    port map (
            O => \N__8385\,
            I => \N__8326\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8384\,
            I => \N__8326\
        );

    \I__1889\ : InMux
    port map (
            O => \N__8383\,
            I => \N__8317\
        );

    \I__1888\ : InMux
    port map (
            O => \N__8382\,
            I => \N__8317\
        );

    \I__1887\ : InMux
    port map (
            O => \N__8381\,
            I => \N__8317\
        );

    \I__1886\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8317\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8377\,
            I => \N__8314\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__8374\,
            I => \N__8311\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8373\,
            I => \N__8304\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8372\,
            I => \N__8304\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8371\,
            I => \N__8304\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__8368\,
            I => \N__8299\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__8365\,
            I => \N__8299\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8362\,
            I => \N__8294\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8357\,
            I => \N__8294\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8354\,
            I => \N__8291\
        );

    \I__1875\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8288\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8285\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__8347\,
            I => \N__8278\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8342\,
            I => \N__8278\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8337\,
            I => \N__8267\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8334\,
            I => \N__8267\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__8331\,
            I => \N__8267\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8326\,
            I => \N__8267\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8317\,
            I => \N__8267\
        );

    \I__1866\ : Span4Mux_v
    port map (
            O => \N__8314\,
            I => \N__8260\
        );

    \I__1865\ : Span4Mux_v
    port map (
            O => \N__8311\,
            I => \N__8260\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8304\,
            I => \N__8260\
        );

    \I__1863\ : Span4Mux_v
    port map (
            O => \N__8299\,
            I => \N__8255\
        );

    \I__1862\ : Span4Mux_v
    port map (
            O => \N__8294\,
            I => \N__8255\
        );

    \I__1861\ : Span4Mux_h
    port map (
            O => \N__8291\,
            I => \N__8248\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8288\,
            I => \N__8248\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__8285\,
            I => \N__8248\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8284\,
            I => \N__8245\
        );

    \I__1857\ : InMux
    port map (
            O => \N__8283\,
            I => \N__8242\
        );

    \I__1856\ : Span4Mux_v
    port map (
            O => \N__8278\,
            I => \N__8239\
        );

    \I__1855\ : Span4Mux_v
    port map (
            O => \N__8267\,
            I => \N__8234\
        );

    \I__1854\ : Span4Mux_h
    port map (
            O => \N__8260\,
            I => \N__8234\
        );

    \I__1853\ : Span4Mux_h
    port map (
            O => \N__8255\,
            I => \N__8229\
        );

    \I__1852\ : Span4Mux_v
    port map (
            O => \N__8248\,
            I => \N__8229\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__8245\,
            I => \CPU_CYCLEm\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8242\,
            I => \CPU_CYCLEm\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__8239\,
            I => \CPU_CYCLEm\
        );

    \I__1848\ : Odrv4
    port map (
            O => \N__8234\,
            I => \CPU_CYCLEm\
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__8229\,
            I => \CPU_CYCLEm\
        );

    \I__1846\ : InMux
    port map (
            O => \N__8218\,
            I => \N__8215\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8215\,
            I => \N__8212\
        );

    \I__1844\ : Sp12to4
    port map (
            O => \N__8212\,
            I => \N__8209\
        );

    \I__1843\ : Span12Mux_v
    port map (
            O => \N__8209\,
            I => \N__8206\
        );

    \I__1842\ : Span12Mux_h
    port map (
            O => \N__8206\,
            I => \N__8203\
        );

    \I__1841\ : Odrv12
    port map (
            O => \N__8203\,
            I => \A_c_20\
        );

    \I__1840\ : IoInMux
    port map (
            O => \N__8200\,
            I => \N__8197\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8197\,
            I => \N__8194\
        );

    \I__1838\ : Span12Mux_s6_v
    port map (
            O => \N__8194\,
            I => \N__8190\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8193\,
            I => \N__8187\
        );

    \I__1836\ : Odrv12
    port map (
            O => \N__8190\,
            I => \BANK0_c\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8187\,
            I => \BANK0_c\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8182\,
            I => \N__8175\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8181\,
            I => \N__8175\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__8180\,
            I => \N__8167\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__8175\,
            I => \N__8164\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__8174\,
            I => \N__8161\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8173\,
            I => \N__8153\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8172\,
            I => \N__8153\
        );

    \I__1827\ : InMux
    port map (
            O => \N__8171\,
            I => \N__8153\
        );

    \I__1826\ : InMux
    port map (
            O => \N__8170\,
            I => \N__8150\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8147\
        );

    \I__1824\ : Span4Mux_h
    port map (
            O => \N__8164\,
            I => \N__8144\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8161\,
            I => \N__8139\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8160\,
            I => \N__8139\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8153\,
            I => \N__8136\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8150\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8147\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__8144\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__8139\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1816\ : Odrv12
    port map (
            O => \N__8136\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8122\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8122\,
            I => \N__8119\
        );

    \I__1813\ : Span4Mux_h
    port map (
            O => \N__8119\,
            I => \N__8116\
        );

    \I__1812\ : Odrv4
    port map (
            O => \N__8116\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__8113\,
            I => \U712_CHIP_RAM.DMA_CYCLE_7_cascade_\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8110\,
            I => \N__8101\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8101\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8101\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8101\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0\
        );

    \I__1806\ : IoInMux
    port map (
            O => \N__8098\,
            I => \N__8095\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__8095\,
            I => \N__8092\
        );

    \I__1804\ : Span4Mux_s2_v
    port map (
            O => \N__8092\,
            I => \N__8088\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8085\
        );

    \I__1802\ : Sp12to4
    port map (
            O => \N__8088\,
            I => \N__8081\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8085\,
            I => \N__8078\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8084\,
            I => \N__8075\
        );

    \I__1799\ : Span12Mux_h
    port map (
            O => \N__8081\,
            I => \N__8072\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__8078\,
            I => \N__8069\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8075\,
            I => \N__8066\
        );

    \I__1796\ : Span12Mux_v
    port map (
            O => \N__8072\,
            I => \N__8062\
        );

    \I__1795\ : Span4Mux_h
    port map (
            O => \N__8069\,
            I => \N__8057\
        );

    \I__1794\ : Span4Mux_h
    port map (
            O => \N__8066\,
            I => \N__8057\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8054\
        );

    \I__1792\ : Odrv12
    port map (
            O => \N__8062\,
            I => \DBENn_c\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__8057\,
            I => \DBENn_c\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8054\,
            I => \DBENn_c\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8047\,
            I => \N__8044\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8044\,
            I => \N__8040\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8043\,
            I => \N__8037\
        );

    \I__1786\ : Span4Mux_h
    port map (
            O => \N__8040\,
            I => \N__8032\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__8037\,
            I => \N__8032\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__8032\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1783\ : InMux
    port map (
            O => \N__8029\,
            I => \N__8024\
        );

    \I__1782\ : InMux
    port map (
            O => \N__8028\,
            I => \N__8020\
        );

    \I__1781\ : CascadeMux
    port map (
            O => \N__8027\,
            I => \N__8017\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8024\,
            I => \N__8014\
        );

    \I__1779\ : InMux
    port map (
            O => \N__8023\,
            I => \N__8010\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__8020\,
            I => \N__8007\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8017\,
            I => \N__8004\
        );

    \I__1776\ : Span4Mux_h
    port map (
            O => \N__8014\,
            I => \N__8001\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8013\,
            I => \N__7998\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__8010\,
            I => \N__7993\
        );

    \I__1773\ : Span4Mux_v
    port map (
            O => \N__8007\,
            I => \N__7993\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8004\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__8001\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__7998\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__7993\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1768\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7981\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__7981\,
            I => \U712_CHIP_RAM.N_148\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__7978\,
            I => \N__7972\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__7977\,
            I => \N__7969\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__7976\,
            I => \N__7960\
        );

    \I__1763\ : CascadeMux
    port map (
            O => \N__7975\,
            I => \N__7957\
        );

    \I__1762\ : InMux
    port map (
            O => \N__7972\,
            I => \N__7953\
        );

    \I__1761\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7950\
        );

    \I__1760\ : InMux
    port map (
            O => \N__7968\,
            I => \N__7946\
        );

    \I__1759\ : InMux
    port map (
            O => \N__7967\,
            I => \N__7942\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__7966\,
            I => \N__7937\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__7965\,
            I => \N__7934\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__7964\,
            I => \N__7931\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__7963\,
            I => \N__7928\
        );

    \I__1754\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7921\
        );

    \I__1753\ : InMux
    port map (
            O => \N__7957\,
            I => \N__7921\
        );

    \I__1752\ : InMux
    port map (
            O => \N__7956\,
            I => \N__7921\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__7953\,
            I => \N__7918\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__7950\,
            I => \N__7915\
        );

    \I__1749\ : InMux
    port map (
            O => \N__7949\,
            I => \N__7912\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__7946\,
            I => \N__7909\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__7945\,
            I => \N__7900\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__7942\,
            I => \N__7895\
        );

    \I__1745\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7892\
        );

    \I__1744\ : InMux
    port map (
            O => \N__7940\,
            I => \N__7885\
        );

    \I__1743\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7885\
        );

    \I__1742\ : InMux
    port map (
            O => \N__7934\,
            I => \N__7885\
        );

    \I__1741\ : InMux
    port map (
            O => \N__7931\,
            I => \N__7882\
        );

    \I__1740\ : InMux
    port map (
            O => \N__7928\,
            I => \N__7879\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__7921\,
            I => \N__7868\
        );

    \I__1738\ : Span4Mux_v
    port map (
            O => \N__7918\,
            I => \N__7868\
        );

    \I__1737\ : Span4Mux_v
    port map (
            O => \N__7915\,
            I => \N__7868\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__7912\,
            I => \N__7868\
        );

    \I__1735\ : Span4Mux_h
    port map (
            O => \N__7909\,
            I => \N__7868\
        );

    \I__1734\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7865\
        );

    \I__1733\ : InMux
    port map (
            O => \N__7907\,
            I => \N__7860\
        );

    \I__1732\ : InMux
    port map (
            O => \N__7906\,
            I => \N__7860\
        );

    \I__1731\ : InMux
    port map (
            O => \N__7905\,
            I => \N__7853\
        );

    \I__1730\ : InMux
    port map (
            O => \N__7904\,
            I => \N__7853\
        );

    \I__1729\ : InMux
    port map (
            O => \N__7903\,
            I => \N__7853\
        );

    \I__1728\ : InMux
    port map (
            O => \N__7900\,
            I => \N__7846\
        );

    \I__1727\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7846\
        );

    \I__1726\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7846\
        );

    \I__1725\ : Odrv4
    port map (
            O => \N__7895\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__7892\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__7885\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__7882\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__7879\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1720\ : Odrv4
    port map (
            O => \N__7868\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__7865\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__7860\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__7853\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__7846\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1715\ : IoInMux
    port map (
            O => \N__7825\,
            I => \N__7822\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__7822\,
            I => \N__7819\
        );

    \I__1713\ : Span4Mux_s3_h
    port map (
            O => \N__7819\,
            I => \N__7816\
        );

    \I__1712\ : Sp12to4
    port map (
            O => \N__7816\,
            I => \N__7813\
        );

    \I__1711\ : Span12Mux_v
    port map (
            O => \N__7813\,
            I => \N__7809\
        );

    \I__1710\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7806\
        );

    \I__1709\ : Odrv12
    port map (
            O => \N__7809\,
            I => \CLK_EN_c\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__7806\,
            I => \CLK_EN_c\
        );

    \I__1707\ : InMux
    port map (
            O => \N__7801\,
            I => \N__7794\
        );

    \I__1706\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7794\
        );

    \I__1705\ : InMux
    port map (
            O => \N__7799\,
            I => \N__7791\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__7794\,
            I => \N__7788\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__7791\,
            I => \N__7785\
        );

    \I__1702\ : Span12Mux_h
    port map (
            O => \N__7788\,
            I => \N__7782\
        );

    \I__1701\ : Span12Mux_h
    port map (
            O => \N__7785\,
            I => \N__7779\
        );

    \I__1700\ : Span12Mux_v
    port map (
            O => \N__7782\,
            I => \N__7776\
        );

    \I__1699\ : Span12Mux_v
    port map (
            O => \N__7779\,
            I => \N__7773\
        );

    \I__1698\ : Odrv12
    port map (
            O => \N__7776\,
            I => \CASLn_c\
        );

    \I__1697\ : Odrv12
    port map (
            O => \N__7773\,
            I => \CASLn_c\
        );

    \I__1696\ : InMux
    port map (
            O => \N__7768\,
            I => \N__7763\
        );

    \I__1695\ : InMux
    port map (
            O => \N__7767\,
            I => \N__7758\
        );

    \I__1694\ : InMux
    port map (
            O => \N__7766\,
            I => \N__7758\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__7763\,
            I => \N__7755\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__7758\,
            I => \N__7752\
        );

    \I__1691\ : Span4Mux_v
    port map (
            O => \N__7755\,
            I => \N__7749\
        );

    \I__1690\ : Sp12to4
    port map (
            O => \N__7752\,
            I => \N__7746\
        );

    \I__1689\ : Sp12to4
    port map (
            O => \N__7749\,
            I => \N__7743\
        );

    \I__1688\ : Span12Mux_v
    port map (
            O => \N__7746\,
            I => \N__7740\
        );

    \I__1687\ : Span12Mux_h
    port map (
            O => \N__7743\,
            I => \N__7737\
        );

    \I__1686\ : Span12Mux_h
    port map (
            O => \N__7740\,
            I => \N__7734\
        );

    \I__1685\ : Span12Mux_v
    port map (
            O => \N__7737\,
            I => \N__7731\
        );

    \I__1684\ : Odrv12
    port map (
            O => \N__7734\,
            I => \CASUn_c\
        );

    \I__1683\ : Odrv12
    port map (
            O => \N__7731\,
            I => \CASUn_c\
        );

    \I__1682\ : InMux
    port map (
            O => \N__7726\,
            I => \N__7722\
        );

    \I__1681\ : InMux
    port map (
            O => \N__7725\,
            I => \N__7718\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__7722\,
            I => \N__7715\
        );

    \I__1679\ : InMux
    port map (
            O => \N__7721\,
            I => \N__7712\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__7718\,
            I => \N__7709\
        );

    \I__1677\ : Odrv4
    port map (
            O => \N__7715\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__7712\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1675\ : Odrv4
    port map (
            O => \N__7709\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1674\ : InMux
    port map (
            O => \N__7702\,
            I => \N__7699\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__7699\,
            I => \N__7693\
        );

    \I__1672\ : InMux
    port map (
            O => \N__7698\,
            I => \N__7690\
        );

    \I__1671\ : InMux
    port map (
            O => \N__7697\,
            I => \N__7687\
        );

    \I__1670\ : InMux
    port map (
            O => \N__7696\,
            I => \N__7684\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__7693\,
            I => \N__7679\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__7690\,
            I => \N__7676\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__7687\,
            I => \N__7673\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__7684\,
            I => \N__7670\
        );

    \I__1665\ : InMux
    port map (
            O => \N__7683\,
            I => \N__7667\
        );

    \I__1664\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7664\
        );

    \I__1663\ : Odrv4
    port map (
            O => \N__7679\,
            I => \DMA_CYCLEm\
        );

    \I__1662\ : Odrv12
    port map (
            O => \N__7676\,
            I => \DMA_CYCLEm\
        );

    \I__1661\ : Odrv4
    port map (
            O => \N__7673\,
            I => \DMA_CYCLEm\
        );

    \I__1660\ : Odrv4
    port map (
            O => \N__7670\,
            I => \DMA_CYCLEm\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__7667\,
            I => \DMA_CYCLEm\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__7664\,
            I => \DMA_CYCLEm\
        );

    \I__1657\ : InMux
    port map (
            O => \N__7651\,
            I => \N__7647\
        );

    \I__1656\ : InMux
    port map (
            O => \N__7650\,
            I => \N__7644\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__7647\,
            I => \N__7639\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__7644\,
            I => \N__7636\
        );

    \I__1653\ : InMux
    port map (
            O => \N__7643\,
            I => \N__7633\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__7642\,
            I => \N__7630\
        );

    \I__1651\ : Sp12to4
    port map (
            O => \N__7639\,
            I => \N__7627\
        );

    \I__1650\ : Span4Mux_h
    port map (
            O => \N__7636\,
            I => \N__7622\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__7633\,
            I => \N__7622\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7630\,
            I => \N__7619\
        );

    \I__1647\ : Odrv12
    port map (
            O => \N__7627\,
            I => \REG_CYCLEm\
        );

    \I__1646\ : Odrv4
    port map (
            O => \N__7622\,
            I => \REG_CYCLEm\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__7619\,
            I => \REG_CYCLEm\
        );

    \I__1644\ : IoInMux
    port map (
            O => \N__7612\,
            I => \N__7609\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7609\,
            I => \N__7606\
        );

    \I__1642\ : Span4Mux_s2_v
    port map (
            O => \N__7606\,
            I => \N__7603\
        );

    \I__1641\ : Span4Mux_v
    port map (
            O => \N__7603\,
            I => \N__7600\
        );

    \I__1640\ : Sp12to4
    port map (
            O => \N__7600\,
            I => \N__7597\
        );

    \I__1639\ : Span12Mux_h
    port map (
            O => \N__7597\,
            I => \N__7594\
        );

    \I__1638\ : Odrv12
    port map (
            O => \N__7594\,
            I => \DRDENn_c\
        );

    \I__1637\ : InMux
    port map (
            O => \N__7591\,
            I => \N__7585\
        );

    \I__1636\ : InMux
    port map (
            O => \N__7590\,
            I => \N__7582\
        );

    \I__1635\ : InMux
    port map (
            O => \N__7589\,
            I => \N__7579\
        );

    \I__1634\ : InMux
    port map (
            O => \N__7588\,
            I => \N__7576\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7585\,
            I => \N__7570\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__7582\,
            I => \N__7570\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__7579\,
            I => \N__7566\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__7576\,
            I => \N__7563\
        );

    \I__1629\ : InMux
    port map (
            O => \N__7575\,
            I => \N__7560\
        );

    \I__1628\ : Span4Mux_v
    port map (
            O => \N__7570\,
            I => \N__7557\
        );

    \I__1627\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7554\
        );

    \I__1626\ : Span4Mux_h
    port map (
            O => \N__7566\,
            I => \N__7547\
        );

    \I__1625\ : Span4Mux_h
    port map (
            O => \N__7563\,
            I => \N__7547\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7560\,
            I => \N__7547\
        );

    \I__1623\ : Span4Mux_h
    port map (
            O => \N__7557\,
            I => \N__7544\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__7554\,
            I => \N__7539\
        );

    \I__1621\ : Sp12to4
    port map (
            O => \N__7547\,
            I => \N__7539\
        );

    \I__1620\ : Sp12to4
    port map (
            O => \N__7544\,
            I => \N__7534\
        );

    \I__1619\ : Span12Mux_v
    port map (
            O => \N__7539\,
            I => \N__7534\
        );

    \I__1618\ : Span12Mux_h
    port map (
            O => \N__7534\,
            I => \N__7531\
        );

    \I__1617\ : Odrv12
    port map (
            O => \N__7531\,
            I => \RESETn_c\
        );

    \I__1616\ : IoInMux
    port map (
            O => \N__7528\,
            I => \N__7525\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__7525\,
            I => \N__7522\
        );

    \I__1614\ : Span12Mux_s0_v
    port map (
            O => \N__7522\,
            I => \N__7519\
        );

    \I__1613\ : Odrv12
    port map (
            O => \N__7519\,
            I => \RESETn_c_i\
        );

    \I__1612\ : IoInMux
    port map (
            O => \N__7516\,
            I => \N__7513\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__7513\,
            I => \N__7510\
        );

    \I__1610\ : IoSpan4Mux
    port map (
            O => \N__7510\,
            I => \N__7507\
        );

    \I__1609\ : Sp12to4
    port map (
            O => \N__7507\,
            I => \N__7504\
        );

    \I__1608\ : Span12Mux_s9_v
    port map (
            O => \N__7504\,
            I => \N__7501\
        );

    \I__1607\ : Odrv12
    port map (
            O => \N__7501\,
            I => \RASn_c\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7498\,
            I => \N__7495\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__7495\,
            I => \N__7492\
        );

    \I__1604\ : Sp12to4
    port map (
            O => \N__7492\,
            I => \N__7489\
        );

    \I__1603\ : Span12Mux_v
    port map (
            O => \N__7489\,
            I => \N__7486\
        );

    \I__1602\ : Span12Mux_h
    port map (
            O => \N__7486\,
            I => \N__7483\
        );

    \I__1601\ : Odrv12
    port map (
            O => \N__7483\,
            I => \A_c_16\
        );

    \I__1600\ : CascadeMux
    port map (
            O => \N__7480\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7477\,
            I => \N__7474\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__7474\,
            I => \N__7471\
        );

    \I__1597\ : Sp12to4
    port map (
            O => \N__7471\,
            I => \N__7468\
        );

    \I__1596\ : Span12Mux_v
    port map (
            O => \N__7468\,
            I => \N__7465\
        );

    \I__1595\ : Span12Mux_h
    port map (
            O => \N__7465\,
            I => \N__7462\
        );

    \I__1594\ : Odrv12
    port map (
            O => \N__7462\,
            I => \A_c_18\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__7459\,
            I => \U712_CHIP_RAM.N_313_cascade_\
        );

    \I__1592\ : IoInMux
    port map (
            O => \N__7456\,
            I => \N__7453\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__7453\,
            I => \N__7450\
        );

    \I__1590\ : Span4Mux_s2_h
    port map (
            O => \N__7450\,
            I => \N__7447\
        );

    \I__1589\ : Span4Mux_v
    port map (
            O => \N__7447\,
            I => \N__7444\
        );

    \I__1588\ : Sp12to4
    port map (
            O => \N__7444\,
            I => \N__7441\
        );

    \I__1587\ : Span12Mux_h
    port map (
            O => \N__7441\,
            I => \N__7438\
        );

    \I__1586\ : Odrv12
    port map (
            O => \N__7438\,
            I => \CMA_c_7\
        );

    \I__1585\ : InMux
    port map (
            O => \N__7435\,
            I => \N__7432\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7432\,
            I => \N__7429\
        );

    \I__1583\ : Span4Mux_v
    port map (
            O => \N__7429\,
            I => \N__7426\
        );

    \I__1582\ : Span4Mux_v
    port map (
            O => \N__7426\,
            I => \N__7423\
        );

    \I__1581\ : Sp12to4
    port map (
            O => \N__7423\,
            I => \N__7420\
        );

    \I__1580\ : Span12Mux_h
    port map (
            O => \N__7420\,
            I => \N__7417\
        );

    \I__1579\ : Odrv12
    port map (
            O => \N__7417\,
            I => \A_c_17\
        );

    \I__1578\ : IoInMux
    port map (
            O => \N__7414\,
            I => \N__7411\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7411\,
            I => \N__7408\
        );

    \I__1576\ : IoSpan4Mux
    port map (
            O => \N__7408\,
            I => \N__7405\
        );

    \I__1575\ : IoSpan4Mux
    port map (
            O => \N__7405\,
            I => \N__7402\
        );

    \I__1574\ : Sp12to4
    port map (
            O => \N__7402\,
            I => \N__7399\
        );

    \I__1573\ : Span12Mux_s7_h
    port map (
            O => \N__7399\,
            I => \N__7396\
        );

    \I__1572\ : Odrv12
    port map (
            O => \N__7396\,
            I => \CMA_c_8\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7393\,
            I => \N__7387\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7392\,
            I => \N__7387\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7387\,
            I => \U712_CHIP_RAM.CMA_5_i_0_8\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__7384\,
            I => \N__7381\
        );

    \I__1567\ : InMux
    port map (
            O => \N__7381\,
            I => \N__7378\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7378\,
            I => \N__7375\
        );

    \I__1565\ : Span4Mux_v
    port map (
            O => \N__7375\,
            I => \N__7372\
        );

    \I__1564\ : Span4Mux_v
    port map (
            O => \N__7372\,
            I => \N__7369\
        );

    \I__1563\ : Sp12to4
    port map (
            O => \N__7369\,
            I => \N__7366\
        );

    \I__1562\ : Span12Mux_h
    port map (
            O => \N__7366\,
            I => \N__7363\
        );

    \I__1561\ : Odrv12
    port map (
            O => \N__7363\,
            I => \A_c_19\
        );

    \I__1560\ : IoInMux
    port map (
            O => \N__7360\,
            I => \N__7357\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7357\,
            I => \N__7354\
        );

    \I__1558\ : Span4Mux_s3_h
    port map (
            O => \N__7354\,
            I => \N__7351\
        );

    \I__1557\ : Sp12to4
    port map (
            O => \N__7351\,
            I => \N__7348\
        );

    \I__1556\ : Span12Mux_s11_v
    port map (
            O => \N__7348\,
            I => \N__7345\
        );

    \I__1555\ : Odrv12
    port map (
            O => \N__7345\,
            I => \CMA_c_9\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7342\,
            I => \N__7339\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__7339\,
            I => \N__7336\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__7336\,
            I => \U712_CHIP_RAM.N_309\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7322\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7315\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7331\,
            I => \N__7315\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7330\,
            I => \N__7312\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7329\,
            I => \N__7301\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7328\,
            I => \N__7301\
        );

    \I__1545\ : InMux
    port map (
            O => \N__7327\,
            I => \N__7301\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7326\,
            I => \N__7301\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7301\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__7322\,
            I => \N__7298\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7321\,
            I => \N__7295\
        );

    \I__1540\ : InMux
    port map (
            O => \N__7320\,
            I => \N__7291\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__7315\,
            I => \N__7284\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7312\,
            I => \N__7284\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__7301\,
            I => \N__7284\
        );

    \I__1536\ : Span4Mux_v
    port map (
            O => \N__7298\,
            I => \N__7279\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__7295\,
            I => \N__7279\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7274\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__7291\,
            I => \N__7271\
        );

    \I__1532\ : Span4Mux_h
    port map (
            O => \N__7284\,
            I => \N__7268\
        );

    \I__1531\ : Span4Mux_h
    port map (
            O => \N__7279\,
            I => \N__7265\
        );

    \I__1530\ : InMux
    port map (
            O => \N__7278\,
            I => \N__7262\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7277\,
            I => \N__7259\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7274\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1527\ : Odrv12
    port map (
            O => \N__7271\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__7268\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__7265\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7262\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7259\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1522\ : IoInMux
    port map (
            O => \N__7246\,
            I => \N__7243\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7243\,
            I => \N__7240\
        );

    \I__1520\ : Span4Mux_s3_h
    port map (
            O => \N__7240\,
            I => \N__7237\
        );

    \I__1519\ : Span4Mux_v
    port map (
            O => \N__7237\,
            I => \N__7234\
        );

    \I__1518\ : Sp12to4
    port map (
            O => \N__7234\,
            I => \N__7231\
        );

    \I__1517\ : Span12Mux_h
    port map (
            O => \N__7231\,
            I => \N__7228\
        );

    \I__1516\ : Odrv12
    port map (
            O => \N__7228\,
            I => \CMA_c_3\
        );

    \I__1515\ : CEMux
    port map (
            O => \N__7225\,
            I => \N__7222\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__7222\,
            I => \N__7219\
        );

    \I__1513\ : Span4Mux_v
    port map (
            O => \N__7219\,
            I => \N__7213\
        );

    \I__1512\ : CEMux
    port map (
            O => \N__7218\,
            I => \N__7210\
        );

    \I__1511\ : CEMux
    port map (
            O => \N__7217\,
            I => \N__7207\
        );

    \I__1510\ : CEMux
    port map (
            O => \N__7216\,
            I => \N__7204\
        );

    \I__1509\ : Span4Mux_h
    port map (
            O => \N__7213\,
            I => \N__7196\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7210\,
            I => \N__7196\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7207\,
            I => \N__7196\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7204\,
            I => \N__7193\
        );

    \I__1505\ : CEMux
    port map (
            O => \N__7203\,
            I => \N__7190\
        );

    \I__1504\ : Span4Mux_v
    port map (
            O => \N__7196\,
            I => \N__7187\
        );

    \I__1503\ : Span4Mux_v
    port map (
            O => \N__7193\,
            I => \N__7184\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7190\,
            I => \N__7179\
        );

    \I__1501\ : Span4Mux_v
    port map (
            O => \N__7187\,
            I => \N__7179\
        );

    \I__1500\ : Odrv4
    port map (
            O => \N__7184\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__7179\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1498\ : CascadeMux
    port map (
            O => \N__7174\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_cascade_\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7171\,
            I => \N__7166\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7170\,
            I => \N__7161\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7169\,
            I => \N__7161\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7166\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__7161\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7152\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7155\,
            I => \N__7148\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__7152\,
            I => \N__7141\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7151\,
            I => \N__7138\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7148\,
            I => \N__7134\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7147\,
            I => \N__7131\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7146\,
            I => \N__7122\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7122\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7144\,
            I => \N__7122\
        );

    \I__1483\ : Span4Mux_h
    port map (
            O => \N__7141\,
            I => \N__7119\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7138\,
            I => \N__7116\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7137\,
            I => \N__7113\
        );

    \I__1480\ : Span4Mux_h
    port map (
            O => \N__7134\,
            I => \N__7108\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7131\,
            I => \N__7108\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7103\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7129\,
            I => \N__7103\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__7122\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1475\ : Odrv4
    port map (
            O => \N__7119\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1474\ : Odrv12
    port map (
            O => \N__7116\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7113\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1472\ : Odrv4
    port map (
            O => \N__7108\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7103\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1470\ : CascadeMux
    port map (
            O => \N__7090\,
            I => \N__7086\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7089\,
            I => \N__7082\
        );

    \I__1468\ : InMux
    port map (
            O => \N__7086\,
            I => \N__7079\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7085\,
            I => \N__7076\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7082\,
            I => \N__7073\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7079\,
            I => \N__7067\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7076\,
            I => \N__7067\
        );

    \I__1463\ : Span4Mux_v
    port map (
            O => \N__7073\,
            I => \N__7064\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7072\,
            I => \N__7061\
        );

    \I__1461\ : Odrv4
    port map (
            O => \N__7067\,
            I => \U712_CHIP_RAM.N_428\
        );

    \I__1460\ : Odrv4
    port map (
            O => \N__7064\,
            I => \U712_CHIP_RAM.N_428\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7061\,
            I => \U712_CHIP_RAM.N_428\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7054\,
            I => \N__7051\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7051\,
            I => \N__7048\
        );

    \I__1456\ : Span4Mux_h
    port map (
            O => \N__7048\,
            I => \N__7045\
        );

    \I__1455\ : Odrv4
    port map (
            O => \N__7045\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7042\,
            I => \N__7038\
        );

    \I__1453\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7035\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__7038\,
            I => \N__7032\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7035\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__7032\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7027\,
            I => \N__7021\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7026\,
            I => \N__7015\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7025\,
            I => \N__7012\
        );

    \I__1446\ : InMux
    port map (
            O => \N__7024\,
            I => \N__7007\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7021\,
            I => \N__7004\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__7020\,
            I => \N__7001\
        );

    \I__1443\ : InMux
    port map (
            O => \N__7019\,
            I => \N__6995\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7018\,
            I => \N__6995\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7015\,
            I => \N__6990\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__7012\,
            I => \N__6990\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7011\,
            I => \N__6985\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7010\,
            I => \N__6985\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7007\,
            I => \N__6980\
        );

    \I__1436\ : Span4Mux_v
    port map (
            O => \N__7004\,
            I => \N__6980\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7001\,
            I => \N__6975\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6975\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__6995\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1432\ : Odrv4
    port map (
            O => \N__6990\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__6985\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1430\ : Odrv4
    port map (
            O => \N__6980\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__6975\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__6964\,
            I => \N__6958\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6963\,
            I => \N__6955\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6962\,
            I => \N__6949\
        );

    \I__1425\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6946\
        );

    \I__1424\ : InMux
    port map (
            O => \N__6958\,
            I => \N__6943\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__6955\,
            I => \N__6940\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__6954\,
            I => \N__6937\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__6953\,
            I => \N__6934\
        );

    \I__1420\ : InMux
    port map (
            O => \N__6952\,
            I => \N__6930\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__6949\,
            I => \N__6927\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__6946\,
            I => \N__6920\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__6943\,
            I => \N__6920\
        );

    \I__1416\ : Span4Mux_h
    port map (
            O => \N__6940\,
            I => \N__6920\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6913\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6913\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6933\,
            I => \N__6913\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6930\,
            I => \U712_CHIP_RAM.N_275\
        );

    \I__1411\ : Odrv4
    port map (
            O => \N__6927\,
            I => \U712_CHIP_RAM.N_275\
        );

    \I__1410\ : Odrv4
    port map (
            O => \N__6920\,
            I => \U712_CHIP_RAM.N_275\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__6913\,
            I => \U712_CHIP_RAM.N_275\
        );

    \I__1408\ : InMux
    port map (
            O => \N__6904\,
            I => \N__6901\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__6901\,
            I => \N__6898\
        );

    \I__1406\ : Span4Mux_h
    port map (
            O => \N__6898\,
            I => \N__6895\
        );

    \I__1405\ : Odrv4
    port map (
            O => \N__6895\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_0_a2_0_0\
        );

    \I__1404\ : InMux
    port map (
            O => \N__6892\,
            I => \N__6889\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__6889\,
            I => \N__6885\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6888\,
            I => \N__6881\
        );

    \I__1401\ : Span4Mux_h
    port map (
            O => \N__6885\,
            I => \N__6878\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6884\,
            I => \N__6875\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__6881\,
            I => \N__6872\
        );

    \I__1398\ : Odrv4
    port map (
            O => \N__6878\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_0_a2_0\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__6875\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_0_a2_0\
        );

    \I__1396\ : Odrv4
    port map (
            O => \N__6872\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_0_a2_0\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__6865\,
            I => \U712_CHIP_RAM.N_375_cascade_\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__6862\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_cascade_\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6859\,
            I => \N__6855\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6858\,
            I => \N__6852\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6855\,
            I => \N__6846\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6852\,
            I => \N__6840\
        );

    \I__1389\ : InMux
    port map (
            O => \N__6851\,
            I => \N__6833\
        );

    \I__1388\ : InMux
    port map (
            O => \N__6850\,
            I => \N__6833\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6833\
        );

    \I__1386\ : Span4Mux_v
    port map (
            O => \N__6846\,
            I => \N__6830\
        );

    \I__1385\ : InMux
    port map (
            O => \N__6845\,
            I => \N__6825\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6844\,
            I => \N__6825\
        );

    \I__1383\ : InMux
    port map (
            O => \N__6843\,
            I => \N__6822\
        );

    \I__1382\ : Odrv4
    port map (
            O => \N__6840\,
            I => \U712_CHIP_RAM.N_263\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__6833\,
            I => \U712_CHIP_RAM.N_263\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__6830\,
            I => \U712_CHIP_RAM.N_263\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6825\,
            I => \U712_CHIP_RAM.N_263\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6822\,
            I => \U712_CHIP_RAM.N_263\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6811\,
            I => \N__6808\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__6808\,
            I => \N__6801\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6807\,
            I => \N__6798\
        );

    \I__1374\ : CascadeMux
    port map (
            O => \N__6806\,
            I => \N__6791\
        );

    \I__1373\ : InMux
    port map (
            O => \N__6805\,
            I => \N__6786\
        );

    \I__1372\ : InMux
    port map (
            O => \N__6804\,
            I => \N__6783\
        );

    \I__1371\ : Span4Mux_h
    port map (
            O => \N__6801\,
            I => \N__6780\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__6798\,
            I => \N__6777\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6797\,
            I => \N__6774\
        );

    \I__1368\ : InMux
    port map (
            O => \N__6796\,
            I => \N__6767\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6795\,
            I => \N__6767\
        );

    \I__1366\ : InMux
    port map (
            O => \N__6794\,
            I => \N__6767\
        );

    \I__1365\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6760\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6790\,
            I => \N__6760\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6789\,
            I => \N__6760\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__6786\,
            I => \N__6757\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6783\,
            I => \U712_CHIP_RAM.N_267\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__6780\,
            I => \U712_CHIP_RAM.N_267\
        );

    \I__1359\ : Odrv4
    port map (
            O => \N__6777\,
            I => \U712_CHIP_RAM.N_267\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__6774\,
            I => \U712_CHIP_RAM.N_267\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__6767\,
            I => \U712_CHIP_RAM.N_267\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__6760\,
            I => \U712_CHIP_RAM.N_267\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__6757\,
            I => \U712_CHIP_RAM.N_267\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__6742\,
            I => \N__6737\
        );

    \I__1353\ : InMux
    port map (
            O => \N__6741\,
            I => \N__6734\
        );

    \I__1352\ : InMux
    port map (
            O => \N__6740\,
            I => \N__6731\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6728\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6734\,
            I => \U712_CHIP_RAM.N_270\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6731\,
            I => \U712_CHIP_RAM.N_270\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__6728\,
            I => \U712_CHIP_RAM.N_270\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6721\,
            I => \N__6718\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__6718\,
            I => \N__6713\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6717\,
            I => \N__6708\
        );

    \I__1344\ : InMux
    port map (
            O => \N__6716\,
            I => \N__6708\
        );

    \I__1343\ : Span4Mux_v
    port map (
            O => \N__6713\,
            I => \N__6702\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6708\,
            I => \N__6702\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6707\,
            I => \N__6697\
        );

    \I__1340\ : Span4Mux_h
    port map (
            O => \N__6702\,
            I => \N__6694\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6701\,
            I => \N__6689\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6700\,
            I => \N__6689\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6697\,
            I => \U712_CHIP_RAM.N_289\
        );

    \I__1336\ : Odrv4
    port map (
            O => \N__6694\,
            I => \U712_CHIP_RAM.N_289\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__6689\,
            I => \U712_CHIP_RAM.N_289\
        );

    \I__1334\ : CEMux
    port map (
            O => \N__6682\,
            I => \N__6679\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__6679\,
            I => \N__6676\
        );

    \I__1332\ : Odrv12
    port map (
            O => \N__6676\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_0\
        );

    \I__1331\ : InMux
    port map (
            O => \N__6673\,
            I => \N__6670\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__6670\,
            I => \N__6667\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__6667\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_3\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__6664\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0_i_0_cascade_\
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__6661\,
            I => \N__6654\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6660\,
            I => \N__6642\
        );

    \I__1325\ : InMux
    port map (
            O => \N__6659\,
            I => \N__6642\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6658\,
            I => \N__6637\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6657\,
            I => \N__6637\
        );

    \I__1322\ : InMux
    port map (
            O => \N__6654\,
            I => \N__6634\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6631\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6652\,
            I => \N__6624\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6624\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6650\,
            I => \N__6624\
        );

    \I__1317\ : InMux
    port map (
            O => \N__6649\,
            I => \N__6617\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6648\,
            I => \N__6617\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6647\,
            I => \N__6617\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__6642\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6637\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6634\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__6631\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__6624\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6617\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1308\ : CascadeMux
    port map (
            O => \N__6604\,
            I => \U712_CHIP_RAM.N_275_cascade_\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__6601\,
            I => \N__6596\
        );

    \I__1306\ : InMux
    port map (
            O => \N__6600\,
            I => \N__6593\
        );

    \I__1305\ : InMux
    port map (
            O => \N__6599\,
            I => \N__6590\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6583\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6593\,
            I => \N__6578\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__6590\,
            I => \N__6567\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6589\,
            I => \N__6564\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6588\,
            I => \N__6557\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6587\,
            I => \N__6557\
        );

    \I__1298\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6557\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6583\,
            I => \N__6554\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6549\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6581\,
            I => \N__6549\
        );

    \I__1294\ : Span4Mux_h
    port map (
            O => \N__6578\,
            I => \N__6546\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6543\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6538\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6575\,
            I => \N__6538\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6574\,
            I => \N__6531\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6573\,
            I => \N__6531\
        );

    \I__1288\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6531\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6526\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6570\,
            I => \N__6526\
        );

    \I__1285\ : Odrv4
    port map (
            O => \N__6567\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__6564\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6557\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1282\ : Odrv4
    port map (
            O => \N__6554\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6549\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1280\ : Odrv4
    port map (
            O => \N__6546\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6543\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__6538\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6531\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__6526\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__6505\,
            I => \U712_CHIP_RAM.N_423_cascade_\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6502\,
            I => \N__6498\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6501\,
            I => \N__6495\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6498\,
            I => \U712_CHIP_RAM.N_265\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__6495\,
            I => \U712_CHIP_RAM.N_265\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6490\,
            I => \N__6486\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6489\,
            I => \N__6483\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6486\,
            I => \U712_CHIP_RAM.N_303\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__6483\,
            I => \U712_CHIP_RAM.N_303\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6475\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6475\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a3_0_0\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6472\,
            I => \N__6469\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__6469\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGURED_e_1\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6466\,
            I => \N__6462\
        );

    \I__1261\ : InMux
    port map (
            O => \N__6465\,
            I => \N__6459\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6462\,
            I => \U712_CHIP_RAM.N_276_i\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6459\,
            I => \U712_CHIP_RAM.N_276_i\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6454\,
            I => \N__6450\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6453\,
            I => \N__6447\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__6450\,
            I => \N__6444\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__6447\,
            I => \N__6441\
        );

    \I__1254\ : Span4Mux_v
    port map (
            O => \N__6444\,
            I => \N__6438\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__6441\,
            I => \N__6435\
        );

    \I__1252\ : Span4Mux_v
    port map (
            O => \N__6438\,
            I => \N__6432\
        );

    \I__1251\ : Span4Mux_v
    port map (
            O => \N__6435\,
            I => \N__6429\
        );

    \I__1250\ : Sp12to4
    port map (
            O => \N__6432\,
            I => \N__6426\
        );

    \I__1249\ : Sp12to4
    port map (
            O => \N__6429\,
            I => \N__6423\
        );

    \I__1248\ : Span12Mux_h
    port map (
            O => \N__6426\,
            I => \N__6420\
        );

    \I__1247\ : Span12Mux_h
    port map (
            O => \N__6423\,
            I => \N__6417\
        );

    \I__1246\ : Odrv12
    port map (
            O => \N__6420\,
            I => \DRA_c_6\
        );

    \I__1245\ : Odrv12
    port map (
            O => \N__6417\,
            I => \DRA_c_6\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6412\,
            I => \N__6409\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__6409\,
            I => \N__6406\
        );

    \I__1242\ : Odrv4
    port map (
            O => \N__6406\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6403\,
            I => \N__6400\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__6400\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6394\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6394\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__6391\,
            I => \N__6387\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6384\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6387\,
            I => \N__6379\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6384\,
            I => \N__6376\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6383\,
            I => \N__6373\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6382\,
            I => \N__6370\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__6379\,
            I => \U712_CHIP_RAM.N_336\
        );

    \I__1230\ : Odrv4
    port map (
            O => \N__6376\,
            I => \U712_CHIP_RAM.N_336\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__6373\,
            I => \U712_CHIP_RAM.N_336\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__6370\,
            I => \U712_CHIP_RAM.N_336\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6361\,
            I => \N__6358\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6358\,
            I => \N__6355\
        );

    \I__1225\ : Odrv4
    port map (
            O => \N__6355\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_1\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__6352\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_1_cascade_\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6346\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__6346\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_3_1\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__6343\,
            I => \N__6340\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6340\,
            I => \N__6337\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6337\,
            I => \N__6334\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__6334\,
            I => \U712_CHIP_RAM.N_369\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6331\,
            I => \N__6328\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__6328\,
            I => \N__6324\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6321\
        );

    \I__1214\ : Odrv12
    port map (
            O => \N__6324\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c2\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__6321\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c2\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__6316\,
            I => \N__6313\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6308\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6303\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6303\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__6308\,
            I => \U712_CHIP_RAM.DMA_CYCLE_START_RNIQU7BEZ0\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6303\,
            I => \U712_CHIP_RAM.DMA_CYCLE_START_RNIQU7BEZ0\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6295\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6295\,
            I => \U712_CHIP_RAM.N_307\
        );

    \I__1204\ : IoInMux
    port map (
            O => \N__6292\,
            I => \N__6289\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6289\,
            I => \N__6286\
        );

    \I__1202\ : Odrv12
    port map (
            O => \N__6286\,
            I => \CMA_c_1\
        );

    \I__1201\ : IoInMux
    port map (
            O => \N__6283\,
            I => \N__6280\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6280\,
            I => \N__6277\
        );

    \I__1199\ : Span4Mux_s2_v
    port map (
            O => \N__6277\,
            I => \N__6274\
        );

    \I__1198\ : Span4Mux_v
    port map (
            O => \N__6274\,
            I => \N__6271\
        );

    \I__1197\ : Span4Mux_v
    port map (
            O => \N__6271\,
            I => \N__6268\
        );

    \I__1196\ : Span4Mux_h
    port map (
            O => \N__6268\,
            I => \N__6265\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__6265\,
            I => \CMA_c_10\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6262\,
            I => \N__6259\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6259\,
            I => \U712_CHIP_RAM.N_311\
        );

    \I__1192\ : IoInMux
    port map (
            O => \N__6256\,
            I => \N__6253\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__6253\,
            I => \N__6250\
        );

    \I__1190\ : Span12Mux_s4_h
    port map (
            O => \N__6250\,
            I => \N__6247\
        );

    \I__1189\ : Span12Mux_h
    port map (
            O => \N__6247\,
            I => \N__6244\
        );

    \I__1188\ : Odrv12
    port map (
            O => \N__6244\,
            I => \CMA_c_5\
        );

    \I__1187\ : IoInMux
    port map (
            O => \N__6241\,
            I => \N__6238\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6238\,
            I => \N__6235\
        );

    \I__1185\ : IoSpan4Mux
    port map (
            O => \N__6235\,
            I => \N__6232\
        );

    \I__1184\ : Span4Mux_s2_v
    port map (
            O => \N__6232\,
            I => \N__6229\
        );

    \I__1183\ : Span4Mux_v
    port map (
            O => \N__6229\,
            I => \N__6226\
        );

    \I__1182\ : Span4Mux_v
    port map (
            O => \N__6226\,
            I => \N__6223\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__6223\,
            I => \CMA_c_0\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6220\,
            I => \N__6217\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6217\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6211\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6211\,
            I => \N__6208\
        );

    \I__1176\ : Span12Mux_v
    port map (
            O => \N__6208\,
            I => \N__6205\
        );

    \I__1175\ : Span12Mux_h
    port map (
            O => \N__6205\,
            I => \N__6202\
        );

    \I__1174\ : Odrv12
    port map (
            O => \N__6202\,
            I => \A_c_15\
        );

    \I__1173\ : CascadeMux
    port map (
            O => \N__6199\,
            I => \N__6196\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6196\,
            I => \N__6193\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6193\,
            I => \N__6190\
        );

    \I__1170\ : Span4Mux_v
    port map (
            O => \N__6190\,
            I => \N__6187\
        );

    \I__1169\ : Span4Mux_v
    port map (
            O => \N__6187\,
            I => \N__6184\
        );

    \I__1168\ : Sp12to4
    port map (
            O => \N__6184\,
            I => \N__6181\
        );

    \I__1167\ : Span12Mux_h
    port map (
            O => \N__6181\,
            I => \N__6178\
        );

    \I__1166\ : Odrv12
    port map (
            O => \N__6178\,
            I => \A_c_8\
        );

    \I__1165\ : InMux
    port map (
            O => \N__6175\,
            I => \N__6172\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__6172\,
            I => \U712_CHIP_RAM.N_312\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6169\,
            I => \N__6166\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__6166\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6163\,
            I => \N__6160\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__6160\,
            I => \N__6157\
        );

    \I__1159\ : Span12Mux_v
    port map (
            O => \N__6157\,
            I => \N__6154\
        );

    \I__1158\ : Span12Mux_h
    port map (
            O => \N__6154\,
            I => \N__6151\
        );

    \I__1157\ : Odrv12
    port map (
            O => \N__6151\,
            I => \A_c_9\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__6148\,
            I => \N__6145\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6145\,
            I => \N__6142\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6142\,
            I => \N__6139\
        );

    \I__1153\ : Span12Mux_v
    port map (
            O => \N__6139\,
            I => \N__6136\
        );

    \I__1152\ : Span12Mux_h
    port map (
            O => \N__6136\,
            I => \N__6133\
        );

    \I__1151\ : Span12Mux_v
    port map (
            O => \N__6133\,
            I => \N__6130\
        );

    \I__1150\ : Odrv12
    port map (
            O => \N__6130\,
            I => \A_c_2\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6127\,
            I => \N__6124\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6124\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__6121\,
            I => \N__6118\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6118\,
            I => \N__6115\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6115\,
            I => \U712_CHIP_RAM.N_306\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6112\,
            I => \N__6109\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6109\,
            I => \N__6105\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6108\,
            I => \N__6102\
        );

    \I__1141\ : Sp12to4
    port map (
            O => \N__6105\,
            I => \N__6097\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__6102\,
            I => \N__6097\
        );

    \I__1139\ : Span12Mux_v
    port map (
            O => \N__6097\,
            I => \N__6094\
        );

    \I__1138\ : Span12Mux_h
    port map (
            O => \N__6094\,
            I => \N__6091\
        );

    \I__1137\ : Odrv12
    port map (
            O => \N__6091\,
            I => \DRA_c_4\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6085\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6085\,
            I => \N__6082\
        );

    \I__1134\ : Odrv12
    port map (
            O => \N__6082\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6079\,
            I => \N__6072\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6072\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6069\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__6072\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6069\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6064\,
            I => \N__6058\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6063\,
            I => \N__6058\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6058\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__1125\ : IoInMux
    port map (
            O => \N__6055\,
            I => \N__6052\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6052\,
            I => \N__6049\
        );

    \I__1123\ : Span12Mux_s7_v
    port map (
            O => \N__6049\,
            I => \N__6046\
        );

    \I__1122\ : Span12Mux_h
    port map (
            O => \N__6046\,
            I => \N__6043\
        );

    \I__1121\ : Odrv12
    port map (
            O => \N__6043\,
            I => \U712_REG_SM_un1_UDSn_i\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6040\,
            I => \N__6036\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6039\,
            I => \N__6032\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6036\,
            I => \N__6029\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6026\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6032\,
            I => \N__6022\
        );

    \I__1115\ : Span4Mux_v
    port map (
            O => \N__6029\,
            I => \N__6019\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6026\,
            I => \N__6016\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6025\,
            I => \N__6013\
        );

    \I__1112\ : Span4Mux_v
    port map (
            O => \N__6022\,
            I => \N__6010\
        );

    \I__1111\ : Sp12to4
    port map (
            O => \N__6019\,
            I => \N__6001\
        );

    \I__1110\ : Sp12to4
    port map (
            O => \N__6016\,
            I => \N__6001\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6013\,
            I => \N__6001\
        );

    \I__1108\ : Sp12to4
    port map (
            O => \N__6010\,
            I => \N__6001\
        );

    \I__1107\ : Span12Mux_h
    port map (
            O => \N__6001\,
            I => \N__5998\
        );

    \I__1106\ : Span12Mux_v
    port map (
            O => \N__5998\,
            I => \N__5995\
        );

    \I__1105\ : Odrv12
    port map (
            O => \N__5995\,
            I => \RnW_c\
        );

    \I__1104\ : IoInMux
    port map (
            O => \N__5992\,
            I => \N__5989\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5989\,
            I => \N__5985\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__5988\,
            I => \N__5982\
        );

    \I__1101\ : Span12Mux_s1_v
    port map (
            O => \N__5985\,
            I => \N__5978\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5982\,
            I => \N__5975\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__5981\,
            I => \N__5972\
        );

    \I__1098\ : Span12Mux_v
    port map (
            O => \N__5978\,
            I => \N__5969\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5975\,
            I => \N__5966\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5963\
        );

    \I__1095\ : Odrv12
    port map (
            O => \N__5969\,
            I => \DBDIR_c\
        );

    \I__1094\ : Odrv12
    port map (
            O => \N__5966\,
            I => \DBDIR_c\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5963\,
            I => \DBDIR_c\
        );

    \I__1092\ : IoInMux
    port map (
            O => \N__5956\,
            I => \N__5953\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5953\,
            I => \N__5950\
        );

    \I__1090\ : Span12Mux_s7_h
    port map (
            O => \N__5950\,
            I => \N__5947\
        );

    \I__1089\ : Span12Mux_v
    port map (
            O => \N__5947\,
            I => \N__5944\
        );

    \I__1088\ : Odrv12
    port map (
            O => \N__5944\,
            I => \N_208\
        );

    \I__1087\ : IoInMux
    port map (
            O => \N__5941\,
            I => \N__5938\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5938\,
            I => \N__5935\
        );

    \I__1085\ : Span12Mux_s6_v
    port map (
            O => \N__5935\,
            I => \N__5932\
        );

    \I__1084\ : Odrv12
    port map (
            O => \N__5932\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5929\,
            I => \N__5926\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__5926\,
            I => \N__5923\
        );

    \I__1081\ : Span4Mux_h
    port map (
            O => \N__5923\,
            I => \N__5920\
        );

    \I__1080\ : Odrv4
    port map (
            O => \N__5920\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5917\,
            I => \N__5914\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__5914\,
            I => \N__5911\
        );

    \I__1077\ : Span4Mux_v
    port map (
            O => \N__5911\,
            I => \N__5908\
        );

    \I__1076\ : Sp12to4
    port map (
            O => \N__5908\,
            I => \N__5905\
        );

    \I__1075\ : Span12Mux_h
    port map (
            O => \N__5905\,
            I => \N__5902\
        );

    \I__1074\ : Odrv12
    port map (
            O => \N__5902\,
            I => \A_c_10\
        );

    \I__1073\ : CascadeMux
    port map (
            O => \N__5899\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_\
        );

    \I__1072\ : InMux
    port map (
            O => \N__5896\,
            I => \N__5893\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__5893\,
            I => \N__5890\
        );

    \I__1070\ : Span4Mux_v
    port map (
            O => \N__5890\,
            I => \N__5887\
        );

    \I__1069\ : Sp12to4
    port map (
            O => \N__5887\,
            I => \N__5884\
        );

    \I__1068\ : Span12Mux_h
    port map (
            O => \N__5884\,
            I => \N__5881\
        );

    \I__1067\ : Span12Mux_v
    port map (
            O => \N__5881\,
            I => \N__5878\
        );

    \I__1066\ : Odrv12
    port map (
            O => \N__5878\,
            I => \A_c_3\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5872\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__5872\,
            I => \N__5869\
        );

    \I__1063\ : Odrv4
    port map (
            O => \N__5869\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5863\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5863\,
            I => \N__5860\
        );

    \I__1060\ : Span4Mux_v
    port map (
            O => \N__5860\,
            I => \N__5857\
        );

    \I__1059\ : Sp12to4
    port map (
            O => \N__5857\,
            I => \N__5854\
        );

    \I__1058\ : Span12Mux_h
    port map (
            O => \N__5854\,
            I => \N__5851\
        );

    \I__1057\ : Odrv12
    port map (
            O => \N__5851\,
            I => \A_c_14\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__5848\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5_cascade_\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5845\,
            I => \N__5842\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5842\,
            I => \N__5839\
        );

    \I__1053\ : Span4Mux_h
    port map (
            O => \N__5839\,
            I => \N__5836\
        );

    \I__1052\ : Span4Mux_v
    port map (
            O => \N__5836\,
            I => \N__5833\
        );

    \I__1051\ : Span4Mux_v
    port map (
            O => \N__5833\,
            I => \N__5830\
        );

    \I__1050\ : Sp12to4
    port map (
            O => \N__5830\,
            I => \N__5827\
        );

    \I__1049\ : Odrv12
    port map (
            O => \N__5827\,
            I => \A_c_7\
        );

    \I__1048\ : IoInMux
    port map (
            O => \N__5824\,
            I => \N__5821\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5821\,
            I => \N__5818\
        );

    \I__1046\ : IoSpan4Mux
    port map (
            O => \N__5818\,
            I => \N__5815\
        );

    \I__1045\ : Span4Mux_s3_h
    port map (
            O => \N__5815\,
            I => \N__5812\
        );

    \I__1044\ : Span4Mux_v
    port map (
            O => \N__5812\,
            I => \N__5809\
        );

    \I__1043\ : Span4Mux_h
    port map (
            O => \N__5809\,
            I => \N__5806\
        );

    \I__1042\ : Sp12to4
    port map (
            O => \N__5806\,
            I => \N__5803\
        );

    \I__1041\ : Odrv12
    port map (
            O => \N__5803\,
            I => \CMA_c_6\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__5800\,
            I => \N__5797\
        );

    \I__1039\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5790\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5796\,
            I => \N__5790\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5795\,
            I => \N__5787\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5790\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5787\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__1034\ : InMux
    port map (
            O => \N__5782\,
            I => \N__5778\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5781\,
            I => \N__5775\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5778\,
            I => \N__5770\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__5775\,
            I => \N__5767\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5774\,
            I => \N__5762\
        );

    \I__1029\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5762\
        );

    \I__1028\ : Odrv12
    port map (
            O => \N__5770\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1027\ : Odrv4
    port map (
            O => \N__5767\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__5762\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5755\,
            I => \N__5749\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5754\,
            I => \N__5746\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5753\,
            I => \N__5741\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5752\,
            I => \N__5741\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__5749\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5746\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5741\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1018\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5731\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5731\,
            I => \U712_REG_SM.DS_EN_RNOZ0Z_2\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__1015\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5722\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5722\,
            I => \N__5719\
        );

    \I__1013\ : Odrv4
    port map (
            O => \N__5719\,
            I => \U712_REG_SM.N_210\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5716\,
            I => \N__5713\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__5713\,
            I => \U712_REG_SM.N_355\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5710\,
            I => \N__5707\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__5707\,
            I => \N__5704\
        );

    \I__1008\ : Span4Mux_h
    port map (
            O => \N__5704\,
            I => \N__5698\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5693\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5702\,
            I => \N__5693\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5690\
        );

    \I__1004\ : Odrv4
    port map (
            O => \N__5698\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5693\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__5690\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__5683\,
            I => \N__5679\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5682\,
            I => \N__5673\
        );

    \I__999\ : InMux
    port map (
            O => \N__5679\,
            I => \N__5673\
        );

    \I__998\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5670\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5673\,
            I => \N__5667\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5670\,
            I => \U712_REG_SM.N_279\
        );

    \I__995\ : Odrv4
    port map (
            O => \N__5667\,
            I => \U712_REG_SM.N_279\
        );

    \I__994\ : InMux
    port map (
            O => \N__5662\,
            I => \N__5659\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5659\,
            I => \N__5656\
        );

    \I__992\ : Span4Mux_h
    port map (
            O => \N__5656\,
            I => \N__5651\
        );

    \I__991\ : InMux
    port map (
            O => \N__5655\,
            I => \N__5646\
        );

    \I__990\ : InMux
    port map (
            O => \N__5654\,
            I => \N__5646\
        );

    \I__989\ : Odrv4
    port map (
            O => \N__5651\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5646\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__5641\,
            I => \N__5638\
        );

    \I__986\ : InMux
    port map (
            O => \N__5638\,
            I => \N__5634\
        );

    \I__985\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5631\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5634\,
            I => \REG_TACK\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5631\,
            I => \REG_TACK\
        );

    \I__982\ : InMux
    port map (
            O => \N__5626\,
            I => \N__5623\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5623\,
            I => \N__5617\
        );

    \I__980\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5612\
        );

    \I__979\ : InMux
    port map (
            O => \N__5621\,
            I => \N__5612\
        );

    \I__978\ : InMux
    port map (
            O => \N__5620\,
            I => \N__5609\
        );

    \I__977\ : Span4Mux_h
    port map (
            O => \N__5617\,
            I => \N__5606\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5612\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__5609\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__974\ : Odrv4
    port map (
            O => \N__5606\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__973\ : InMux
    port map (
            O => \N__5599\,
            I => \N__5592\
        );

    \I__972\ : InMux
    port map (
            O => \N__5598\,
            I => \N__5592\
        );

    \I__971\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5589\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5592\,
            I => \U712_REG_SM.N_301\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__5589\,
            I => \U712_REG_SM.N_301\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__5584\,
            I => \U712_REG_SM.N_302_cascade_\
        );

    \I__967\ : InMux
    port map (
            O => \N__5581\,
            I => \N__5575\
        );

    \I__966\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5575\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__5575\,
            I => \N__5572\
        );

    \I__964\ : Odrv12
    port map (
            O => \N__5572\,
            I => \U712_REG_SM.LDS_OUT_2_0_a2_0_a2Z0Z_0\
        );

    \I__963\ : InMux
    port map (
            O => \N__5569\,
            I => \N__5562\
        );

    \I__962\ : InMux
    port map (
            O => \N__5568\,
            I => \N__5562\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__5567\,
            I => \N__5558\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__5562\,
            I => \N__5553\
        );

    \I__959\ : InMux
    port map (
            O => \N__5561\,
            I => \N__5548\
        );

    \I__958\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5548\
        );

    \I__957\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5543\
        );

    \I__956\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5543\
        );

    \I__955\ : Span4Mux_h
    port map (
            O => \N__5553\,
            I => \N__5540\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5548\,
            I => \N__5535\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5543\,
            I => \N__5535\
        );

    \I__952\ : Span4Mux_v
    port map (
            O => \N__5540\,
            I => \N__5532\
        );

    \I__951\ : Sp12to4
    port map (
            O => \N__5535\,
            I => \N__5529\
        );

    \I__950\ : Sp12to4
    port map (
            O => \N__5532\,
            I => \N__5524\
        );

    \I__949\ : Span12Mux_v
    port map (
            O => \N__5529\,
            I => \N__5524\
        );

    \I__948\ : Odrv12
    port map (
            O => \N__5524\,
            I => \A_c_0\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__5521\,
            I => \N__5518\
        );

    \I__946\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5515\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__5515\,
            I => \U712_REG_SM.N_302\
        );

    \I__944\ : InMux
    port map (
            O => \N__5512\,
            I => \N__5506\
        );

    \I__943\ : InMux
    port map (
            O => \N__5511\,
            I => \N__5506\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5506\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__941\ : IoInMux
    port map (
            O => \N__5503\,
            I => \N__5500\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5500\,
            I => \N__5497\
        );

    \I__939\ : Span4Mux_s2_v
    port map (
            O => \N__5497\,
            I => \N__5494\
        );

    \I__938\ : Sp12to4
    port map (
            O => \N__5494\,
            I => \N__5491\
        );

    \I__937\ : Span12Mux_h
    port map (
            O => \N__5491\,
            I => \N__5488\
        );

    \I__936\ : Span12Mux_v
    port map (
            O => \N__5488\,
            I => \N__5485\
        );

    \I__935\ : Odrv12
    port map (
            O => \N__5485\,
            I => \U712_REG_SM_un1_LDSn_i\
        );

    \I__934\ : InMux
    port map (
            O => \N__5482\,
            I => \N__5479\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__5479\,
            I => \N__5476\
        );

    \I__932\ : Span4Mux_v
    port map (
            O => \N__5476\,
            I => \N__5473\
        );

    \I__931\ : Odrv4
    port map (
            O => \N__5473\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1\
        );

    \I__930\ : InMux
    port map (
            O => \N__5470\,
            I => \N__5467\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5467\,
            I => \N__5464\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__5464\,
            I => \U712_CHIP_RAM.N_427\
        );

    \I__927\ : InMux
    port map (
            O => \N__5461\,
            I => \N__5458\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5458\,
            I => \CPU_TACKm\
        );

    \I__925\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5450\
        );

    \I__924\ : InMux
    port map (
            O => \N__5454\,
            I => \N__5447\
        );

    \I__923\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5444\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__5450\,
            I => \N__5437\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__5447\,
            I => \N__5437\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__5444\,
            I => \N__5437\
        );

    \I__919\ : Odrv12
    port map (
            O => \N__5437\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__918\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5430\
        );

    \I__917\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5427\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5430\,
            I => \N__5424\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__5427\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__914\ : Odrv12
    port map (
            O => \N__5424\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__5419\,
            I => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__5416\,
            I => \N__5412\
        );

    \I__911\ : InMux
    port map (
            O => \N__5415\,
            I => \N__5408\
        );

    \I__910\ : InMux
    port map (
            O => \N__5412\,
            I => \N__5405\
        );

    \I__909\ : InMux
    port map (
            O => \N__5411\,
            I => \N__5402\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__5408\,
            I => \N__5399\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5405\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5402\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__905\ : Odrv4
    port map (
            O => \N__5399\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__5392\,
            I => \U712_CYCLE_TERM.N_298_i_0_en_cascade_\
        );

    \I__903\ : CEMux
    port map (
            O => \N__5389\,
            I => \N__5386\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5386\,
            I => \N__5383\
        );

    \I__901\ : Odrv12
    port map (
            O => \N__5383\,
            I => \U712_CYCLE_TERM.N_298_i_0_en_0\
        );

    \I__900\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5373\
        );

    \I__899\ : InMux
    port map (
            O => \N__5379\,
            I => \N__5373\
        );

    \I__898\ : InMux
    port map (
            O => \N__5378\,
            I => \N__5370\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5373\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5370\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__5365\,
            I => \N__5362\
        );

    \I__894\ : InMux
    port map (
            O => \N__5362\,
            I => \N__5358\
        );

    \I__893\ : InMux
    port map (
            O => \N__5361\,
            I => \N__5355\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5358\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__5355\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__5350\,
            I => \N__5347\
        );

    \I__889\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5342\
        );

    \I__888\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5339\
        );

    \I__887\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5336\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5342\,
            I => \N__5333\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5339\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5336\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__883\ : Odrv4
    port map (
            O => \N__5333\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__882\ : InMux
    port map (
            O => \N__5326\,
            I => \N__5320\
        );

    \I__881\ : InMux
    port map (
            O => \N__5325\,
            I => \N__5313\
        );

    \I__880\ : InMux
    port map (
            O => \N__5324\,
            I => \N__5313\
        );

    \I__879\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5313\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__5320\,
            I => \N__5310\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5313\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__876\ : Odrv4
    port map (
            O => \N__5310\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__5305\,
            I => \U712_CHIP_RAM.N_267_cascade_\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__5302\,
            I => \U712_CHIP_RAM.N_204_cascade_\
        );

    \I__873\ : CEMux
    port map (
            O => \N__5299\,
            I => \N__5296\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5296\,
            I => \N__5293\
        );

    \I__871\ : Span4Mux_v
    port map (
            O => \N__5293\,
            I => \N__5290\
        );

    \I__870\ : Odrv4
    port map (
            O => \N__5290\,
            I => \U712_CHIP_RAM.N_204_0_0\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__5287\,
            I => \U712_CHIP_RAM.N_340_cascade_\
        );

    \I__868\ : InMux
    port map (
            O => \N__5284\,
            I => \N__5274\
        );

    \I__867\ : InMux
    port map (
            O => \N__5283\,
            I => \N__5274\
        );

    \I__866\ : InMux
    port map (
            O => \N__5282\,
            I => \N__5274\
        );

    \I__865\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5271\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5274\,
            I => \U712_CHIP_RAM.N_278\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5271\,
            I => \U712_CHIP_RAM.N_278\
        );

    \I__862\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5263\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5263\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_1_0\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__5260\,
            I => \U712_CHIP_RAM.N_417_cascade_\
        );

    \I__859\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5254\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5254\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__857\ : SRMux
    port map (
            O => \N__5251\,
            I => \N__5248\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__5248\,
            I => \N__5245\
        );

    \I__855\ : Span4Mux_h
    port map (
            O => \N__5245\,
            I => \N__5242\
        );

    \I__854\ : Odrv4
    port map (
            O => \N__5242\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__853\ : CascadeMux
    port map (
            O => \N__5239\,
            I => \U712_CHIP_RAM.REFRESH_RST_cascade_\
        );

    \I__852\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5233\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5233\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__5230\,
            I => \N__5227\
        );

    \I__849\ : InMux
    port map (
            O => \N__5227\,
            I => \N__5222\
        );

    \I__848\ : InMux
    port map (
            O => \N__5226\,
            I => \N__5217\
        );

    \I__847\ : InMux
    port map (
            O => \N__5225\,
            I => \N__5217\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5222\,
            I => \N__5212\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5217\,
            I => \N__5212\
        );

    \I__844\ : Odrv4
    port map (
            O => \N__5212\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__843\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5205\
        );

    \I__842\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5202\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5205\,
            I => \N__5197\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5202\,
            I => \N__5197\
        );

    \I__839\ : Span4Mux_v
    port map (
            O => \N__5197\,
            I => \N__5194\
        );

    \I__838\ : Sp12to4
    port map (
            O => \N__5194\,
            I => \N__5191\
        );

    \I__837\ : Span12Mux_h
    port map (
            O => \N__5191\,
            I => \N__5188\
        );

    \I__836\ : Span12Mux_v
    port map (
            O => \N__5188\,
            I => \N__5185\
        );

    \I__835\ : Odrv12
    port map (
            O => \N__5185\,
            I => \AWEn_c\
        );

    \I__834\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5179\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__5179\,
            I => \N__5175\
        );

    \I__832\ : IoInMux
    port map (
            O => \N__5178\,
            I => \N__5172\
        );

    \I__831\ : Span4Mux_v
    port map (
            O => \N__5175\,
            I => \N__5169\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5172\,
            I => \N__5166\
        );

    \I__829\ : Sp12to4
    port map (
            O => \N__5169\,
            I => \N__5163\
        );

    \I__828\ : Span4Mux_s3_h
    port map (
            O => \N__5166\,
            I => \N__5160\
        );

    \I__827\ : Span12Mux_h
    port map (
            O => \N__5163\,
            I => \N__5155\
        );

    \I__826\ : Sp12to4
    port map (
            O => \N__5160\,
            I => \N__5155\
        );

    \I__825\ : Span12Mux_v
    port map (
            O => \N__5155\,
            I => \N__5152\
        );

    \I__824\ : Odrv12
    port map (
            O => \N__5152\,
            I => \C1_c\
        );

    \I__823\ : InMux
    port map (
            O => \N__5149\,
            I => \N__5140\
        );

    \I__822\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5133\
        );

    \I__821\ : InMux
    port map (
            O => \N__5147\,
            I => \N__5133\
        );

    \I__820\ : InMux
    port map (
            O => \N__5146\,
            I => \N__5133\
        );

    \I__819\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5126\
        );

    \I__818\ : InMux
    port map (
            O => \N__5144\,
            I => \N__5126\
        );

    \I__817\ : InMux
    port map (
            O => \N__5143\,
            I => \N__5126\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5140\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__5133\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__5126\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__813\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5116\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5116\,
            I => \U712_CHIP_RAM.N_308\
        );

    \I__811\ : IoInMux
    port map (
            O => \N__5113\,
            I => \N__5110\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__5110\,
            I => \N__5107\
        );

    \I__809\ : Span12Mux_s8_v
    port map (
            O => \N__5107\,
            I => \N__5104\
        );

    \I__808\ : Odrv12
    port map (
            O => \N__5104\,
            I => \CMA_c_2\
        );

    \I__807\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5098\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5098\,
            I => \U712_CHIP_RAM.N_310\
        );

    \I__805\ : IoInMux
    port map (
            O => \N__5095\,
            I => \N__5092\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5092\,
            I => \N__5089\
        );

    \I__803\ : Span4Mux_s3_h
    port map (
            O => \N__5089\,
            I => \N__5086\
        );

    \I__802\ : Sp12to4
    port map (
            O => \N__5086\,
            I => \N__5083\
        );

    \I__801\ : Span12Mux_s10_v
    port map (
            O => \N__5083\,
            I => \N__5080\
        );

    \I__800\ : Span12Mux_h
    port map (
            O => \N__5080\,
            I => \N__5077\
        );

    \I__799\ : Odrv12
    port map (
            O => \N__5077\,
            I => \CMA_c_4\
        );

    \I__798\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5070\
        );

    \I__797\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5067\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5070\,
            I => \N__5064\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__5067\,
            I => \N__5061\
        );

    \I__794\ : Span4Mux_v
    port map (
            O => \N__5064\,
            I => \N__5058\
        );

    \I__793\ : Span4Mux_v
    port map (
            O => \N__5061\,
            I => \N__5055\
        );

    \I__792\ : Sp12to4
    port map (
            O => \N__5058\,
            I => \N__5052\
        );

    \I__791\ : Sp12to4
    port map (
            O => \N__5055\,
            I => \N__5049\
        );

    \I__790\ : Span12Mux_h
    port map (
            O => \N__5052\,
            I => \N__5046\
        );

    \I__789\ : Span12Mux_v
    port map (
            O => \N__5049\,
            I => \N__5043\
        );

    \I__788\ : Span12Mux_v
    port map (
            O => \N__5046\,
            I => \N__5040\
        );

    \I__787\ : Span12Mux_h
    port map (
            O => \N__5043\,
            I => \N__5037\
        );

    \I__786\ : Odrv12
    port map (
            O => \N__5040\,
            I => \DRA_c_0\
        );

    \I__785\ : Odrv12
    port map (
            O => \N__5037\,
            I => \DRA_c_0\
        );

    \I__784\ : InMux
    port map (
            O => \N__5032\,
            I => \N__5028\
        );

    \I__783\ : InMux
    port map (
            O => \N__5031\,
            I => \N__5025\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5028\,
            I => \N__5022\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5025\,
            I => \N__5019\
        );

    \I__780\ : Span4Mux_v
    port map (
            O => \N__5022\,
            I => \N__5016\
        );

    \I__779\ : Sp12to4
    port map (
            O => \N__5019\,
            I => \N__5013\
        );

    \I__778\ : Sp12to4
    port map (
            O => \N__5016\,
            I => \N__5010\
        );

    \I__777\ : Span12Mux_v
    port map (
            O => \N__5013\,
            I => \N__5007\
        );

    \I__776\ : Span12Mux_h
    port map (
            O => \N__5010\,
            I => \N__5004\
        );

    \I__775\ : Span12Mux_h
    port map (
            O => \N__5007\,
            I => \N__5001\
        );

    \I__774\ : Span12Mux_v
    port map (
            O => \N__5004\,
            I => \N__4998\
        );

    \I__773\ : Odrv12
    port map (
            O => \N__5001\,
            I => \DRA_c_2\
        );

    \I__772\ : Odrv12
    port map (
            O => \N__4998\,
            I => \DRA_c_2\
        );

    \I__771\ : InMux
    port map (
            O => \N__4993\,
            I => \N__4990\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4990\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__769\ : InMux
    port map (
            O => \N__4987\,
            I => \N__4984\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__4984\,
            I => \N__4980\
        );

    \I__767\ : InMux
    port map (
            O => \N__4983\,
            I => \N__4977\
        );

    \I__766\ : Span4Mux_h
    port map (
            O => \N__4980\,
            I => \N__4972\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4977\,
            I => \N__4972\
        );

    \I__764\ : Span4Mux_v
    port map (
            O => \N__4972\,
            I => \N__4969\
        );

    \I__763\ : Sp12to4
    port map (
            O => \N__4969\,
            I => \N__4966\
        );

    \I__762\ : Span12Mux_h
    port map (
            O => \N__4966\,
            I => \N__4963\
        );

    \I__761\ : Span12Mux_v
    port map (
            O => \N__4963\,
            I => \N__4960\
        );

    \I__760\ : Odrv12
    port map (
            O => \N__4960\,
            I => \DRA_c_3\
        );

    \I__759\ : InMux
    port map (
            O => \N__4957\,
            I => \N__4954\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4954\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__757\ : InMux
    port map (
            O => \N__4951\,
            I => \N__4948\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__4948\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__755\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4942\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__4942\,
            I => \N__4938\
        );

    \I__753\ : InMux
    port map (
            O => \N__4941\,
            I => \N__4935\
        );

    \I__752\ : Span4Mux_h
    port map (
            O => \N__4938\,
            I => \N__4930\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4935\,
            I => \N__4930\
        );

    \I__750\ : Span4Mux_h
    port map (
            O => \N__4930\,
            I => \N__4927\
        );

    \I__749\ : Sp12to4
    port map (
            O => \N__4927\,
            I => \N__4924\
        );

    \I__748\ : Span12Mux_v
    port map (
            O => \N__4924\,
            I => \N__4921\
        );

    \I__747\ : Span12Mux_h
    port map (
            O => \N__4921\,
            I => \N__4918\
        );

    \I__746\ : Odrv12
    port map (
            O => \N__4918\,
            I => \DRA_c_5\
        );

    \I__745\ : CascadeMux
    port map (
            O => \N__4915\,
            I => \N__4912\
        );

    \I__744\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4908\
        );

    \I__743\ : InMux
    port map (
            O => \N__4911\,
            I => \N__4904\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4908\,
            I => \N__4901\
        );

    \I__741\ : InMux
    port map (
            O => \N__4907\,
            I => \N__4898\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4904\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__739\ : Odrv12
    port map (
            O => \N__4901\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4898\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__4891\,
            I => \N__4887\
        );

    \I__736\ : InMux
    port map (
            O => \N__4890\,
            I => \N__4883\
        );

    \I__735\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4878\
        );

    \I__734\ : InMux
    port map (
            O => \N__4886\,
            I => \N__4878\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4883\,
            I => \U712_REG_SM.N_273\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4878\,
            I => \U712_REG_SM.N_273\
        );

    \I__731\ : InMux
    port map (
            O => \N__4873\,
            I => \N__4870\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4870\,
            I => \N__4867\
        );

    \I__729\ : Odrv4
    port map (
            O => \N__4867\,
            I => \U712_REG_SM.N_420\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__4864\,
            I => \N__4861\
        );

    \I__727\ : InMux
    port map (
            O => \N__4861\,
            I => \N__4856\
        );

    \I__726\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4853\
        );

    \I__725\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4850\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__4856\,
            I => \U712_REG_SM.N_491\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__4853\,
            I => \U712_REG_SM.N_491\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4850\,
            I => \U712_REG_SM.N_491\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__4843\,
            I => \U712_REG_SM.N_420_cascade_\
        );

    \I__720\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4835\
        );

    \I__719\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4832\
        );

    \I__718\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4829\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4835\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4832\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4829\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__4822\,
            I => \N__4817\
        );

    \I__713\ : InMux
    port map (
            O => \N__4821\,
            I => \N__4812\
        );

    \I__712\ : InMux
    port map (
            O => \N__4820\,
            I => \N__4805\
        );

    \I__711\ : InMux
    port map (
            O => \N__4817\,
            I => \N__4805\
        );

    \I__710\ : InMux
    port map (
            O => \N__4816\,
            I => \N__4805\
        );

    \I__709\ : InMux
    port map (
            O => \N__4815\,
            I => \N__4802\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4812\,
            I => \N__4799\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__4805\,
            I => \U712_REG_SM.N_281\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4802\,
            I => \U712_REG_SM.N_281\
        );

    \I__705\ : Odrv4
    port map (
            O => \N__4799\,
            I => \U712_REG_SM.N_281\
        );

    \I__704\ : CascadeMux
    port map (
            O => \N__4792\,
            I => \U712_REG_SM.N_281_cascade_\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__4789\,
            I => \N__4786\
        );

    \I__702\ : InMux
    port map (
            O => \N__4786\,
            I => \N__4782\
        );

    \I__701\ : InMux
    port map (
            O => \N__4785\,
            I => \N__4779\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4782\,
            I => \U712_REG_SM.N_300\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__4779\,
            I => \U712_REG_SM.N_300\
        );

    \I__698\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4762\
        );

    \I__697\ : InMux
    port map (
            O => \N__4773\,
            I => \N__4762\
        );

    \I__696\ : InMux
    port map (
            O => \N__4772\,
            I => \N__4762\
        );

    \I__695\ : InMux
    port map (
            O => \N__4771\,
            I => \N__4759\
        );

    \I__694\ : InMux
    port map (
            O => \N__4770\,
            I => \N__4754\
        );

    \I__693\ : InMux
    port map (
            O => \N__4769\,
            I => \N__4754\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4762\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__4759\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4754\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__689\ : CascadeMux
    port map (
            O => \N__4747\,
            I => \N__4744\
        );

    \I__688\ : InMux
    port map (
            O => \N__4744\,
            I => \N__4738\
        );

    \I__687\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4738\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4738\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__685\ : InMux
    port map (
            O => \N__4735\,
            I => \N__4731\
        );

    \I__684\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4728\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4731\,
            I => \U712_REG_SM.N_274\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__4728\,
            I => \U712_REG_SM.N_274\
        );

    \I__681\ : InMux
    port map (
            O => \N__4723\,
            I => \N__4717\
        );

    \I__680\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4717\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__4717\,
            I => \U712_REG_SM.N_282\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__4714\,
            I => \U712_REG_SM.N_274_cascade_\
        );

    \I__677\ : CascadeMux
    port map (
            O => \N__4711\,
            I => \N__4707\
        );

    \I__676\ : InMux
    port map (
            O => \N__4710\,
            I => \N__4703\
        );

    \I__675\ : InMux
    port map (
            O => \N__4707\,
            I => \N__4700\
        );

    \I__674\ : InMux
    port map (
            O => \N__4706\,
            I => \N__4697\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4703\,
            I => \U712_REG_SM.N_297\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4700\,
            I => \U712_REG_SM.N_297\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4697\,
            I => \U712_REG_SM.N_297\
        );

    \I__670\ : CascadeMux
    port map (
            O => \N__4690\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6_cascade_\
        );

    \I__669\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4684\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4684\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6\
        );

    \I__667\ : InMux
    port map (
            O => \N__4681\,
            I => \N__4677\
        );

    \I__666\ : InMux
    port map (
            O => \N__4680\,
            I => \N__4674\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4677\,
            I => \U712_REG_SM.N_492\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4674\,
            I => \U712_REG_SM.N_492\
        );

    \I__663\ : InMux
    port map (
            O => \N__4669\,
            I => \N__4660\
        );

    \I__662\ : InMux
    port map (
            O => \N__4668\,
            I => \N__4660\
        );

    \I__661\ : InMux
    port map (
            O => \N__4667\,
            I => \N__4660\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4660\,
            I => \N__4657\
        );

    \I__659\ : Odrv4
    port map (
            O => \N__4657\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c4\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__4654\,
            I => \U712_REG_SM.N_273_cascade_\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__4651\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_\
        );

    \I__656\ : CascadeMux
    port map (
            O => \N__4648\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_\
        );

    \I__655\ : CEMux
    port map (
            O => \N__4645\,
            I => \N__4642\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4642\,
            I => \N__4639\
        );

    \I__653\ : Odrv12
    port map (
            O => \N__4639\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__4636\,
            I => \N__4633\
        );

    \I__651\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4630\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4630\,
            I => \N__4627\
        );

    \I__649\ : Span4Mux_h
    port map (
            O => \N__4627\,
            I => \N__4623\
        );

    \I__648\ : InMux
    port map (
            O => \N__4626\,
            I => \N__4620\
        );

    \I__647\ : Odrv4
    port map (
            O => \N__4623\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__4620\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__645\ : InMux
    port map (
            O => \N__4615\,
            I => \N__4612\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4612\,
            I => \N__4609\
        );

    \I__643\ : Span12Mux_h
    port map (
            O => \N__4609\,
            I => \N__4606\
        );

    \I__642\ : Span12Mux_v
    port map (
            O => \N__4606\,
            I => \N__4603\
        );

    \I__641\ : Odrv12
    port map (
            O => \N__4603\,
            I => \DBRn_c\
        );

    \I__640\ : InMux
    port map (
            O => \N__4600\,
            I => \N__4597\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4597\,
            I => \N__4592\
        );

    \I__638\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4587\
        );

    \I__637\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4587\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__4592\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4587\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__634\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4577\
        );

    \I__633\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4574\
        );

    \I__632\ : InMux
    port map (
            O => \N__4580\,
            I => \N__4571\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4577\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4574\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__4571\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__628\ : InMux
    port map (
            O => \N__4564\,
            I => \N__4561\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__4561\,
            I => \U712_CHIP_RAM.N_139\
        );

    \I__626\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4555\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4555\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_1\
        );

    \I__624\ : CascadeMux
    port map (
            O => \N__4552\,
            I => \U712_CHIP_RAM.SDRAM_CMD_e_1_2_cascade_\
        );

    \I__623\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4545\
        );

    \I__622\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4542\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__4545\,
            I => \U712_CHIP_RAM.N_296\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__4542\,
            I => \U712_CHIP_RAM.N_296\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__4537\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c2_cascade_\
        );

    \I__618\ : CascadeMux
    port map (
            O => \N__4534\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_tz_0_cascade_\
        );

    \I__617\ : InMux
    port map (
            O => \N__4531\,
            I => \N__4522\
        );

    \I__616\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4522\
        );

    \I__615\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4522\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__4522\,
            I => \U712_REG_SM.N_292\
        );

    \I__613\ : InMux
    port map (
            O => \N__4519\,
            I => \N__4510\
        );

    \I__612\ : InMux
    port map (
            O => \N__4518\,
            I => \N__4510\
        );

    \I__611\ : InMux
    port map (
            O => \N__4517\,
            I => \N__4510\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4510\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__609\ : InMux
    port map (
            O => \N__4507\,
            I => \N__4504\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__4504\,
            I => \N__4501\
        );

    \I__607\ : Span12Mux_h
    port map (
            O => \N__4501\,
            I => \N__4498\
        );

    \I__606\ : Odrv12
    port map (
            O => \N__4498\,
            I => \A_c_13\
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__4495\,
            I => \N__4492\
        );

    \I__604\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4489\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__4489\,
            I => \N__4486\
        );

    \I__602\ : Span12Mux_v
    port map (
            O => \N__4486\,
            I => \N__4483\
        );

    \I__601\ : Span12Mux_h
    port map (
            O => \N__4483\,
            I => \N__4480\
        );

    \I__600\ : Odrv12
    port map (
            O => \N__4480\,
            I => \A_c_6\
        );

    \I__599\ : InMux
    port map (
            O => \N__4477\,
            I => \N__4474\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__4474\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__597\ : InMux
    port map (
            O => \N__4471\,
            I => \N__4468\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__4468\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4\
        );

    \I__595\ : CascadeMux
    port map (
            O => \N__4465\,
            I => \N__4462\
        );

    \I__594\ : InMux
    port map (
            O => \N__4462\,
            I => \N__4459\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4459\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__592\ : InMux
    port map (
            O => \N__4456\,
            I => \N__4453\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4453\,
            I => \N__4450\
        );

    \I__590\ : Span12Mux_v
    port map (
            O => \N__4450\,
            I => \N__4447\
        );

    \I__589\ : Span12Mux_h
    port map (
            O => \N__4447\,
            I => \N__4444\
        );

    \I__588\ : Odrv12
    port map (
            O => \N__4444\,
            I => \A_c_4\
        );

    \I__587\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4438\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4438\,
            I => \N__4435\
        );

    \I__585\ : Span12Mux_h
    port map (
            O => \N__4435\,
            I => \N__4432\
        );

    \I__584\ : Odrv12
    port map (
            O => \N__4432\,
            I => \A_c_11\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__4429\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_\
        );

    \I__582\ : InMux
    port map (
            O => \N__4426\,
            I => \N__4423\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__4423\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_2_0\
        );

    \I__580\ : InMux
    port map (
            O => \N__4420\,
            I => \N__4417\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__4417\,
            I => \N__4414\
        );

    \I__578\ : Span4Mux_v
    port map (
            O => \N__4414\,
            I => \N__4411\
        );

    \I__577\ : Sp12to4
    port map (
            O => \N__4411\,
            I => \N__4408\
        );

    \I__576\ : Span12Mux_h
    port map (
            O => \N__4408\,
            I => \N__4405\
        );

    \I__575\ : Odrv12
    port map (
            O => \N__4405\,
            I => \A_c_12\
        );

    \I__574\ : CascadeMux
    port map (
            O => \N__4402\,
            I => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_\
        );

    \I__573\ : InMux
    port map (
            O => \N__4399\,
            I => \N__4396\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4396\,
            I => \N__4393\
        );

    \I__571\ : Span4Mux_v
    port map (
            O => \N__4393\,
            I => \N__4390\
        );

    \I__570\ : Span4Mux_v
    port map (
            O => \N__4390\,
            I => \N__4387\
        );

    \I__569\ : Sp12to4
    port map (
            O => \N__4387\,
            I => \N__4384\
        );

    \I__568\ : Span12Mux_h
    port map (
            O => \N__4384\,
            I => \N__4381\
        );

    \I__567\ : Odrv12
    port map (
            O => \N__4381\,
            I => \A_c_5\
        );

    \I__566\ : InMux
    port map (
            O => \N__4378\,
            I => \N__4372\
        );

    \I__565\ : InMux
    port map (
            O => \N__4377\,
            I => \N__4372\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4372\,
            I => \N__4369\
        );

    \I__563\ : Odrv4
    port map (
            O => \N__4369\,
            I => \U712_REG_SM.N_295\
        );

    \I__562\ : CascadeMux
    port map (
            O => \N__4366\,
            I => \N__4362\
        );

    \I__561\ : CascadeMux
    port map (
            O => \N__4365\,
            I => \N__4359\
        );

    \I__560\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4356\
        );

    \I__559\ : InMux
    port map (
            O => \N__4359\,
            I => \N__4353\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__4356\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__4353\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__556\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4345\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4345\,
            I => \N__4342\
        );

    \I__554\ : Span12Mux_h
    port map (
            O => \N__4342\,
            I => \N__4339\
        );

    \I__553\ : Span12Mux_v
    port map (
            O => \N__4339\,
            I => \N__4336\
        );

    \I__552\ : Odrv12
    port map (
            O => \N__4336\,
            I => \C3_c\
        );

    \I__551\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4330\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4330\,
            I => \U712_REG_SM.N_338\
        );

    \I__549\ : CascadeMux
    port map (
            O => \N__4327\,
            I => \N__4324\
        );

    \I__548\ : InMux
    port map (
            O => \N__4324\,
            I => \N__4321\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4321\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_2_1_0\
        );

    \I__546\ : InMux
    port map (
            O => \N__4318\,
            I => \N__4312\
        );

    \I__545\ : InMux
    port map (
            O => \N__4317\,
            I => \N__4312\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4312\,
            I => \N__4309\
        );

    \I__543\ : Odrv4
    port map (
            O => \N__4309\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0Z0Z_0\
        );

    \I__542\ : InMux
    port map (
            O => \N__4306\,
            I => \N__4302\
        );

    \I__541\ : InMux
    port map (
            O => \N__4305\,
            I => \N__4299\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4302\,
            I => \N__4296\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__4299\,
            I => \N__4293\
        );

    \I__538\ : Span4Mux_h
    port map (
            O => \N__4296\,
            I => \N__4290\
        );

    \I__537\ : Span12Mux_h
    port map (
            O => \N__4293\,
            I => \N__4287\
        );

    \I__536\ : Sp12to4
    port map (
            O => \N__4290\,
            I => \N__4284\
        );

    \I__535\ : Span12Mux_v
    port map (
            O => \N__4287\,
            I => \N__4281\
        );

    \I__534\ : Span12Mux_v
    port map (
            O => \N__4284\,
            I => \N__4278\
        );

    \I__533\ : Odrv12
    port map (
            O => \N__4281\,
            I => \TSn_c\
        );

    \I__532\ : Odrv12
    port map (
            O => \N__4278\,
            I => \TSn_c\
        );

    \I__531\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4270\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__4270\,
            I => \N__4266\
        );

    \I__529\ : IoInMux
    port map (
            O => \N__4269\,
            I => \N__4263\
        );

    \I__528\ : Span12Mux_h
    port map (
            O => \N__4266\,
            I => \N__4260\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4263\,
            I => \N__4257\
        );

    \I__526\ : Span12Mux_v
    port map (
            O => \N__4260\,
            I => \N__4254\
        );

    \I__525\ : IoSpan4Mux
    port map (
            O => \N__4257\,
            I => \N__4251\
        );

    \I__524\ : Odrv12
    port map (
            O => \N__4254\,
            I => \RAMENn_c\
        );

    \I__523\ : Odrv4
    port map (
            O => \N__4251\,
            I => \RAMENn_c\
        );

    \I__522\ : InMux
    port map (
            O => \N__4246\,
            I => \N__4243\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4243\,
            I => \N__4240\
        );

    \I__520\ : Span4Mux_v
    port map (
            O => \N__4240\,
            I => \N__4237\
        );

    \I__519\ : Span4Mux_h
    port map (
            O => \N__4237\,
            I => \N__4234\
        );

    \I__518\ : Odrv4
    port map (
            O => \N__4234\,
            I => \TACK_EN_i_ess\
        );

    \I__517\ : IoInMux
    port map (
            O => \N__4231\,
            I => \N__4228\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4228\,
            I => \N__4224\
        );

    \I__515\ : IoInMux
    port map (
            O => \N__4227\,
            I => \N__4221\
        );

    \I__514\ : Span4Mux_s3_v
    port map (
            O => \N__4224\,
            I => \N__4218\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4221\,
            I => \N__4215\
        );

    \I__512\ : Span4Mux_h
    port map (
            O => \N__4218\,
            I => \N__4212\
        );

    \I__511\ : Span4Mux_s3_v
    port map (
            O => \N__4215\,
            I => \N__4209\
        );

    \I__510\ : Span4Mux_h
    port map (
            O => \N__4212\,
            I => \N__4206\
        );

    \I__509\ : Span4Mux_h
    port map (
            O => \N__4209\,
            I => \N__4203\
        );

    \I__508\ : Sp12to4
    port map (
            O => \N__4206\,
            I => \N__4200\
        );

    \I__507\ : Sp12to4
    port map (
            O => \N__4203\,
            I => \N__4197\
        );

    \I__506\ : Span12Mux_v
    port map (
            O => \N__4200\,
            I => \N__4191\
        );

    \I__505\ : Span12Mux_v
    port map (
            O => \N__4197\,
            I => \N__4191\
        );

    \I__504\ : InMux
    port map (
            O => \N__4196\,
            I => \N__4188\
        );

    \I__503\ : Odrv12
    port map (
            O => \N__4191\,
            I => \ASn_c\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4188\,
            I => \ASn_c\
        );

    \I__501\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4180\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4180\,
            I => \U712_BYTE_ENABLE.N_383\
        );

    \I__499\ : InMux
    port map (
            O => \N__4177\,
            I => \N__4174\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4174\,
            I => \U712_BYTE_ENABLE.N_379\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__4171\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_0_cascade_\
        );

    \I__496\ : IoInMux
    port map (
            O => \N__4168\,
            I => \N__4165\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4165\,
            I => \N__4162\
        );

    \I__494\ : Span4Mux_s3_h
    port map (
            O => \N__4162\,
            I => \N__4159\
        );

    \I__493\ : Span4Mux_v
    port map (
            O => \N__4159\,
            I => \N__4156\
        );

    \I__492\ : Sp12to4
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__491\ : Span12Mux_h
    port map (
            O => \N__4153\,
            I => \N__4150\
        );

    \I__490\ : Span12Mux_v
    port map (
            O => \N__4150\,
            I => \N__4147\
        );

    \I__489\ : Odrv12
    port map (
            O => \N__4147\,
            I => \N_48_i\
        );

    \I__488\ : InMux
    port map (
            O => \N__4144\,
            I => \N__4137\
        );

    \I__487\ : InMux
    port map (
            O => \N__4143\,
            I => \N__4137\
        );

    \I__486\ : CascadeMux
    port map (
            O => \N__4142\,
            I => \N__4134\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__4137\,
            I => \N__4131\
        );

    \I__484\ : InMux
    port map (
            O => \N__4134\,
            I => \N__4128\
        );

    \I__483\ : Span4Mux_v
    port map (
            O => \N__4131\,
            I => \N__4125\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4128\,
            I => \N__4122\
        );

    \I__481\ : Span4Mux_h
    port map (
            O => \N__4125\,
            I => \N__4119\
        );

    \I__480\ : Span4Mux_v
    port map (
            O => \N__4122\,
            I => \N__4116\
        );

    \I__479\ : Sp12to4
    port map (
            O => \N__4119\,
            I => \N__4111\
        );

    \I__478\ : Sp12to4
    port map (
            O => \N__4116\,
            I => \N__4111\
        );

    \I__477\ : Span12Mux_s9_h
    port map (
            O => \N__4111\,
            I => \N__4108\
        );

    \I__476\ : Span12Mux_v
    port map (
            O => \N__4108\,
            I => \N__4105\
        );

    \I__475\ : Odrv12
    port map (
            O => \N__4105\,
            I => \SIZ_c_1\
        );

    \I__474\ : InMux
    port map (
            O => \N__4102\,
            I => \N__4099\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__4099\,
            I => \U712_BYTE_ENABLE.N_381\
        );

    \I__472\ : CascadeMux
    port map (
            O => \N__4096\,
            I => \U712_BYTE_ENABLE.N_376_cascade_\
        );

    \I__471\ : IoInMux
    port map (
            O => \N__4093\,
            I => \N__4090\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4090\,
            I => \N__4087\
        );

    \I__469\ : IoSpan4Mux
    port map (
            O => \N__4087\,
            I => \N__4084\
        );

    \I__468\ : Sp12to4
    port map (
            O => \N__4084\,
            I => \N__4081\
        );

    \I__467\ : Span12Mux_s9_h
    port map (
            O => \N__4081\,
            I => \N__4078\
        );

    \I__466\ : Span12Mux_v
    port map (
            O => \N__4078\,
            I => \N__4075\
        );

    \I__465\ : Odrv12
    port map (
            O => \N__4075\,
            I => \N_47_i\
        );

    \I__464\ : CascadeMux
    port map (
            O => \N__4072\,
            I => \N__4069\
        );

    \I__463\ : InMux
    port map (
            O => \N__4069\,
            I => \N__4063\
        );

    \I__462\ : InMux
    port map (
            O => \N__4068\,
            I => \N__4063\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4063\,
            I => \N__4058\
        );

    \I__460\ : InMux
    port map (
            O => \N__4062\,
            I => \N__4055\
        );

    \I__459\ : InMux
    port map (
            O => \N__4061\,
            I => \N__4052\
        );

    \I__458\ : Span4Mux_h
    port map (
            O => \N__4058\,
            I => \N__4045\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4055\,
            I => \N__4045\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__4052\,
            I => \N__4045\
        );

    \I__455\ : Span4Mux_h
    port map (
            O => \N__4045\,
            I => \N__4042\
        );

    \I__454\ : Sp12to4
    port map (
            O => \N__4042\,
            I => \N__4039\
        );

    \I__453\ : Span12Mux_v
    port map (
            O => \N__4039\,
            I => \N__4036\
        );

    \I__452\ : Odrv12
    port map (
            O => \N__4036\,
            I => \A_c_1\
        );

    \I__451\ : InMux
    port map (
            O => \N__4033\,
            I => \N__4030\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4030\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_0\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__4027\,
            I => \N__4022\
        );

    \I__448\ : InMux
    port map (
            O => \N__4026\,
            I => \N__4015\
        );

    \I__447\ : InMux
    port map (
            O => \N__4025\,
            I => \N__4015\
        );

    \I__446\ : InMux
    port map (
            O => \N__4022\,
            I => \N__4015\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4015\,
            I => \U712_BYTE_ENABLE.N_376\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__4012\,
            I => \U712_BYTE_ENABLE.N_377_cascade_\
        );

    \I__443\ : IoInMux
    port map (
            O => \N__4009\,
            I => \N__4006\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4006\,
            I => \N__4003\
        );

    \I__441\ : IoSpan4Mux
    port map (
            O => \N__4003\,
            I => \N__4000\
        );

    \I__440\ : IoSpan4Mux
    port map (
            O => \N__4000\,
            I => \N__3997\
        );

    \I__439\ : Span4Mux_s3_h
    port map (
            O => \N__3997\,
            I => \N__3994\
        );

    \I__438\ : Sp12to4
    port map (
            O => \N__3994\,
            I => \N__3991\
        );

    \I__437\ : Span12Mux_s11_h
    port map (
            O => \N__3991\,
            I => \N__3988\
        );

    \I__436\ : Odrv12
    port map (
            O => \N__3988\,
            I => \N_49_i\
        );

    \I__435\ : InMux
    port map (
            O => \N__3985\,
            I => \N__3982\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3982\,
            I => \N__3979\
        );

    \I__433\ : Span4Mux_v
    port map (
            O => \N__3979\,
            I => \N__3975\
        );

    \I__432\ : InMux
    port map (
            O => \N__3978\,
            I => \N__3972\
        );

    \I__431\ : Sp12to4
    port map (
            O => \N__3975\,
            I => \N__3967\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3972\,
            I => \N__3967\
        );

    \I__429\ : Span12Mux_h
    port map (
            O => \N__3967\,
            I => \N__3964\
        );

    \I__428\ : Span12Mux_v
    port map (
            O => \N__3964\,
            I => \N__3961\
        );

    \I__427\ : Odrv12
    port map (
            O => \N__3961\,
            I => \SIZ_c_0\
        );

    \I__426\ : InMux
    port map (
            O => \N__3958\,
            I => \N__3954\
        );

    \I__425\ : InMux
    port map (
            O => \N__3957\,
            I => \N__3951\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3954\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__3951\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__422\ : InMux
    port map (
            O => \N__3946\,
            I => \N__3942\
        );

    \I__421\ : InMux
    port map (
            O => \N__3945\,
            I => \N__3939\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3942\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3939\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__418\ : InMux
    port map (
            O => \N__3934\,
            I => \N__3930\
        );

    \I__417\ : InMux
    port map (
            O => \N__3933\,
            I => \N__3927\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3930\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3927\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__414\ : InMux
    port map (
            O => \N__3922\,
            I => \N__3918\
        );

    \I__413\ : InMux
    port map (
            O => \N__3921\,
            I => \N__3915\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__3918\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__3915\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__410\ : InMux
    port map (
            O => \N__3910\,
            I => \N__3906\
        );

    \I__409\ : InMux
    port map (
            O => \N__3909\,
            I => \N__3903\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3906\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__3903\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__3898\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_\
        );

    \I__405\ : InMux
    port map (
            O => \N__3895\,
            I => \N__3892\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__3892\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__403\ : InMux
    port map (
            O => \N__3889\,
            I => \N__3879\
        );

    \I__402\ : InMux
    port map (
            O => \N__3888\,
            I => \N__3879\
        );

    \I__401\ : InMux
    port map (
            O => \N__3887\,
            I => \N__3879\
        );

    \I__400\ : InMux
    port map (
            O => \N__3886\,
            I => \N__3876\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3879\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3876\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__397\ : CascadeMux
    port map (
            O => \N__3871\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0_cascade_\
        );

    \I__396\ : InMux
    port map (
            O => \N__3868\,
            I => \N__3862\
        );

    \I__395\ : InMux
    port map (
            O => \N__3867\,
            I => \N__3862\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3862\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__393\ : InMux
    port map (
            O => \N__3859\,
            I => \N__3854\
        );

    \I__392\ : InMux
    port map (
            O => \N__3858\,
            I => \N__3849\
        );

    \I__391\ : InMux
    port map (
            O => \N__3857\,
            I => \N__3849\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3854\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__3849\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__388\ : IoInMux
    port map (
            O => \N__3844\,
            I => \N__3841\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__3841\,
            I => \N__3838\
        );

    \I__386\ : Span12Mux_s0_v
    port map (
            O => \N__3838\,
            I => \N__3835\
        );

    \I__385\ : Span12Mux_v
    port map (
            O => \N__3835\,
            I => \N__3832\
        );

    \I__384\ : Odrv12
    port map (
            O => \N__3832\,
            I => \N_46_i\
        );

    \I__383\ : InMux
    port map (
            O => \N__3829\,
            I => \bfn_8_8_0_\
        );

    \I__382\ : InMux
    port map (
            O => \N__3826\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__381\ : InMux
    port map (
            O => \N__3823\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__380\ : InMux
    port map (
            O => \N__3820\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__379\ : InMux
    port map (
            O => \N__3817\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__378\ : InMux
    port map (
            O => \N__3814\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__377\ : InMux
    port map (
            O => \N__3811\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__376\ : InMux
    port map (
            O => \N__3808\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__375\ : ClkMux
    port map (
            O => \N__3805\,
            I => \N__3802\
        );

    \I__374\ : GlobalMux
    port map (
            O => \N__3802\,
            I => \N__3799\
        );

    \I__373\ : gio2CtrlBuf
    port map (
            O => \N__3799\,
            I => \C1_c_g\
        );

    \I__372\ : InMux
    port map (
            O => \N__3796\,
            I => \N__3792\
        );

    \I__371\ : InMux
    port map (
            O => \N__3795\,
            I => \N__3789\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__3792\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__3789\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__368\ : InMux
    port map (
            O => \N__3784\,
            I => \N__3780\
        );

    \I__367\ : InMux
    port map (
            O => \N__3783\,
            I => \N__3777\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__3780\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__3777\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__364\ : CascadeMux
    port map (
            O => \N__3772\,
            I => \N__3768\
        );

    \I__363\ : InMux
    port map (
            O => \N__3771\,
            I => \N__3765\
        );

    \I__362\ : InMux
    port map (
            O => \N__3768\,
            I => \N__3762\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__3765\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3762\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__359\ : IoInMux
    port map (
            O => \N__3757\,
            I => \N__3754\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3754\,
            I => \N__3751\
        );

    \I__357\ : Span4Mux_s2_v
    port map (
            O => \N__3751\,
            I => \N__3748\
        );

    \I__356\ : Span4Mux_v
    port map (
            O => \N__3748\,
            I => \N__3745\
        );

    \I__355\ : Odrv4
    port map (
            O => \N__3745\,
            I => \CLK80_OUT_i_i\
        );

    \I__354\ : IoInMux
    port map (
            O => \N__3742\,
            I => \N__3739\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__3739\,
            I => \N__3736\
        );

    \I__352\ : Span4Mux_s1_h
    port map (
            O => \N__3736\,
            I => \N__3733\
        );

    \I__351\ : Span4Mux_h
    port map (
            O => \N__3733\,
            I => \N__3730\
        );

    \I__350\ : Sp12to4
    port map (
            O => \N__3730\,
            I => \N__3727\
        );

    \I__349\ : Span12Mux_v
    port map (
            O => \N__3727\,
            I => \N__3724\
        );

    \I__348\ : Odrv12
    port map (
            O => \N__3724\,
            I => \N_882_i\
        );

    \I__347\ : IoInMux
    port map (
            O => \N__3721\,
            I => \N__3718\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__3718\,
            I => \N__3715\
        );

    \I__345\ : Odrv12
    port map (
            O => \N__3715\,
            I => \CLK40_OUT_i_i\
        );

    \I__344\ : InMux
    port map (
            O => \N__3712\,
            I => \N__3709\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3709\,
            I => \N__3706\
        );

    \I__342\ : Span4Mux_h
    port map (
            O => \N__3706\,
            I => \N__3703\
        );

    \I__341\ : Sp12to4
    port map (
            O => \N__3703\,
            I => \N__3700\
        );

    \I__340\ : Span12Mux_v
    port map (
            O => \N__3700\,
            I => \N__3697\
        );

    \I__339\ : Odrv12
    port map (
            O => \N__3697\,
            I => \REGSPACEn_c\
        );

    \I__338\ : InMux
    port map (
            O => \N__3694\,
            I => \N__3688\
        );

    \I__337\ : InMux
    port map (
            O => \N__3693\,
            I => \N__3681\
        );

    \I__336\ : InMux
    port map (
            O => \N__3692\,
            I => \N__3681\
        );

    \I__335\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3681\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__3688\,
            I => \N__3678\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__3681\,
            I => \N__3675\
        );

    \I__332\ : Span4Mux_v
    port map (
            O => \N__3678\,
            I => \N__3672\
        );

    \I__331\ : Span4Mux_v
    port map (
            O => \N__3675\,
            I => \N__3669\
        );

    \I__330\ : Span4Mux_v
    port map (
            O => \N__3672\,
            I => \N__3666\
        );

    \I__329\ : Span4Mux_v
    port map (
            O => \N__3669\,
            I => \N__3663\
        );

    \I__328\ : Sp12to4
    port map (
            O => \N__3666\,
            I => \N__3658\
        );

    \I__327\ : Sp12to4
    port map (
            O => \N__3663\,
            I => \N__3658\
        );

    \I__326\ : Span12Mux_h
    port map (
            O => \N__3658\,
            I => \N__3655\
        );

    \I__325\ : Odrv12
    port map (
            O => \N__3655\,
            I => \CLK40_OUT_i\
        );

    \I__324\ : IoInMux
    port map (
            O => \N__3652\,
            I => \N__3649\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__3649\,
            I => \N__3646\
        );

    \I__322\ : IoSpan4Mux
    port map (
            O => \N__3646\,
            I => \N__3643\
        );

    \I__321\ : Span4Mux_s0_h
    port map (
            O => \N__3643\,
            I => \N__3640\
        );

    \I__320\ : Sp12to4
    port map (
            O => \N__3640\,
            I => \N__3636\
        );

    \I__319\ : CascadeMux
    port map (
            O => \N__3639\,
            I => \N__3633\
        );

    \I__318\ : Span12Mux_v
    port map (
            O => \N__3636\,
            I => \N__3630\
        );

    \I__317\ : InMux
    port map (
            O => \N__3633\,
            I => \N__3627\
        );

    \I__316\ : Odrv12
    port map (
            O => \N__3630\,
            I => \TACK_OUTn\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__3627\,
            I => \TACK_OUTn\
        );

    \I__314\ : IoInMux
    port map (
            O => \N__3622\,
            I => \N__3619\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__3619\,
            I => \N__3616\
        );

    \I__312\ : Span12Mux_s9_v
    port map (
            O => \N__3616\,
            I => \N__3613\
        );

    \I__311\ : Odrv12
    port map (
            O => \N__3613\,
            I => \VBENn_c\
        );

    \I__310\ : IoInMux
    port map (
            O => \N__3610\,
            I => \N__3607\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__3607\,
            I => \N__3604\
        );

    \I__308\ : IoSpan4Mux
    port map (
            O => \N__3604\,
            I => \N__3601\
        );

    \I__307\ : Span4Mux_s2_v
    port map (
            O => \N__3601\,
            I => \N__3598\
        );

    \I__306\ : Sp12to4
    port map (
            O => \N__3598\,
            I => \N__3595\
        );

    \I__305\ : Span12Mux_v
    port map (
            O => \N__3595\,
            I => \N__3592\
        );

    \I__304\ : Odrv12
    port map (
            O => \N__3592\,
            I => \CLK40_IN_c\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7528\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5178\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9229\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4246\,
            lcout => \N_882_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK40C_obuf_RNO_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3694\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_srsts_0_i_o3_0_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4306\,
            in2 => \_gnd_net_\,
            in3 => \N__3712\,
            lcout => \U712_REG_SM.N_295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__3888\,
            in1 => \N__5455\,
            in2 => \N__5416\,
            in3 => \N__3691\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9224\,
            ce => 'H',
            sr => \N__9034\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__3692\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3889\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9224\,
            ce => 'H',
            sr => \N__9034\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111010000"
        )
    port map (
            in0 => \N__3887\,
            in1 => \N__3693\,
            in2 => \N__3639\,
            in3 => \N__3859\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9224\,
            ce => 'H',
            sr => \N__9034\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__5557\,
            in1 => \N__4062\,
            in2 => \N__4142\,
            in3 => \N__8401\,
            lcout => \U712_BYTE_ENABLE.N_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8399\,
            in1 => \N__4061\,
            in2 => \_gnd_net_\,
            in3 => \N__5556\,
            lcout => \U712_BYTE_ENABLE.N_381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_0_a2_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8403\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7651\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3958\,
            in2 => \_gnd_net_\,
            in3 => \N__3829\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__3805\,
            ce => 'H',
            sr => \N__5251\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3784\,
            in2 => \_gnd_net_\,
            in3 => \N__3826\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__3805\,
            ce => 'H',
            sr => \N__5251\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3796\,
            in2 => \_gnd_net_\,
            in3 => \N__3823\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__3805\,
            ce => 'H',
            sr => \N__5251\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3910\,
            in2 => \_gnd_net_\,
            in3 => \N__3820\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__3805\,
            ce => 'H',
            sr => \N__5251\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3771\,
            in2 => \_gnd_net_\,
            in3 => \N__3817\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__3805\,
            ce => 'H',
            sr => \N__5251\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3934\,
            in2 => \_gnd_net_\,
            in3 => \N__3814\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__3805\,
            ce => 'H',
            sr => \N__5251\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3946\,
            in2 => \_gnd_net_\,
            in3 => \N__3811\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__3805\,
            ce => 'H',
            sr => \N__5251\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3922\,
            in2 => \_gnd_net_\,
            in3 => \N__3808\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3805\,
            ce => 'H',
            sr => \N__5251\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__3795\,
            in1 => \N__3783\,
            in2 => \N__3772\,
            in3 => \N__3957\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3945\,
            in2 => \_gnd_net_\,
            in3 => \N__3933\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111111101111"
        )
    port map (
            in0 => \N__3921\,
            in1 => \N__3909\,
            in2 => \N__3898\,
            in3 => \N__3895\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9218\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001001100"
        )
    port map (
            in0 => \N__7968\,
            in1 => \N__7151\,
            in2 => \N__6601\,
            in3 => \N__8023\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3857\,
            in2 => \_gnd_net_\,
            in3 => \N__3867\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__3886\,
            in1 => \N__5453\,
            in2 => \N__3871\,
            in3 => \N__5433\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9221\,
            ce => 'H',
            sr => \N__9030\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3868\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9221\,
            ce => 'H',
            sr => \N__9030\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3858\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9221\,
            ce => 'H',
            sr => \N__9030\
        );

    \U712_BYTE_ENABLE.N_46_i_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__4317\,
            in1 => \N__4183\,
            in2 => \N__4027\,
            in3 => \N__7800\,
            lcout => \N_46_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__4143\,
            in1 => \N__4068\,
            in2 => \N__5567\,
            in3 => \N__8397\,
            lcout => \U712_BYTE_ENABLE.N_383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_0_0_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7698\,
            in2 => \_gnd_net_\,
            in3 => \N__8091\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_0\,
            ltout => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_48_i_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100011"
        )
    port map (
            in0 => \N__7801\,
            in1 => \N__4177\,
            in2 => \N__4171\,
            in3 => \N__4025\,
            lcout => \N_48_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__8398\,
            in1 => \N__4144\,
            in2 => \_gnd_net_\,
            in3 => \N__3985\,
            lcout => \U712_BYTE_ENABLE.N_376\,
            ltout => \U712_BYTE_ENABLE.N_376_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_47_i_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__4102\,
            in1 => \N__4318\,
            in2 => \N__4096\,
            in3 => \N__7766\,
            lcout => \N_47_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_0_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5561\,
            in2 => \N__4072\,
            in3 => \N__8400\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_377_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_49_i_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__4033\,
            in1 => \N__4026\,
            in2 => \N__4012\,
            in3 => \N__7767\,
            lcout => \N_49_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDS_OUT_2_0_a2_0_a2_0_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3978\,
            in2 => \_gnd_net_\,
            in3 => \N__6039\,
            lcout => \U712_REG_SM.LDS_OUT_2_0_a2_0_a2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4945\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9196\,
            ce => \N__8593\,
            sr => \N__9047\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5031\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9196\,
            ce => \N__8593\,
            sr => \N__9047\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5074\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9202\,
            ce => \N__8592\,
            sr => \N__9042\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4987\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9202\,
            ce => \N__8592\,
            sr => \N__9042\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__7591\,
            in1 => \N__6859\,
            in2 => \N__4327\,
            in3 => \N__6811\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__8402\,
            in1 => \N__8013\,
            in2 => \_gnd_net_\,
            in3 => \N__6600\,
            lcout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0_0_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7702\,
            in2 => \_gnd_net_\,
            in3 => \N__8084\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__4564\,
            in1 => \N__6892\,
            in2 => \N__8027\,
            in3 => \N__6721\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9213\,
            ce => 'H',
            sr => \N__9031\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010001"
        )
    port map (
            in0 => \N__4305\,
            in1 => \N__4273\,
            in2 => \N__8404\,
            in3 => \N__4582\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9213\,
            ce => 'H',
            sr => \N__9031\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__7590\,
            in1 => \N__5454\,
            in2 => \_gnd_net_\,
            in3 => \N__5411\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9219\,
            ce => \N__5389\,
            sr => \N__9021\
        );

    \U712_REG_SM.REGENn_1_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111110100010"
        )
    port map (
            in0 => \N__4196\,
            in1 => \N__4873\,
            in2 => \N__4822\,
            in3 => \N__4681\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9222\,
            ce => 'H',
            sr => \N__9015\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__4377\,
            in1 => \N__4680\,
            in2 => \N__4365\,
            in3 => \N__4820\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9222\,
            ce => 'H',
            sr => \N__9015\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__5621\,
            in1 => \N__4378\,
            in2 => \N__4366\,
            in3 => \N__5598\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9222\,
            ce => 'H',
            sr => \N__9015\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__5599\,
            in1 => \N__4911\,
            in2 => \N__4711\,
            in3 => \N__5622\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9222\,
            ce => 'H',
            sr => \N__9015\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__4816\,
            in1 => \N__4840\,
            in2 => \N__4864\,
            in3 => \N__4333\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9222\,
            ce => 'H',
            sr => \N__9015\
        );

    \U712_REG_SM.C3_SYNC_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4348\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9222\,
            ce => 'H',
            sr => \N__9015\
        );

    \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__4890\,
            in1 => \N__4600\,
            in2 => \N__4636\,
            in3 => \N__4735\,
            lcout => \U712_REG_SM.N_292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5701\,
            in2 => \_gnd_net_\,
            in3 => \N__4785\,
            lcout => \U712_REG_SM.N_338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__4531\,
            in1 => \N__5655\,
            in2 => \N__5683\,
            in3 => \N__4518\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9225\,
            ce => 'H',
            sr => \N__9002\
        );

    \U712_REG_SM.REG_CYCLE_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111010"
        )
    port map (
            in0 => \N__4517\,
            in1 => \N__5702\,
            in2 => \N__7642\,
            in3 => \N__4529\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9225\,
            ce => 'H',
            sr => \N__9002\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010101000"
        )
    port map (
            in0 => \N__4530\,
            in1 => \N__4519\,
            in2 => \N__4915\,
            in3 => \N__4710\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9225\,
            ce => 'H',
            sr => \N__9002\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__5654\,
            in1 => \N__5682\,
            in2 => \N__4789\,
            in3 => \N__5703\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9225\,
            ce => 'H',
            sr => \N__9002\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__4507\,
            in1 => \N__8396\,
            in2 => \N__4495\,
            in3 => \N__4471\,
            lcout => \U712_CHIP_RAM.N_310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__4477\,
            in1 => \N__8371\,
            in2 => \N__8868\,
            in3 => \N__4951\,
            lcout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__8372\,
            in1 => \N__4993\,
            in2 => \N__4465\,
            in3 => \N__8848\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__4456\,
            in1 => \N__4441\,
            in2 => \N__4429\,
            in3 => \N__8373\,
            lcout => \U712_CHIP_RAM.N_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111100010"
        )
    port map (
            in0 => \N__4549\,
            in1 => \N__5226\,
            in2 => \N__8512\,
            in3 => \N__4426\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9197\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__6088\,
            in1 => \N__8390\,
            in2 => \N__8869\,
            in3 => \N__4957\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8391\,
            in1 => \N__4420\,
            in2 => \N__4402\,
            in3 => \N__4399\,
            lcout => \U712_CHIP_RAM.N_309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000101000011"
        )
    port map (
            in0 => \N__6599\,
            in1 => \N__6858\,
            in2 => \N__7977\,
            in3 => \N__7155\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_e_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000101"
        )
    port map (
            in0 => \N__5225\,
            in1 => \N__6390\,
            in2 => \N__4552\,
            in3 => \N__7294\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9197\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_3_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__4548\,
            in1 => \N__6574\,
            in2 => \N__6391\,
            in3 => \N__6673\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9203\,
            ce => \N__4645\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQDMA1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__7941\,
            in1 => \N__7156\,
            in2 => \_gnd_net_\,
            in3 => \N__7089\,
            lcout => \U712_CHIP_RAM.N_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_1_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7904\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6573\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c2\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__6651\,
            in1 => \N__7024\,
            in2 => \N__4537\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7903\,
            in1 => \N__6572\,
            in2 => \_gnd_net_\,
            in3 => \N__6650\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6652\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7905\,
            lcout => \U712_CHIP_RAM.N_427\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__7027\,
            in1 => \N__6797\,
            in2 => \N__6661\,
            in3 => \N__6741\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_tz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIN8RQ7_3_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__7589\,
            in1 => \N__4558\,
            in2 => \N__4534\,
            in3 => \N__6962\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIBUNAE_0_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__6382\,
            in1 => \N__6502\,
            in2 => \N__4651\,
            in3 => \N__7949\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_sbtinv_3_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4648\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__4626\,
            in1 => \N__4595\,
            in2 => \_gnd_net_\,
            in3 => \N__4580\,
            lcout => \U712_CHIP_RAM.N_278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4596\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM_DBR_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9210\,
            ce => 'H',
            sr => \N__9022\
        );

    \U712_CHIP_RAM.DBR_SYNC_0_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4615\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM_DBR_SYNC_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9210\,
            ce => 'H',
            sr => \N__9022\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100110000"
        )
    port map (
            in0 => \N__6040\,
            in1 => \N__5208\,
            in2 => \N__8174\,
            in3 => \N__4581\,
            lcout => \U712_CHIP_RAM.N_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIRB433_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6653\,
            in1 => \N__5281\,
            in2 => \N__6742\,
            in3 => \N__8160\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__5324\,
            in1 => \N__5346\,
            in2 => \N__9094\,
            in3 => \N__4669\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4667\,
            in1 => \N__5345\,
            in2 => \_gnd_net_\,
            in3 => \N__5323\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_15_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__9089\,
            in1 => \_gnd_net_\,
            in2 => \N__4690\,
            in3 => \N__5379\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__5380\,
            in1 => \N__4687\,
            in2 => \N__5365\,
            in3 => \N__9090\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4838\,
            in2 => \_gnd_net_\,
            in3 => \N__4859\,
            lcout => \U712_REG_SM.N_492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__4668\,
            in1 => \N__9085\,
            in2 => \_gnd_net_\,
            in3 => \N__5325\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNICU4F1_2_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__5754\,
            in1 => \N__5146\,
            in2 => \N__5800\,
            in3 => \N__4772\,
            lcout => \U712_REG_SM.N_491\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI90BP_0_2_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5753\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5796\,
            lcout => \U712_REG_SM.N_273\,
            ltout => \U712_REG_SM.N_273_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_1_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4821\,
            in1 => \N__5147\,
            in2 => \N__4654\,
            in3 => \N__4773\,
            lcout => \U712_REG_SM.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4886\,
            in2 => \_gnd_net_\,
            in3 => \N__4734\,
            lcout => \U712_REG_SM.N_279\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5795\,
            in2 => \_gnd_net_\,
            in3 => \N__5752\,
            lcout => \U712_REG_SM.N_282\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4907\,
            in2 => \_gnd_net_\,
            in3 => \N__4706\,
            lcout => \U712_REG_SM.N_355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNINB3L1_1_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__5620\,
            in1 => \N__4774\,
            in2 => \N__4891\,
            in3 => \N__5148\,
            lcout => \U712_REG_SM.N_420\,
            ltout => \U712_REG_SM.N_420_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_2_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001010000"
        )
    port map (
            in0 => \N__4815\,
            in1 => \N__4860\,
            in2 => \N__4843\,
            in3 => \N__4839\,
            lcout => \U712_REG_SM.DS_EN_RNOZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_2_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4770\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9223\,
            ce => 'H',
            sr => \N__9003\
        );

    \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5773\,
            in2 => \_gnd_net_\,
            in3 => \N__4743\,
            lcout => \U712_REG_SM.N_281\,
            ltout => \U712_REG_SM.N_281_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_0_1_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4771\,
            in1 => \N__5144\,
            in2 => \N__4792\,
            in3 => \N__4722\,
            lcout => \U712_REG_SM.N_300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_1_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5145\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9223\,
            ce => 'H',
            sr => \N__9003\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__5774\,
            in1 => \N__4769\,
            in2 => \N__4747\,
            in3 => \N__5143\,
            lcout => \U712_REG_SM.N_274\,
            ltout => \U712_REG_SM.N_274_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__4723\,
            in1 => \_gnd_net_\,
            in2 => \N__4714\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.N_297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_0_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5182\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9223\,
            ce => 'H',
            sr => \N__9003\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__6025\,
            in1 => \N__5781\,
            in2 => \_gnd_net_\,
            in3 => \N__5149\,
            lcout => \U712_REG_SM.N_210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__5119\,
            in1 => \N__7331\,
            in2 => \_gnd_net_\,
            in3 => \N__8510\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9185\,
            ce => \N__7216\,
            sr => \N__9043\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__5101\,
            in1 => \N__7332\,
            in2 => \_gnd_net_\,
            in3 => \N__8511\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9185\,
            ce => \N__7216\,
            sr => \N__9043\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5073\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9189\,
            ce => \N__8551\,
            sr => \N__9036\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5032\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9189\,
            ce => \N__8551\,
            sr => \N__9036\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4983\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9189\,
            ce => \N__8551\,
            sr => \N__9036\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6112\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9189\,
            ce => \N__8551\,
            sr => \N__9036\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4941\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9189\,
            ce => \N__8551\,
            sr => \N__9036\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6454\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9189\,
            ce => \N__8551\,
            sr => \N__9036\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010011"
        )
    port map (
            in0 => \N__5257\,
            in1 => \N__6397\,
            in2 => \N__8862\,
            in3 => \N__8353\,
            lcout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNITDMK_3_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8758\,
            in1 => \N__7277\,
            in2 => \N__8486\,
            in3 => \N__8835\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => \U712_CHIP_RAM.REFRESH_RST_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNI9T531_3_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__8836\,
            in1 => \N__8759\,
            in2 => \N__5239\,
            in3 => \N__7278\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__8837\,
            in1 => \N__6403\,
            in2 => \N__8395\,
            in3 => \N__5236\,
            lcout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111001010"
        )
    port map (
            in0 => \N__6361\,
            in1 => \N__8841\,
            in2 => \N__5230\,
            in3 => \N__6349\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBDIR_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011000111110000"
        )
    port map (
            in0 => \N__6717\,
            in1 => \N__5209\,
            in2 => \N__5981\,
            in3 => \N__6884\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9198\,
            ce => 'H',
            sr => \N__9023\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI3EN62_0_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__8171\,
            in1 => \N__6933\,
            in2 => \_gnd_net_\,
            in3 => \N__5282\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI3EN62_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__5283\,
            in1 => \_gnd_net_\,
            in2 => \N__6953\,
            in3 => \N__8172\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_340_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIQU7BE_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111010"
        )
    port map (
            in0 => \N__6489\,
            in1 => \_gnd_net_\,
            in2 => \N__5287\,
            in3 => \N__6716\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_START_RNIQU7BEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__5284\,
            in1 => \_gnd_net_\,
            in2 => \N__6954\,
            in3 => \N__8173\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a2_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011011"
        )
    port map (
            in0 => \N__6707\,
            in1 => \N__5266\,
            in2 => \N__7945\,
            in3 => \N__6490\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7000\,
            in2 => \_gnd_net_\,
            in3 => \N__6647\,
            lcout => \U712_CHIP_RAM.N_263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7588\,
            in2 => \_gnd_net_\,
            in3 => \N__6805\,
            lcout => \U712_CHIP_RAM.N_336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6311\,
            in1 => \N__6327\,
            in2 => \_gnd_net_\,
            in3 => \N__6649\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOO5O1_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6648\,
            in1 => \N__6575\,
            in2 => \N__7020\,
            in3 => \N__7137\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_417_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIN7BL3_1_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__7072\,
            in1 => \N__6843\,
            in2 => \N__5260\,
            in3 => \N__6571\,
            lcout => \U712_CHIP_RAM.N_265\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7899\,
            in1 => \N__6576\,
            in2 => \_gnd_net_\,
            in3 => \N__6312\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6570\,
            in2 => \_gnd_net_\,
            in3 => \N__7898\,
            lcout => \U712_CHIP_RAM.N_270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__5482\,
            in1 => \N__5470\,
            in2 => \N__6343\,
            in3 => \N__6804\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9211\,
            ce => \N__5299\,
            sr => \N__9010\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5637\,
            in2 => \_gnd_net_\,
            in3 => \N__5461\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__7575\,
            in1 => \N__5434\,
            in2 => \N__5419\,
            in3 => \N__5415\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_298_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5392\,
            in3 => \N__9084\,
            lcout => \U712_CYCLE_TERM.N_298_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5378\,
            in1 => \N__5361\,
            in2 => \N__5350\,
            in3 => \N__5326\,
            lcout => \U712_CHIP_RAM.N_267\,
            ltout => \U712_CHIP_RAM.N_267_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__7025\,
            in1 => \N__6465\,
            in2 => \N__5305\,
            in3 => \N__6963\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__9083\,
            in1 => \_gnd_net_\,
            in2 => \N__5302\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_204_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_1_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__6577\,
            in1 => \N__7908\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_276_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_2_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5755\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9215\,
            ce => 'H',
            sr => \N__9004\
        );

    \U712_REG_SM.C3_SYNC_1_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5782\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9215\,
            ce => 'H',
            sr => \N__9004\
        );

    \U712_REG_SM.DS_EN_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__6077\,
            in1 => \N__5734\,
            in2 => \N__5728\,
            in3 => \N__5716\,
            lcout => \U712_REG_SM.DS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9215\,
            ce => 'H',
            sr => \N__9004\
        );

    \U712_REG_SM.REG_TACK_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101010000"
        )
    port map (
            in0 => \N__5710\,
            in1 => \N__5678\,
            in2 => \N__5641\,
            in3 => \N__5662\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9215\,
            ce => 'H',
            sr => \N__9004\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__8047\,
            in1 => \N__7726\,
            in2 => \N__8180\,
            in3 => \N__7682\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9215\,
            ce => 'H',
            sr => \N__9004\
        );

    \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5626\,
            in2 => \_gnd_net_\,
            in3 => \N__5597\,
            lcout => \U712_REG_SM.N_302\,
            ltout => \U712_REG_SM.N_302_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDS_OUT_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001101"
        )
    port map (
            in0 => \N__5580\,
            in1 => \N__5568\,
            in2 => \N__5584\,
            in3 => \N__5511\,
            lcout => \U712_REG_SM.LDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9220\,
            ce => 'H',
            sr => \N__8997\
        );

    \U712_REG_SM.UDS_OUT_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100000111"
        )
    port map (
            in0 => \N__5581\,
            in1 => \N__5569\,
            in2 => \N__5521\,
            in3 => \N__6063\,
            lcout => \U712_REG_SM.UDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9220\,
            ce => 'H',
            sr => \N__8997\
        );

    \U712_REG_SM.LDS_OUT_RNIL31J_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5512\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6078\,
            lcout => \U712_REG_SM_un1_LDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_RNIUP9B_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6079\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6064\,
            lcout => \U712_REG_SM_un1_UDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_i_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001010"
        )
    port map (
            in0 => \N__7696\,
            in1 => \N__6035\,
            in2 => \N__5988\,
            in3 => \N__7643\,
            lcout => \N_208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__5929\,
            in1 => \N__8380\,
            in2 => \N__8901\,
            in3 => \N__8692\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8382\,
            in1 => \N__5917\,
            in2 => \N__5899\,
            in3 => \N__5896\,
            lcout => \U712_CHIP_RAM.N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__6412\,
            in1 => \N__8381\,
            in2 => \N__8902\,
            in3 => \N__5875\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8383\,
            in1 => \N__5866\,
            in2 => \N__5848\,
            in3 => \N__5845\,
            lcout => \U712_CHIP_RAM.N_311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__7326\,
            in1 => \N__6175\,
            in2 => \_gnd_net_\,
            in3 => \N__8522\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9182\,
            ce => \N__7225\,
            sr => \N__9033\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000101"
        )
    port map (
            in0 => \N__8896\,
            in1 => \N__6298\,
            in2 => \N__8528\,
            in3 => \N__7328\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9182\,
            ce => \N__7225\,
            sr => \N__9033\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7325\,
            in1 => \N__8521\,
            in2 => \N__8905\,
            in3 => \N__8773\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9182\,
            ce => \N__7225\,
            sr => \N__9033\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000101"
        )
    port map (
            in0 => \N__8897\,
            in1 => \N__6262\,
            in2 => \N__8529\,
            in3 => \N__7329\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9182\,
            ce => \N__7225\,
            sr => \N__9033\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__8514\,
            in1 => \_gnd_net_\,
            in2 => \N__6121\,
            in3 => \N__7327\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9182\,
            ce => \N__7225\,
            sr => \N__9033\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001010101"
        )
    port map (
            in0 => \N__6220\,
            in1 => \N__6214\,
            in2 => \N__6199\,
            in3 => \N__8385\,
            lcout => \U712_CHIP_RAM.N_312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIV62J1_3_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9092\,
            in2 => \_gnd_net_\,
            in3 => \N__6169\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__7321\,
            in1 => \N__8852\,
            in2 => \_gnd_net_\,
            in3 => \N__8513\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__6163\,
            in1 => \N__8384\,
            in2 => \N__6148\,
            in3 => \N__6127\,
            lcout => \U712_CHIP_RAM.N_306\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6108\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9188\,
            ce => \N__8581\,
            sr => \N__9020\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6453\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9188\,
            ce => \N__8581\,
            sr => \N__9020\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8679\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9188\,
            ce => \N__8581\,
            sr => \N__9020\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8722\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9188\,
            ce => \N__8581\,
            sr => \N__9020\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111100"
        )
    port map (
            in0 => \N__7145\,
            in1 => \N__6383\,
            in2 => \N__7964\,
            in3 => \N__6851\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__6961\,
            in1 => \N__7085\,
            in2 => \_gnd_net_\,
            in3 => \N__6587\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110001"
        )
    port map (
            in0 => \N__7146\,
            in1 => \N__7940\,
            in2 => \N__6352\,
            in3 => \N__6589\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6849\,
            in1 => \N__6807\,
            in2 => \N__7965\,
            in3 => \N__8028\,
            lcout => \U712_CHIP_RAM.N_369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__6331\,
            in1 => \N__6660\,
            in2 => \N__6316\,
            in3 => \N__7019\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9191\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6588\,
            in1 => \N__7018\,
            in2 => \_gnd_net_\,
            in3 => \N__6659\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGURED_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_3_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101001011010"
        )
    port map (
            in0 => \N__6850\,
            in1 => \N__6586\,
            in2 => \N__7966\,
            in3 => \N__7144\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111110"
        )
    port map (
            in0 => \N__6952\,
            in1 => \N__6582\,
            in2 => \N__7963\,
            in3 => \N__6658\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_3_0_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__6790\,
            in1 => \_gnd_net_\,
            in2 => \N__6664\,
            in3 => \N__7011\,
            lcout => \U712_CHIP_RAM.N_148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__7042\,
            in1 => \N__7129\,
            in2 => \_gnd_net_\,
            in3 => \N__7171\,
            lcout => \U712_CHIP_RAM.N_275\,
            ltout => \U712_CHIP_RAM.N_275_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_3_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__7010\,
            in1 => \N__6657\,
            in2 => \N__6604\,
            in3 => \N__6581\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_423_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJ42D8_0_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101010"
        )
    port map (
            in0 => \N__9082\,
            in1 => \N__6478\,
            in2 => \N__6505\,
            in3 => \N__6501\,
            lcout => \U712_CHIP_RAM.N_303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6789\,
            in2 => \_gnd_net_\,
            in3 => \N__7906\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_0_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__7907\,
            in1 => \N__6472\,
            in2 => \N__6806\,
            in3 => \N__7130\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9195\,
            ce => 'H',
            sr => \N__9006\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6796\,
            in1 => \N__6845\,
            in2 => \N__7090\,
            in3 => \N__6466\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011111010"
        )
    port map (
            in0 => \N__7170\,
            in1 => \_gnd_net_\,
            in2 => \N__7174\,
            in3 => \N__6701\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9201\,
            ce => 'H',
            sr => \N__8998\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__7041\,
            in1 => \N__7169\,
            in2 => \_gnd_net_\,
            in3 => \N__7147\,
            lcout => \U712_CHIP_RAM.N_428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7054\,
            in1 => \N__7683\,
            in2 => \_gnd_net_\,
            in3 => \N__8284\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9201\,
            ce => 'H',
            sr => \N__8998\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_3_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__6795\,
            in1 => \N__7026\,
            in2 => \N__6964\,
            in3 => \N__6904\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_375_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_3_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__6888\,
            in1 => \_gnd_net_\,
            in2 => \N__6865\,
            in3 => \N__6700\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9081\,
            in1 => \_gnd_net_\,
            in2 => \N__6862\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__6844\,
            in1 => \N__6794\,
            in2 => \_gnd_net_\,
            in3 => \N__6740\,
            lcout => \U712_CHIP_RAM.N_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7967\,
            in2 => \_gnd_net_\,
            in3 => \N__8170\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9206\,
            ce => \N__6682\,
            sr => \N__8996\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7569\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RASn_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7333\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9183\,
            ce => 'H',
            sr => \N__9048\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__8602\,
            in1 => \N__8386\,
            in2 => \N__8903\,
            in3 => \N__8641\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_i_m3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__7498\,
            in1 => \N__8387\,
            in2 => \N__7480\,
            in3 => \N__7477\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_313_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__7330\,
            in1 => \_gnd_net_\,
            in2 => \N__7459\,
            in3 => \N__8527\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9186\,
            ce => \N__7217\,
            sr => \N__9044\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__7435\,
            in1 => \N__7392\,
            in2 => \N__8635\,
            in3 => \N__8388\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9190\,
            ce => \N__7203\,
            sr => \N__9037\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__9280\,
            in1 => \N__7393\,
            in2 => \N__7384\,
            in3 => \N__8389\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9190\,
            ce => \N__7203\,
            sr => \N__9037\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__7342\,
            in1 => \N__7320\,
            in2 => \_gnd_net_\,
            in3 => \N__8523\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9193\,
            ce => \N__7218\,
            sr => \N__9032\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__9091\,
            in1 => \N__8043\,
            in2 => \_gnd_net_\,
            in3 => \N__7725\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__8182\,
            in1 => \N__8283\,
            in2 => \N__7976\,
            in3 => \N__8109\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9205\,
            ce => 'H',
            sr => \N__9016\
        );

    \U712_CHIP_RAM.BANK0_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__8218\,
            in1 => \N__8193\,
            in2 => \N__7975\,
            in3 => \N__8108\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9205\,
            ce => 'H',
            sr => \N__9016\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8181\,
            in2 => \_gnd_net_\,
            in3 => \N__7956\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.DMA_CYCLE_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101111111001100"
        )
    port map (
            in0 => \N__8125\,
            in1 => \N__8065\,
            in2 => \N__8113\,
            in3 => \N__8110\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9205\,
            ce => 'H',
            sr => \N__9016\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7721\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9212\,
            ce => 'H',
            sr => \N__9011\
        );

    \U712_CHIP_RAM.CLK_EN_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111100100011"
        )
    port map (
            in0 => \N__8029\,
            in1 => \N__7984\,
            in2 => \N__7978\,
            in3 => \N__7812\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9212\,
            ce => 'H',
            sr => \N__9011\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7799\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7768\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9216\,
            ce => 'H',
            sr => \N__9005\
        );

    \U712_BUFFERS.un1_DRDENn_0_a2_0_a2_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7697\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7650\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_14_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8904\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9184\,
            ce => 'H',
            sr => \N__9050\
        );

    \U712_CHIP_RAM.CRCSn_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8772\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9187\,
            ce => 'H',
            sr => \N__9049\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8718\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9194\,
            ce => \N__8547\,
            sr => \N__9045\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8680\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9194\,
            ce => \N__8547\,
            sr => \N__9045\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8626\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9194\,
            ce => \N__8547\,
            sr => \N__9045\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8625\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9199\,
            ce => \N__8585\,
            sr => \N__9038\
        );

    \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__9093\,
            in1 => \N__9235\,
            in2 => \_gnd_net_\,
            in3 => \N__9246\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8530\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9200\,
            ce => 'H',
            sr => \N__9051\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8416\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9276\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9217\,
            ce => 'H',
            sr => \N__9046\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9247\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9217\,
            ce => 'H',
            sr => \N__9046\
        );
end \INTERFACE\;

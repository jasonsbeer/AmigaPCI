// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 6 2025 19:31:10

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    TT,
    TM,
    A,
    D,
    RESETn,
    OVL,
    CONFIGENn,
    PIO_S0,
    PORTSIZE,
    TICK60,
    CIACS0n,
    CPUCONFn,
    CLK6,
    CLK_CIA,
    BUFENn,
    AUTOBOOT,
    RnW,
    PIO_P2,
    CIACS1n,
    BRIDGE_ENn,
    PIO_S1,
    ATA_MODE_S,
    PIO_P0,
    TICK50,
    TCIn,
    TBIn,
    RAMSPACEn,
    CLK40_IN,
    CLK28_IN,
    REGSPACEn,
    TSn,
    RTC_ENn,
    PIO_S2,
    ATA_ENn,
    TACKn,
    ATA_MODE_P,
    ROMENn,
    PIO_P1);

    input [1:0] TT;
    input [1:0] TM;
    input [31:1] A;
    inout [7:4] D;
    input RESETn;
    input OVL;
    output CONFIGENn;
    output PIO_S0;
    output PORTSIZE;
    output TICK60;
    output CIACS0n;
    input CPUCONFn;
    input CLK6;
    output CLK_CIA;
    output BUFENn;
    input AUTOBOOT;
    input RnW;
    output PIO_P2;
    output CIACS1n;
    output BRIDGE_ENn;
    output PIO_S1;
    input ATA_MODE_S;
    output PIO_P0;
    output TICK50;
    output TCIn;
    output TBIn;
    output RAMSPACEn;
    input CLK40_IN;
    input CLK28_IN;
    output REGSPACEn;
    input TSn;
    output RTC_ENn;
    output PIO_S2;
    output ATA_ENn;
    inout TACKn;
    input ATA_MODE_P;
    output ROMENn;
    output PIO_P1;

    wire N__12507;
    wire N__12506;
    wire N__12505;
    wire N__12497;
    wire N__12496;
    wire N__12495;
    wire N__12487;
    wire N__12486;
    wire N__12485;
    wire N__12476;
    wire N__12475;
    wire N__12474;
    wire N__12467;
    wire N__12466;
    wire N__12465;
    wire N__12458;
    wire N__12457;
    wire N__12456;
    wire N__12449;
    wire N__12448;
    wire N__12447;
    wire N__12440;
    wire N__12439;
    wire N__12438;
    wire N__12431;
    wire N__12430;
    wire N__12429;
    wire N__12422;
    wire N__12421;
    wire N__12420;
    wire N__12413;
    wire N__12412;
    wire N__12411;
    wire N__12404;
    wire N__12403;
    wire N__12402;
    wire N__12395;
    wire N__12394;
    wire N__12393;
    wire N__12386;
    wire N__12385;
    wire N__12384;
    wire N__12377;
    wire N__12376;
    wire N__12375;
    wire N__12368;
    wire N__12367;
    wire N__12366;
    wire N__12359;
    wire N__12358;
    wire N__12357;
    wire N__12350;
    wire N__12349;
    wire N__12348;
    wire N__12341;
    wire N__12340;
    wire N__12339;
    wire N__12332;
    wire N__12331;
    wire N__12330;
    wire N__12323;
    wire N__12322;
    wire N__12321;
    wire N__12314;
    wire N__12313;
    wire N__12312;
    wire N__12305;
    wire N__12304;
    wire N__12303;
    wire N__12296;
    wire N__12295;
    wire N__12294;
    wire N__12287;
    wire N__12286;
    wire N__12285;
    wire N__12278;
    wire N__12277;
    wire N__12276;
    wire N__12269;
    wire N__12268;
    wire N__12267;
    wire N__12260;
    wire N__12259;
    wire N__12258;
    wire N__12251;
    wire N__12250;
    wire N__12249;
    wire N__12242;
    wire N__12241;
    wire N__12240;
    wire N__12233;
    wire N__12232;
    wire N__12231;
    wire N__12224;
    wire N__12223;
    wire N__12222;
    wire N__12215;
    wire N__12214;
    wire N__12213;
    wire N__12206;
    wire N__12205;
    wire N__12204;
    wire N__12197;
    wire N__12196;
    wire N__12195;
    wire N__12188;
    wire N__12187;
    wire N__12186;
    wire N__12179;
    wire N__12178;
    wire N__12177;
    wire N__12170;
    wire N__12169;
    wire N__12168;
    wire N__12161;
    wire N__12160;
    wire N__12159;
    wire N__12152;
    wire N__12151;
    wire N__12150;
    wire N__12143;
    wire N__12142;
    wire N__12141;
    wire N__12134;
    wire N__12133;
    wire N__12132;
    wire N__12125;
    wire N__12124;
    wire N__12123;
    wire N__12116;
    wire N__12115;
    wire N__12114;
    wire N__12107;
    wire N__12106;
    wire N__12105;
    wire N__12098;
    wire N__12097;
    wire N__12096;
    wire N__12089;
    wire N__12088;
    wire N__12087;
    wire N__12080;
    wire N__12079;
    wire N__12078;
    wire N__12071;
    wire N__12070;
    wire N__12069;
    wire N__12062;
    wire N__12061;
    wire N__12060;
    wire N__12053;
    wire N__12052;
    wire N__12051;
    wire N__12044;
    wire N__12043;
    wire N__12042;
    wire N__12035;
    wire N__12034;
    wire N__12033;
    wire N__12026;
    wire N__12025;
    wire N__12024;
    wire N__12017;
    wire N__12016;
    wire N__12015;
    wire N__12008;
    wire N__12007;
    wire N__12006;
    wire N__11999;
    wire N__11998;
    wire N__11997;
    wire N__11990;
    wire N__11989;
    wire N__11988;
    wire N__11981;
    wire N__11980;
    wire N__11979;
    wire N__11972;
    wire N__11971;
    wire N__11970;
    wire N__11963;
    wire N__11962;
    wire N__11961;
    wire N__11954;
    wire N__11953;
    wire N__11952;
    wire N__11945;
    wire N__11944;
    wire N__11943;
    wire N__11936;
    wire N__11935;
    wire N__11934;
    wire N__11927;
    wire N__11926;
    wire N__11925;
    wire N__11918;
    wire N__11917;
    wire N__11916;
    wire N__11909;
    wire N__11908;
    wire N__11907;
    wire N__11890;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11878;
    wire N__11875;
    wire N__11872;
    wire N__11869;
    wire N__11866;
    wire N__11865;
    wire N__11862;
    wire N__11859;
    wire N__11854;
    wire N__11853;
    wire N__11852;
    wire N__11851;
    wire N__11850;
    wire N__11849;
    wire N__11848;
    wire N__11847;
    wire N__11846;
    wire N__11827;
    wire N__11824;
    wire N__11821;
    wire N__11820;
    wire N__11817;
    wire N__11814;
    wire N__11809;
    wire N__11806;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11794;
    wire N__11791;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11779;
    wire N__11776;
    wire N__11773;
    wire N__11770;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11758;
    wire N__11755;
    wire N__11752;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11740;
    wire N__11737;
    wire N__11734;
    wire N__11731;
    wire N__11730;
    wire N__11727;
    wire N__11724;
    wire N__11719;
    wire N__11716;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11704;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11683;
    wire N__11680;
    wire N__11677;
    wire N__11674;
    wire N__11673;
    wire N__11670;
    wire N__11667;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11638;
    wire N__11637;
    wire N__11634;
    wire N__11633;
    wire N__11628;
    wire N__11625;
    wire N__11620;
    wire N__11619;
    wire N__11618;
    wire N__11617;
    wire N__11614;
    wire N__11611;
    wire N__11606;
    wire N__11603;
    wire N__11596;
    wire N__11595;
    wire N__11592;
    wire N__11589;
    wire N__11584;
    wire N__11581;
    wire N__11580;
    wire N__11577;
    wire N__11574;
    wire N__11569;
    wire N__11566;
    wire N__11565;
    wire N__11562;
    wire N__11559;
    wire N__11554;
    wire N__11551;
    wire N__11548;
    wire N__11547;
    wire N__11544;
    wire N__11541;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11520;
    wire N__11517;
    wire N__11514;
    wire N__11509;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11487;
    wire N__11484;
    wire N__11481;
    wire N__11476;
    wire N__11473;
    wire N__11472;
    wire N__11469;
    wire N__11466;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11424;
    wire N__11421;
    wire N__11418;
    wire N__11413;
    wire N__11410;
    wire N__11409;
    wire N__11406;
    wire N__11403;
    wire N__11398;
    wire N__11395;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11383;
    wire N__11380;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11368;
    wire N__11365;
    wire N__11362;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11335;
    wire N__11332;
    wire N__11329;
    wire N__11328;
    wire N__11325;
    wire N__11324;
    wire N__11323;
    wire N__11322;
    wire N__11321;
    wire N__11320;
    wire N__11319;
    wire N__11316;
    wire N__11307;
    wire N__11300;
    wire N__11293;
    wire N__11292;
    wire N__11291;
    wire N__11290;
    wire N__11289;
    wire N__11288;
    wire N__11287;
    wire N__11286;
    wire N__11283;
    wire N__11274;
    wire N__11267;
    wire N__11260;
    wire N__11259;
    wire N__11258;
    wire N__11257;
    wire N__11254;
    wire N__11253;
    wire N__11250;
    wire N__11249;
    wire N__11248;
    wire N__11247;
    wire N__11244;
    wire N__11241;
    wire N__11236;
    wire N__11233;
    wire N__11224;
    wire N__11215;
    wire N__11214;
    wire N__11211;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11194;
    wire N__11193;
    wire N__11192;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11180;
    wire N__11177;
    wire N__11170;
    wire N__11167;
    wire N__11166;
    wire N__11163;
    wire N__11160;
    wire N__11155;
    wire N__11152;
    wire N__11151;
    wire N__11148;
    wire N__11145;
    wire N__11140;
    wire N__11137;
    wire N__11136;
    wire N__11133;
    wire N__11130;
    wire N__11125;
    wire N__11122;
    wire N__11119;
    wire N__11116;
    wire N__11113;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11101;
    wire N__11098;
    wire N__11097;
    wire N__11094;
    wire N__11091;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11077;
    wire N__11076;
    wire N__11075;
    wire N__11074;
    wire N__11073;
    wire N__11070;
    wire N__11069;
    wire N__11068;
    wire N__11059;
    wire N__11052;
    wire N__11047;
    wire N__11046;
    wire N__11045;
    wire N__11044;
    wire N__11043;
    wire N__11042;
    wire N__11041;
    wire N__11038;
    wire N__11035;
    wire N__11032;
    wire N__11025;
    wire N__11018;
    wire N__11011;
    wire N__11008;
    wire N__11005;
    wire N__11002;
    wire N__10999;
    wire N__10998;
    wire N__10997;
    wire N__10996;
    wire N__10995;
    wire N__10994;
    wire N__10993;
    wire N__10992;
    wire N__10989;
    wire N__10982;
    wire N__10973;
    wire N__10966;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10956;
    wire N__10953;
    wire N__10950;
    wire N__10945;
    wire N__10944;
    wire N__10943;
    wire N__10942;
    wire N__10937;
    wire N__10932;
    wire N__10927;
    wire N__10926;
    wire N__10925;
    wire N__10924;
    wire N__10919;
    wire N__10914;
    wire N__10909;
    wire N__10908;
    wire N__10907;
    wire N__10904;
    wire N__10903;
    wire N__10900;
    wire N__10895;
    wire N__10890;
    wire N__10885;
    wire N__10884;
    wire N__10883;
    wire N__10882;
    wire N__10881;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10866;
    wire N__10861;
    wire N__10852;
    wire N__10851;
    wire N__10848;
    wire N__10845;
    wire N__10840;
    wire N__10837;
    wire N__10836;
    wire N__10835;
    wire N__10834;
    wire N__10833;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10825;
    wire N__10824;
    wire N__10823;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10809;
    wire N__10808;
    wire N__10803;
    wire N__10796;
    wire N__10793;
    wire N__10788;
    wire N__10783;
    wire N__10780;
    wire N__10777;
    wire N__10776;
    wire N__10773;
    wire N__10768;
    wire N__10767;
    wire N__10764;
    wire N__10759;
    wire N__10756;
    wire N__10753;
    wire N__10752;
    wire N__10751;
    wire N__10746;
    wire N__10745;
    wire N__10742;
    wire N__10741;
    wire N__10740;
    wire N__10739;
    wire N__10730;
    wire N__10725;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10714;
    wire N__10711;
    wire N__10708;
    wire N__10705;
    wire N__10702;
    wire N__10699;
    wire N__10696;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10686;
    wire N__10683;
    wire N__10676;
    wire N__10669;
    wire N__10666;
    wire N__10663;
    wire N__10656;
    wire N__10649;
    wire N__10642;
    wire N__10639;
    wire N__10636;
    wire N__10633;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10615;
    wire N__10612;
    wire N__10609;
    wire N__10608;
    wire N__10605;
    wire N__10602;
    wire N__10597;
    wire N__10594;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10579;
    wire N__10578;
    wire N__10577;
    wire N__10574;
    wire N__10571;
    wire N__10568;
    wire N__10561;
    wire N__10560;
    wire N__10557;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10540;
    wire N__10537;
    wire N__10536;
    wire N__10535;
    wire N__10534;
    wire N__10533;
    wire N__10532;
    wire N__10529;
    wire N__10524;
    wire N__10519;
    wire N__10516;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10498;
    wire N__10497;
    wire N__10492;
    wire N__10489;
    wire N__10486;
    wire N__10483;
    wire N__10480;
    wire N__10479;
    wire N__10478;
    wire N__10477;
    wire N__10468;
    wire N__10465;
    wire N__10462;
    wire N__10461;
    wire N__10460;
    wire N__10459;
    wire N__10456;
    wire N__10451;
    wire N__10448;
    wire N__10441;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10431;
    wire N__10428;
    wire N__10425;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10417;
    wire N__10414;
    wire N__10409;
    wire N__10404;
    wire N__10399;
    wire N__10396;
    wire N__10393;
    wire N__10392;
    wire N__10391;
    wire N__10390;
    wire N__10389;
    wire N__10388;
    wire N__10387;
    wire N__10384;
    wire N__10381;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10363;
    wire N__10360;
    wire N__10359;
    wire N__10358;
    wire N__10357;
    wire N__10356;
    wire N__10353;
    wire N__10352;
    wire N__10351;
    wire N__10350;
    wire N__10349;
    wire N__10348;
    wire N__10345;
    wire N__10342;
    wire N__10339;
    wire N__10336;
    wire N__10303;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10288;
    wire N__10285;
    wire N__10284;
    wire N__10283;
    wire N__10280;
    wire N__10275;
    wire N__10270;
    wire N__10269;
    wire N__10268;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10256;
    wire N__10249;
    wire N__10248;
    wire N__10245;
    wire N__10242;
    wire N__10237;
    wire N__10234;
    wire N__10231;
    wire N__10230;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10210;
    wire N__10207;
    wire N__10204;
    wire N__10203;
    wire N__10202;
    wire N__10201;
    wire N__10198;
    wire N__10195;
    wire N__10192;
    wire N__10191;
    wire N__10188;
    wire N__10185;
    wire N__10180;
    wire N__10175;
    wire N__10168;
    wire N__10165;
    wire N__10162;
    wire N__10159;
    wire N__10156;
    wire N__10155;
    wire N__10152;
    wire N__10149;
    wire N__10146;
    wire N__10143;
    wire N__10138;
    wire N__10135;
    wire N__10134;
    wire N__10133;
    wire N__10132;
    wire N__10131;
    wire N__10126;
    wire N__10123;
    wire N__10118;
    wire N__10111;
    wire N__10110;
    wire N__10107;
    wire N__10106;
    wire N__10105;
    wire N__10104;
    wire N__10101;
    wire N__10098;
    wire N__10093;
    wire N__10090;
    wire N__10081;
    wire N__10080;
    wire N__10077;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10059;
    wire N__10056;
    wire N__10053;
    wire N__10048;
    wire N__10045;
    wire N__10042;
    wire N__10039;
    wire N__10036;
    wire N__10035;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10015;
    wire N__10014;
    wire N__10011;
    wire N__10008;
    wire N__10005;
    wire N__10002;
    wire N__9999;
    wire N__9988;
    wire N__9985;
    wire N__9982;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9970;
    wire N__9969;
    wire N__9966;
    wire N__9963;
    wire N__9962;
    wire N__9957;
    wire N__9954;
    wire N__9949;
    wire N__9948;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9930;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9919;
    wire N__9916;
    wire N__9911;
    wire N__9908;
    wire N__9901;
    wire N__9898;
    wire N__9897;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9879;
    wire N__9874;
    wire N__9873;
    wire N__9870;
    wire N__9867;
    wire N__9862;
    wire N__9859;
    wire N__9856;
    wire N__9855;
    wire N__9852;
    wire N__9849;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9799;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9787;
    wire N__9786;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9776;
    wire N__9773;
    wire N__9768;
    wire N__9763;
    wire N__9760;
    wire N__9759;
    wire N__9756;
    wire N__9753;
    wire N__9750;
    wire N__9747;
    wire N__9742;
    wire N__9739;
    wire N__9736;
    wire N__9735;
    wire N__9734;
    wire N__9733;
    wire N__9732;
    wire N__9731;
    wire N__9730;
    wire N__9729;
    wire N__9728;
    wire N__9727;
    wire N__9726;
    wire N__9703;
    wire N__9700;
    wire N__9697;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9687;
    wire N__9684;
    wire N__9681;
    wire N__9676;
    wire N__9675;
    wire N__9674;
    wire N__9673;
    wire N__9670;
    wire N__9665;
    wire N__9662;
    wire N__9655;
    wire N__9654;
    wire N__9653;
    wire N__9652;
    wire N__9649;
    wire N__9646;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9628;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9616;
    wire N__9613;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9601;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9591;
    wire N__9588;
    wire N__9583;
    wire N__9580;
    wire N__9577;
    wire N__9576;
    wire N__9575;
    wire N__9572;
    wire N__9567;
    wire N__9562;
    wire N__9561;
    wire N__9558;
    wire N__9555;
    wire N__9550;
    wire N__9549;
    wire N__9548;
    wire N__9545;
    wire N__9540;
    wire N__9535;
    wire N__9532;
    wire N__9529;
    wire N__9528;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9511;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9499;
    wire N__9498;
    wire N__9497;
    wire N__9494;
    wire N__9493;
    wire N__9492;
    wire N__9489;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9475;
    wire N__9472;
    wire N__9469;
    wire N__9466;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9450;
    wire N__9447;
    wire N__9440;
    wire N__9437;
    wire N__9432;
    wire N__9427;
    wire N__9424;
    wire N__9421;
    wire N__9418;
    wire N__9417;
    wire N__9416;
    wire N__9415;
    wire N__9414;
    wire N__9413;
    wire N__9412;
    wire N__9401;
    wire N__9396;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9355;
    wire N__9354;
    wire N__9351;
    wire N__9348;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9324;
    wire N__9319;
    wire N__9316;
    wire N__9315;
    wire N__9312;
    wire N__9309;
    wire N__9304;
    wire N__9303;
    wire N__9298;
    wire N__9297;
    wire N__9296;
    wire N__9295;
    wire N__9292;
    wire N__9291;
    wire N__9286;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9276;
    wire N__9271;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9202;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9136;
    wire N__9133;
    wire N__9130;
    wire N__9127;
    wire N__9126;
    wire N__9125;
    wire N__9124;
    wire N__9121;
    wire N__9116;
    wire N__9111;
    wire N__9106;
    wire N__9105;
    wire N__9100;
    wire N__9097;
    wire N__9094;
    wire N__9093;
    wire N__9092;
    wire N__9091;
    wire N__9090;
    wire N__9079;
    wire N__9076;
    wire N__9075;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9064;
    wire N__9055;
    wire N__9052;
    wire N__9051;
    wire N__9050;
    wire N__9047;
    wire N__9046;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9028;
    wire N__9025;
    wire N__9024;
    wire N__9023;
    wire N__9022;
    wire N__9019;
    wire N__9016;
    wire N__9011;
    wire N__9004;
    wire N__9003;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8988;
    wire N__8987;
    wire N__8982;
    wire N__8979;
    wire N__8974;
    wire N__8971;
    wire N__8968;
    wire N__8965;
    wire N__8964;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8941;
    wire N__8940;
    wire N__8937;
    wire N__8934;
    wire N__8929;
    wire N__8926;
    wire N__8925;
    wire N__8922;
    wire N__8919;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8881;
    wire N__8878;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8866;
    wire N__8863;
    wire N__8860;
    wire N__8859;
    wire N__8856;
    wire N__8853;
    wire N__8850;
    wire N__8845;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8806;
    wire N__8803;
    wire N__8802;
    wire N__8799;
    wire N__8796;
    wire N__8795;
    wire N__8790;
    wire N__8789;
    wire N__8788;
    wire N__8787;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8770;
    wire N__8761;
    wire N__8758;
    wire N__8755;
    wire N__8754;
    wire N__8753;
    wire N__8752;
    wire N__8751;
    wire N__8750;
    wire N__8749;
    wire N__8746;
    wire N__8743;
    wire N__8740;
    wire N__8737;
    wire N__8730;
    wire N__8719;
    wire N__8716;
    wire N__8713;
    wire N__8710;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8698;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8683;
    wire N__8680;
    wire N__8677;
    wire N__8676;
    wire N__8671;
    wire N__8668;
    wire N__8667;
    wire N__8664;
    wire N__8663;
    wire N__8662;
    wire N__8661;
    wire N__8658;
    wire N__8657;
    wire N__8656;
    wire N__8653;
    wire N__8650;
    wire N__8641;
    wire N__8638;
    wire N__8629;
    wire N__8628;
    wire N__8627;
    wire N__8626;
    wire N__8625;
    wire N__8624;
    wire N__8623;
    wire N__8620;
    wire N__8617;
    wire N__8614;
    wire N__8611;
    wire N__8602;
    wire N__8599;
    wire N__8590;
    wire N__8589;
    wire N__8588;
    wire N__8585;
    wire N__8580;
    wire N__8575;
    wire N__8572;
    wire N__8571;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8547;
    wire N__8546;
    wire N__8545;
    wire N__8544;
    wire N__8543;
    wire N__8542;
    wire N__8539;
    wire N__8538;
    wire N__8537;
    wire N__8536;
    wire N__8533;
    wire N__8532;
    wire N__8531;
    wire N__8528;
    wire N__8523;
    wire N__8522;
    wire N__8517;
    wire N__8514;
    wire N__8509;
    wire N__8506;
    wire N__8505;
    wire N__8502;
    wire N__8497;
    wire N__8492;
    wire N__8489;
    wire N__8488;
    wire N__8485;
    wire N__8478;
    wire N__8475;
    wire N__8466;
    wire N__8463;
    wire N__8460;
    wire N__8455;
    wire N__8450;
    wire N__8445;
    wire N__8442;
    wire N__8437;
    wire N__8434;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8421;
    wire N__8420;
    wire N__8419;
    wire N__8418;
    wire N__8413;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8399;
    wire N__8394;
    wire N__8389;
    wire N__8388;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8341;
    wire N__8338;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8321;
    wire N__8316;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8304;
    wire N__8301;
    wire N__8298;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8253;
    wire N__8252;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8241;
    wire N__8238;
    wire N__8237;
    wire N__8236;
    wire N__8233;
    wire N__8230;
    wire N__8227;
    wire N__8224;
    wire N__8223;
    wire N__8222;
    wire N__8221;
    wire N__8218;
    wire N__8217;
    wire N__8216;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8202;
    wire N__8199;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8183;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8167;
    wire N__8164;
    wire N__8159;
    wire N__8156;
    wire N__8153;
    wire N__8150;
    wire N__8145;
    wire N__8138;
    wire N__8131;
    wire N__8128;
    wire N__8127;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8119;
    wire N__8116;
    wire N__8113;
    wire N__8110;
    wire N__8107;
    wire N__8098;
    wire N__8097;
    wire N__8096;
    wire N__8093;
    wire N__8092;
    wire N__8089;
    wire N__8086;
    wire N__8083;
    wire N__8080;
    wire N__8077;
    wire N__8068;
    wire N__8065;
    wire N__8062;
    wire N__8059;
    wire N__8056;
    wire N__8055;
    wire N__8052;
    wire N__8049;
    wire N__8044;
    wire N__8041;
    wire N__8040;
    wire N__8037;
    wire N__8034;
    wire N__8033;
    wire N__8032;
    wire N__8031;
    wire N__8030;
    wire N__8029;
    wire N__8028;
    wire N__8025;
    wire N__8022;
    wire N__8019;
    wire N__8018;
    wire N__8017;
    wire N__8014;
    wire N__8011;
    wire N__8010;
    wire N__8005;
    wire N__8004;
    wire N__8001;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7983;
    wire N__7980;
    wire N__7977;
    wire N__7974;
    wire N__7973;
    wire N__7970;
    wire N__7969;
    wire N__7964;
    wire N__7961;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7933;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7914;
    wire N__7909;
    wire N__7906;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7885;
    wire N__7882;
    wire N__7879;
    wire N__7878;
    wire N__7877;
    wire N__7876;
    wire N__7871;
    wire N__7870;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7851;
    wire N__7848;
    wire N__7845;
    wire N__7842;
    wire N__7839;
    wire N__7838;
    wire N__7835;
    wire N__7830;
    wire N__7825;
    wire N__7824;
    wire N__7823;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7813;
    wire N__7810;
    wire N__7805;
    wire N__7802;
    wire N__7789;
    wire N__7786;
    wire N__7783;
    wire N__7780;
    wire N__7779;
    wire N__7778;
    wire N__7777;
    wire N__7774;
    wire N__7771;
    wire N__7770;
    wire N__7767;
    wire N__7764;
    wire N__7761;
    wire N__7758;
    wire N__7755;
    wire N__7750;
    wire N__7747;
    wire N__7742;
    wire N__7739;
    wire N__7736;
    wire N__7735;
    wire N__7734;
    wire N__7731;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7710;
    wire N__7707;
    wire N__7702;
    wire N__7699;
    wire N__7696;
    wire N__7693;
    wire N__7690;
    wire N__7687;
    wire N__7684;
    wire N__7681;
    wire N__7678;
    wire N__7675;
    wire N__7672;
    wire N__7669;
    wire N__7666;
    wire N__7665;
    wire N__7662;
    wire N__7661;
    wire N__7660;
    wire N__7659;
    wire N__7658;
    wire N__7655;
    wire N__7654;
    wire N__7651;
    wire N__7648;
    wire N__7645;
    wire N__7640;
    wire N__7635;
    wire N__7630;
    wire N__7625;
    wire N__7622;
    wire N__7621;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7596;
    wire N__7595;
    wire N__7592;
    wire N__7589;
    wire N__7588;
    wire N__7585;
    wire N__7582;
    wire N__7577;
    wire N__7570;
    wire N__7569;
    wire N__7566;
    wire N__7563;
    wire N__7558;
    wire N__7557;
    wire N__7556;
    wire N__7553;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7541;
    wire N__7540;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7525;
    wire N__7522;
    wire N__7517;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7492;
    wire N__7491;
    wire N__7490;
    wire N__7489;
    wire N__7488;
    wire N__7487;
    wire N__7486;
    wire N__7483;
    wire N__7482;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7462;
    wire N__7461;
    wire N__7458;
    wire N__7455;
    wire N__7452;
    wire N__7451;
    wire N__7450;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7428;
    wire N__7421;
    wire N__7418;
    wire N__7415;
    wire N__7414;
    wire N__7411;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7390;
    wire N__7387;
    wire N__7382;
    wire N__7379;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7358;
    wire N__7353;
    wire N__7348;
    wire N__7345;
    wire N__7344;
    wire N__7343;
    wire N__7342;
    wire N__7339;
    wire N__7336;
    wire N__7331;
    wire N__7324;
    wire N__7323;
    wire N__7322;
    wire N__7319;
    wire N__7318;
    wire N__7315;
    wire N__7312;
    wire N__7309;
    wire N__7306;
    wire N__7297;
    wire N__7296;
    wire N__7295;
    wire N__7294;
    wire N__7293;
    wire N__7292;
    wire N__7279;
    wire N__7278;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7267;
    wire N__7266;
    wire N__7265;
    wire N__7264;
    wire N__7261;
    wire N__7258;
    wire N__7247;
    wire N__7240;
    wire N__7237;
    wire N__7236;
    wire N__7235;
    wire N__7234;
    wire N__7231;
    wire N__7224;
    wire N__7219;
    wire N__7218;
    wire N__7217;
    wire N__7214;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7200;
    wire N__7195;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7185;
    wire N__7184;
    wire N__7181;
    wire N__7178;
    wire N__7175;
    wire N__7172;
    wire N__7165;
    wire N__7162;
    wire N__7159;
    wire N__7156;
    wire N__7153;
    wire N__7150;
    wire N__7147;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7125;
    wire N__7122;
    wire N__7117;
    wire N__7114;
    wire N__7111;
    wire N__7110;
    wire N__7109;
    wire N__7106;
    wire N__7103;
    wire N__7100;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7086;
    wire N__7085;
    wire N__7076;
    wire N__7073;
    wire N__7070;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7047;
    wire N__7042;
    wire N__7041;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7030;
    wire N__7029;
    wire N__7026;
    wire N__7023;
    wire N__7020;
    wire N__7017;
    wire N__7014;
    wire N__7013;
    wire N__7010;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6990;
    wire N__6987;
    wire N__6984;
    wire N__6981;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6967;
    wire N__6966;
    wire N__6961;
    wire N__6958;
    wire N__6955;
    wire N__6952;
    wire N__6949;
    wire N__6946;
    wire N__6945;
    wire N__6944;
    wire N__6941;
    wire N__6936;
    wire N__6931;
    wire N__6930;
    wire N__6927;
    wire N__6926;
    wire N__6923;
    wire N__6920;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6900;
    wire N__6895;
    wire N__6892;
    wire N__6891;
    wire N__6888;
    wire N__6885;
    wire N__6880;
    wire N__6877;
    wire N__6874;
    wire N__6873;
    wire N__6870;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6850;
    wire N__6847;
    wire N__6846;
    wire N__6843;
    wire N__6840;
    wire N__6837;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6815;
    wire N__6808;
    wire N__6805;
    wire N__6804;
    wire N__6803;
    wire N__6802;
    wire N__6797;
    wire N__6792;
    wire N__6787;
    wire N__6786;
    wire N__6783;
    wire N__6782;
    wire N__6779;
    wire N__6778;
    wire N__6777;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6765;
    wire N__6760;
    wire N__6757;
    wire N__6748;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6730;
    wire N__6727;
    wire N__6724;
    wire N__6721;
    wire N__6718;
    wire N__6717;
    wire N__6716;
    wire N__6715;
    wire N__6714;
    wire N__6711;
    wire N__6710;
    wire N__6707;
    wire N__6704;
    wire N__6699;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6687;
    wire N__6684;
    wire N__6681;
    wire N__6670;
    wire N__6669;
    wire N__6666;
    wire N__6663;
    wire N__6660;
    wire N__6659;
    wire N__6658;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6621;
    wire N__6620;
    wire N__6619;
    wire N__6616;
    wire N__6611;
    wire N__6608;
    wire N__6607;
    wire N__6604;
    wire N__6599;
    wire N__6596;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6564;
    wire N__6561;
    wire N__6558;
    wire N__6555;
    wire N__6552;
    wire N__6549;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6529;
    wire N__6528;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6507;
    wire N__6504;
    wire N__6499;
    wire N__6496;
    wire N__6493;
    wire N__6490;
    wire N__6487;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6465;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6402;
    wire N__6401;
    wire N__6400;
    wire N__6397;
    wire N__6396;
    wire N__6391;
    wire N__6388;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6376;
    wire N__6373;
    wire N__6372;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6336;
    wire N__6333;
    wire N__6328;
    wire N__6325;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6300;
    wire N__6299;
    wire N__6298;
    wire N__6297;
    wire N__6296;
    wire N__6295;
    wire N__6294;
    wire N__6289;
    wire N__6288;
    wire N__6285;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6271;
    wire N__6270;
    wire N__6267;
    wire N__6262;
    wire N__6257;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6247;
    wire N__6246;
    wire N__6245;
    wire N__6244;
    wire N__6243;
    wire N__6234;
    wire N__6233;
    wire N__6228;
    wire N__6221;
    wire N__6216;
    wire N__6213;
    wire N__6210;
    wire N__6203;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6186;
    wire N__6183;
    wire N__6178;
    wire N__6177;
    wire N__6176;
    wire N__6171;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6160;
    wire N__6159;
    wire N__6158;
    wire N__6155;
    wire N__6154;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6121;
    wire N__6120;
    wire N__6115;
    wire N__6112;
    wire N__6109;
    wire N__6108;
    wire N__6105;
    wire N__6102;
    wire N__6099;
    wire N__6096;
    wire N__6091;
    wire N__6088;
    wire N__6087;
    wire N__6082;
    wire N__6081;
    wire N__6078;
    wire N__6075;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6065;
    wire N__6062;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6050;
    wire N__6047;
    wire N__6040;
    wire N__6037;
    wire N__6036;
    wire N__6033;
    wire N__6032;
    wire N__6027;
    wire N__6026;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6008;
    wire N__6005;
    wire N__6000;
    wire N__5995;
    wire N__5992;
    wire N__5991;
    wire N__5988;
    wire N__5987;
    wire N__5984;
    wire N__5979;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5957;
    wire N__5952;
    wire N__5947;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5924;
    wire N__5923;
    wire N__5922;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5899;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5887;
    wire N__5884;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5872;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5848;
    wire N__5845;
    wire N__5844;
    wire N__5841;
    wire N__5838;
    wire N__5833;
    wire N__5830;
    wire N__5829;
    wire N__5826;
    wire N__5823;
    wire N__5818;
    wire N__5817;
    wire N__5816;
    wire N__5815;
    wire N__5814;
    wire N__5811;
    wire N__5810;
    wire N__5803;
    wire N__5802;
    wire N__5799;
    wire N__5796;
    wire N__5793;
    wire N__5790;
    wire N__5789;
    wire N__5788;
    wire N__5785;
    wire N__5782;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5751;
    wire N__5746;
    wire N__5745;
    wire N__5742;
    wire N__5737;
    wire N__5734;
    wire N__5733;
    wire N__5730;
    wire N__5729;
    wire N__5728;
    wire N__5727;
    wire N__5724;
    wire N__5721;
    wire N__5716;
    wire N__5713;
    wire N__5712;
    wire N__5709;
    wire N__5704;
    wire N__5703;
    wire N__5702;
    wire N__5701;
    wire N__5698;
    wire N__5697;
    wire N__5696;
    wire N__5695;
    wire N__5694;
    wire N__5693;
    wire N__5690;
    wire N__5685;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5667;
    wire N__5664;
    wire N__5659;
    wire N__5644;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5614;
    wire N__5611;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5598;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5581;
    wire N__5580;
    wire N__5579;
    wire N__5578;
    wire N__5577;
    wire N__5576;
    wire N__5575;
    wire N__5570;
    wire N__5565;
    wire N__5564;
    wire N__5561;
    wire N__5560;
    wire N__5559;
    wire N__5556;
    wire N__5555;
    wire N__5552;
    wire N__5547;
    wire N__5544;
    wire N__5543;
    wire N__5542;
    wire N__5541;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5526;
    wire N__5523;
    wire N__5518;
    wire N__5513;
    wire N__5508;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5488;
    wire N__5485;
    wire N__5478;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5466;
    wire N__5465;
    wire N__5464;
    wire N__5459;
    wire N__5456;
    wire N__5455;
    wire N__5452;
    wire N__5451;
    wire N__5450;
    wire N__5449;
    wire N__5448;
    wire N__5445;
    wire N__5442;
    wire N__5437;
    wire N__5434;
    wire N__5433;
    wire N__5432;
    wire N__5431;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5414;
    wire N__5409;
    wire N__5406;
    wire N__5403;
    wire N__5400;
    wire N__5387;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5340;
    wire N__5339;
    wire N__5338;
    wire N__5335;
    wire N__5334;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5315;
    wire N__5312;
    wire N__5307;
    wire N__5304;
    wire N__5301;
    wire N__5298;
    wire N__5293;
    wire N__5292;
    wire N__5291;
    wire N__5288;
    wire N__5283;
    wire N__5280;
    wire N__5279;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5259;
    wire N__5256;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5242;
    wire N__5241;
    wire N__5240;
    wire N__5239;
    wire N__5236;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5202;
    wire N__5199;
    wire N__5194;
    wire N__5191;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5152;
    wire N__5151;
    wire N__5148;
    wire N__5145;
    wire N__5140;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5104;
    wire N__5103;
    wire N__5102;
    wire N__5101;
    wire N__5092;
    wire N__5089;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5071;
    wire N__5070;
    wire N__5065;
    wire N__5062;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5035;
    wire N__5032;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5020;
    wire N__5017;
    wire N__5014;
    wire N__5011;
    wire N__5008;
    wire N__5005;
    wire N__5002;
    wire N__4999;
    wire N__4998;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4981;
    wire N__4978;
    wire N__4975;
    wire N__4974;
    wire N__4973;
    wire N__4968;
    wire N__4967;
    wire N__4966;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4939;
    wire N__4936;
    wire N__4933;
    wire N__4930;
    wire N__4927;
    wire N__4924;
    wire N__4921;
    wire N__4918;
    wire N__4915;
    wire N__4912;
    wire N__4909;
    wire N__4906;
    wire N__4903;
    wire N__4900;
    wire N__4897;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4882;
    wire N__4879;
    wire N__4876;
    wire N__4873;
    wire N__4870;
    wire N__4867;
    wire N__4864;
    wire N__4861;
    wire N__4858;
    wire N__4857;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4846;
    wire N__4839;
    wire N__4836;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4822;
    wire N__4819;
    wire N__4816;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4804;
    wire N__4801;
    wire N__4798;
    wire N__4797;
    wire N__4796;
    wire N__4791;
    wire N__4788;
    wire N__4783;
    wire N__4780;
    wire N__4777;
    wire N__4774;
    wire N__4771;
    wire N__4770;
    wire N__4767;
    wire N__4764;
    wire N__4759;
    wire N__4756;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4744;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4729;
    wire N__4728;
    wire N__4725;
    wire N__4722;
    wire N__4717;
    wire N__4714;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4695;
    wire N__4692;
    wire N__4689;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4672;
    wire N__4669;
    wire N__4666;
    wire N__4663;
    wire N__4660;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4648;
    wire N__4645;
    wire N__4644;
    wire N__4639;
    wire N__4636;
    wire N__4633;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4615;
    wire N__4612;
    wire N__4609;
    wire N__4606;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4584;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4576;
    wire N__4573;
    wire N__4572;
    wire N__4571;
    wire N__4568;
    wire N__4559;
    wire N__4556;
    wire N__4549;
    wire N__4546;
    wire N__4545;
    wire N__4544;
    wire N__4543;
    wire N__4534;
    wire N__4533;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4515;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4479;
    wire N__4476;
    wire N__4473;
    wire N__4470;
    wire N__4465;
    wire N__4462;
    wire N__4459;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4447;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4420;
    wire N__4419;
    wire N__4418;
    wire N__4417;
    wire N__4416;
    wire N__4415;
    wire N__4414;
    wire N__4413;
    wire N__4412;
    wire N__4411;
    wire N__4410;
    wire N__4409;
    wire N__4384;
    wire CLK80_OUT;
    wire PIO_S0_c;
    wire GNDG0;
    wire PIO_P0_c;
    wire VCCG0;
    wire \U409_AUTOCONFIG.N_67_cascade_ ;
    wire \U409_AUTOCONFIG.N_214_1 ;
    wire A_c_6;
    wire A_c_7;
    wire \U409_AUTOCONFIG.un1_A_18Z0Z_0_cascade_ ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_cascade_ ;
    wire \U409_AUTOCONFIG.N_63 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_1_2_0_cascade_ ;
    wire \U409_AUTOCONFIG.N_196_1_cascade_ ;
    wire \U409_AUTOCONFIG.LIDE_OUT_7_0_62_i_i_a3_0 ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5_cascade_ ;
    wire \INVU409_AUTOCONFIG.LIDE_CONFC_net ;
    wire \U409_AUTOCONFIG.ATA_BASE10Z0Z_2 ;
    wire \U409_AUTOCONFIG.ATA_BASE10_cascade_ ;
    wire U409_AUTOCONFIG_D_OUT_0_i_3;
    wire \U409_ADDRESS_DECODE.g0_i_a4_0Z0Z_2_cascade_ ;
    wire \INVU409_AUTOCONFIG.STATE_0C_net ;
    wire \U409_AUTOCONFIG.N_55_cascade_ ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ;
    wire CPUCONFn_c;
    wire \U409_AUTOCONFIG.N_40 ;
    wire \U409_AUTOCONFIG.N_59_1_cascade_ ;
    wire \U409_AUTOCONFIG.N_61 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_2_cascade_ ;
    wire \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ;
    wire \U409_AUTOCONFIG.N_67 ;
    wire \U409_AUTOCONFIG.N_56 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_1_0 ;
    wire \U409_AUTOCONFIG.N_59_1 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_8_sqmuxa ;
    wire \U409_AUTOCONFIG.N_57 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_1 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_8_sqmuxa_cascade_ ;
    wire \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ;
    wire \U409_AUTOCONFIG.LIDE_OUT_7_94_i_i_1_tz_cascade_ ;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7_cascade_ ;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_4 ;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_10 ;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9_cascade_ ;
    wire TT_c_1;
    wire TT_c_0;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8 ;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3 ;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4_cascade_ ;
    wire AUTOCONFIG_SPACE_cascade_;
    wire D_1_i;
    wire \INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ;
    wire U409_AUTOCONFIG_D_OUT_0_i_0;
    wire \U409_TRANSFER_ACK.G_14_0_a7_1_3_cascade_ ;
    wire \U409_AUTOCONFIG.un1_AZ0Z_18 ;
    wire \U409_AUTOCONFIG.STATEZ0Z_0 ;
    wire \U409_ADDRESS_DECODE.g0_i_a4_1Z0Z_3 ;
    wire \U409_ADDRESS_DECODE.g0_i_a4Z0Z_1 ;
    wire \U409_AUTOCONFIG.AC_STARTZ0 ;
    wire \U409_AUTOCONFIG.LIDE_OUTc_0_0 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ1Z_0 ;
    wire \U409_AUTOCONFIG.N_50 ;
    wire \U409_AUTOCONFIG.LIDE_OUTc_0_0_0 ;
    wire \U409_AUTOCONFIG.N_48 ;
    wire \U409_AUTOCONFIG.AC_START_RNI777KZ0Z2 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ;
    wire \INVU409_AUTOCONFIG.LIDE_OUT_0C_net ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_1 ;
    wire U409_AUTOCONFIG_D_OUT_0_i_1;
    wire \U409_AUTOCONFIG.BRIDGE_CONFZ0 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ;
    wire U409_AUTOCONFIG_D_OUT_0_i_2;
    wire BRIDGE_BASE_1;
    wire BRIDGE_BASE_2;
    wire A_c_5;
    wire \U409_AUTOCONFIG.N_68 ;
    wire A_c_4;
    wire \U409_AUTOCONFIG.N_47 ;
    wire AUTOBOOT_c;
    wire \U409_AUTOCONFIG.N_196_1 ;
    wire A_c_2;
    wire A_c_3;
    wire \U409_AUTOCONFIG.N_54 ;
    wire \U409_ADDRESS_DECODE.g2_5_0 ;
    wire \U409_ADDRESS_DECODE.g2_6_0_cascade_ ;
    wire A_c_29;
    wire A_c_30;
    wire A_c_27;
    wire A_c_26;
    wire A_c_25;
    wire A_c_24;
    wire \U409_ADDRESS_DECODE.g2Z0Z_4 ;
    wire \U409_ADDRESS_DECODE.un1_Z2_SPACE_7Z0Z_1_cascade_ ;
    wire \U409_ADDRESS_DECODE.un1_Z2_SPACE_6Z0Z_1 ;
    wire \U409_ADDRESS_DECODE.un1_Z2_SPACE_6Z0Z_0 ;
    wire \U409_ADDRESS_DECODE.un1_Z2_SPACE_7Z0Z_3_cascade_ ;
    wire RnW_c;
    wire \U409_ADDRESS_DECODE.un1_Z2_SPACEZ0_cascade_ ;
    wire \U409_ADDRESS_DECODE.g2Z0Z_10 ;
    wire \U409_ADDRESS_DECODE.g2Z0Z_11_cascade_ ;
    wire \U409_ADDRESS_DECODE.g2Z0Z_9 ;
    wire A_c_1;
    wire \U409_AUTOCONFIG.LIDE_CONFZ0 ;
    wire \U409_AUTOCONFIG.un1_STATE_1_0 ;
    wire BRIDGE_BASE_0;
    wire \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_2_cascade_ ;
    wire CONFIGENn_c;
    wire ATA_BASE_5;
    wire \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_0 ;
    wire \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_4 ;
    wire A_c_31;
    wire U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0_cascade_ ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ;
    wire \U409_ADDRESS_DECODE.g2Z0Z_5 ;
    wire A_c_28;
    wire U409_ADDRESS_DECODE_g2_6;
    wire U409_ADDRESS_DECODE_g2_7_cascade_;
    wire \U409_TRANSFER_ACK.G_14_0_o7_0 ;
    wire U409_ADDRESS_DECODE_un1_RTC_ENn_i;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3 ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3_cascade_ ;
    wire ATA_BASE_2;
    wire \INVU409_AUTOCONFIG.ATA_BASE_2C_net ;
    wire D_in_4;
    wire D_in_5;
    wire D_in_6;
    wire \U409_AUTOCONFIG.LIDE_CONF_RNIHQ9AZ0Z3 ;
    wire \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ;
    wire BRIDGE_BASE_3;
    wire un1_AUTOCONFIG_SPACE;
    wire \U409_AUTOCONFIG.STATE_RNI0FVT2Z0Z_0 ;
    wire D_in_7;
    wire ATA_BASE_3;
    wire \INVU409_AUTOCONFIG.ATA_BASE_7C_net ;
    wire U409_ADDRESS_DECODE_ATA_ROM_d;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net ;
    wire \U409_ADDRESS_DECODE.g0_i_0Z0Z_0 ;
    wire \U409_ADDRESS_DECODE.g0_i_o4Z0Z_1 ;
    wire \U409_ADDRESS_DECODE.g0_i_o4Z0Z_0 ;
    wire U409_ADDRESS_DECODE_ATA_ROM_0_1;
    wire \U409_TRANSFER_ACK.CO1 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ;
    wire TM_c_1;
    wire TM_c_0;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2 ;
    wire \U409_ADDRESS_DECODE.un2_REGSPACEn_0_0_cascade_ ;
    wire A_c_19;
    wire A_c_18;
    wire \U409_ADDRESS_DECODE.REG_SPACEZ0Z_2 ;
    wire \U409_ADDRESS_DECODE.REG_SPACE_3 ;
    wire \U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0 ;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn_i;
    wire A_c_17;
    wire ATA_BASE_1;
    wire U409_ADDRESS_DECODE_un1_Z2_SPACE_7_2;
    wire A_c_16;
    wire A_c_22;
    wire ATA_BASE_0;
    wire ATA_BASE_6;
    wire \U409_TRANSFER_ACK.G_14_0_o7_2_cascade_ ;
    wire \U409_TRANSFER_ACK.G_14_0_o7_4 ;
    wire A_c_20;
    wire ATA_BASE_7;
    wire ATA_BASE_4;
    wire \U409_TRANSFER_ACK.G_14_0_o7_3 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_1_0 ;
    wire \U409_TRANSFER_ACK.N_13 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_cascade_ ;
    wire A_c_23;
    wire \U409_TRANSFER_ACK.N_24 ;
    wire \U409_TRANSFER_ACK.G_14_0_1_1 ;
    wire \U409_TRANSFER_ACK.G_14_0_1_cascade_ ;
    wire \U409_TRANSFER_ACK.G_14_0_o7_6 ;
    wire \U409_TRANSFER_ACK.G_14_0_4_cascade_ ;
    wire \U409_TRANSFER_ACK.g0_0_0_o6_4 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_out ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0_cascade_ ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ;
    wire \U409_TRANSFER_ACK.ROMENn_1_sqmuxa_0_c ;
    wire A_c_21;
    wire U409_ADDRESS_DECODE_ROMEN_1;
    wire OVL_c;
    wire \U409_ADDRESS_DECODE.LOWROMZ0Z_3 ;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn_cascade_;
    wire PORTSIZE_0_i;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_2 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net ;
    wire U409_ADDRESS_DECODE_un1_RTC_ENn;
    wire AUTOVECTOR;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0 ;
    wire AC_TACK;
    wire \U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ;
    wire \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3 ;
    wire \U409_TRANSFER_ACK.ROMENn_1_sqmuxa_d ;
    wire ROMENn_c;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_2 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire TSn_c;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn;
    wire TACKn_in;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn;
    wire BUFENn_c;
    wire U409_ADDRESS_DECODE_un2_REGSPACEn_0;
    wire U409_ADDRESS_DECODE_Z2_SPACE;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn_i;
    wire CIA_ENABLE_cascade_;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_CIACS0n_i;
    wire CIA_ENABLE;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_CIACS1n_i;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ;
    wire RESETn_c_i_g;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ;
    wire \U409_TRANSFER_ACK.N_17_mux ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6 ;
    wire \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ;
    wire TACK_OUTn;
    wire \INVU409_TRANSFER_ACK.TACK_OUTnC_net ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire \U409_ADDRESS_DECODE.un1_Z2_SPACEZ0 ;
    wire U409_ADDRESS_DECODE_ATA_ROM_EN;
    wire U409_ADDRESS_DECODE_un1_ATA_ENn_i;
    wire \U409_CIA.CLK_CIA6_4_cascade_ ;
    wire \U409_CIA.VMA_RNOZ0Z_0_cascade_ ;
    wire \U409_CIA.VMAZ0 ;
    wire AUTOCONFIG_SPACE;
    wire CIA_SPACE;
    wire TACK_EN;
    wire TCIn_1_i;
    wire CONSTANT_ONE_NET;
    wire CLK40_IN_c_g;
    wire GB_BUFFER_CLK40_IN_c_g_THRU_CO;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_3_0 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_6_0_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_1C_net ;
    wire bfn_12_9_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_5 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_6 ;
    wire \U409_CIA.un1_CIA_CLK_COUNT_3_2 ;
    wire \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_6 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_7 ;
    wire \U409_CIA.CLK_CIA6_3_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2 ;
    wire \U409_CIA.CLK_CIA6_4 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3 ;
    wire CLK28_IN_c_g;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire CLK_CIA_c;
    wire \U409_CIA.CLK_CIA_r_1_0 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_0 ;
    wire RESETn_c;
    wire RESETn_c_i;
    wire \U409_TICK.TICK603_10_cascade_ ;
    wire TICK60_c;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_8_cascade_ ;
    wire \U409_TICK.TICK603_11 ;
    wire \U409_TICK.TICK603_14 ;
    wire TICK50_c;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.TICK503_11 ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire bfn_14_5_0_;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire bfn_14_6_0_;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire bfn_14_7_0_;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire bfn_14_8_0_;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire CLK6_c_g;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__10297),
            .RESETB(N__9759),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK40_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__12505),
            .GLOBALBUFFEROUTPUT(CLK40_IN_c_g));
    IO_PAD CLK40_IN_ibuf_gb_io_iopad (
            .OE(N__12507),
            .DIN(N__12506),
            .DOUT(N__12505),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_gb_io_preio (
            .PADOEN(N__12507),
            .PADOUT(N__12506),
            .PADIN(N__12505),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__12495),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__12497),
            .DIN(N__12496),
            .DOUT(N__12495),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__12497),
            .PADOUT(N__12496),
            .PADIN(N__12495),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__12485),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__12487),
            .DIN(N__12486),
            .DOUT(N__12485),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__12487),
            .PADOUT(N__12486),
            .PADIN(N__12485),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__12476),
            .DIN(N__12475),
            .DOUT(N__12474),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__12476),
            .PADOUT(N__12475),
            .PADIN(N__12474),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__12467),
            .DIN(N__12466),
            .DOUT(N__12465),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__12467),
            .PADOUT(N__12466),
            .PADIN(N__12465),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_P1_obuf_iopad (
            .OE(N__12458),
            .DIN(N__12457),
            .DOUT(N__12456),
            .PACKAGEPIN(PIO_P1));
    defparam PIO_P1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_P1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_P1_obuf_preio (
            .PADOEN(N__12458),
            .PADOUT(N__12457),
            .PADIN(N__12456),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9786),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_7_iopad (
            .OE(N__12449),
            .DIN(N__12448),
            .DOUT(N__12447),
            .PACKAGEPIN(D[7]));
    defparam D_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_7_preio (
            .PADOEN(N__12449),
            .PADOUT(N__12448),
            .PADIN(N__12447),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4861),
            .DIN0(D_in_7),
            .DOUT0(N__4603),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__12440),
            .DIN(N__12439),
            .DOUT(N__12438),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__12440),
            .PADOUT(N__12439),
            .PADIN(N__12438),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CPUCONFn_ibuf_iopad (
            .OE(N__12431),
            .DIN(N__12430),
            .DOUT(N__12429),
            .PACKAGEPIN(CPUCONFn));
    defparam CPUCONFn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUCONFn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CPUCONFn_ibuf_preio (
            .PADOEN(N__12431),
            .PADOUT(N__12430),
            .PADIN(N__12429),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CPUCONFn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RTC_ENn_obuf_iopad (
            .OE(N__12422),
            .DIN(N__12421),
            .DOUT(N__12420),
            .PACKAGEPIN(RTC_ENn));
    defparam RTC_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RTC_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RTC_ENn_obuf_preio (
            .PADOEN(N__12422),
            .PADOUT(N__12421),
            .PADIN(N__12420),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6442),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__12413),
            .DIN(N__12412),
            .DOUT(N__12411),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__12413),
            .PADOUT(N__12412),
            .PADIN(N__12411),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ATA_MODE_P_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ATA_MODE_P_ibuf_iopad (
            .OE(N__12404),
            .DIN(N__12403),
            .DOUT(N__12402),
            .PACKAGEPIN(ATA_MODE_P));
    defparam ATA_MODE_P_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ATA_MODE_P_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ATA_MODE_P_ibuf_preio (
            .PADOEN(N__12404),
            .PADOUT(N__12403),
            .PADIN(N__12402),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PIO_P0_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_4_iopad (
            .OE(N__12395),
            .DIN(N__12394),
            .DOUT(N__12393),
            .PACKAGEPIN(D[4]));
    defparam D_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_4_preio (
            .PADOEN(N__12395),
            .PADOUT(N__12394),
            .PADIN(N__12393),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4846),
            .DIN0(D_in_4),
            .DOUT0(N__5020),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__12386),
            .DIN(N__12385),
            .DOUT(N__12384),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__12386),
            .PADOUT(N__12385),
            .PADIN(N__12384),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_1_iopad (
            .OE(N__12377),
            .DIN(N__12376),
            .DOUT(N__12375),
            .PACKAGEPIN(TM[1]));
    defparam TM_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_1_preio (
            .PADOEN(N__12377),
            .PADOUT(N__12376),
            .PADIN(N__12375),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__12368),
            .DIN(N__12367),
            .DOUT(N__12366),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__12368),
            .PADOUT(N__12367),
            .PADIN(N__12366),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_obuf_iopad (
            .OE(N__12359),
            .DIN(N__12358),
            .DOUT(N__12357),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMSPACEn_obuf_preio (
            .PADOEN(N__12359),
            .PADOUT(N__12358),
            .PADIN(N__12357),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7681),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__12350),
            .DIN(N__12349),
            .DOUT(N__12348),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__12350),
            .PADOUT(N__12349),
            .PADIN(N__12348),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ROMENn_obuf_iopad (
            .OE(N__12341),
            .DIN(N__12340),
            .DOUT(N__12339),
            .PACKAGEPIN(ROMENn));
    defparam ROMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ROMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ROMENn_obuf_preio (
            .PADOEN(N__12341),
            .PADOUT(N__12340),
            .PADIN(N__12339),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8833),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__12332),
            .DIN(N__12331),
            .DOUT(N__12330),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__12332),
            .PADOUT(N__12331),
            .PADIN(N__12330),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9874),
            .DIN0(),
            .DOUT0(N__9612),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam AUTOBOOT_ibuf_iopad.PULLUP=1'b1;
    IO_PAD AUTOBOOT_ibuf_iopad (
            .OE(N__12323),
            .DIN(N__12322),
            .DOUT(N__12321),
            .PACKAGEPIN(AUTOBOOT));
    defparam AUTOBOOT_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AUTOBOOT_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AUTOBOOT_ibuf_preio (
            .PADOEN(N__12323),
            .PADOUT(N__12322),
            .PADIN(N__12321),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AUTOBOOT_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__12314),
            .DIN(N__12313),
            .DOUT(N__12312),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__12314),
            .PADOUT(N__12313),
            .PADIN(N__12312),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__12305),
            .DIN(N__12304),
            .DOUT(N__12303),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__12305),
            .PADOUT(N__12304),
            .PADIN(N__12303),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8290),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_P2_obuf_iopad (
            .OE(N__12296),
            .DIN(N__12295),
            .DOUT(N__12294),
            .PACKAGEPIN(PIO_P2));
    defparam PIO_P2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_P2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_P2_obuf_preio (
            .PADOEN(N__12296),
            .PADOUT(N__12295),
            .PADIN(N__12294),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9785),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__12287),
            .DIN(N__12286),
            .DOUT(N__12285),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__12287),
            .PADOUT(N__12286),
            .PADIN(N__12285),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BRIDGE_ENn_obuf_iopad (
            .OE(N__12278),
            .DIN(N__12277),
            .DOUT(N__12276),
            .PACKAGEPIN(BRIDGE_ENn));
    defparam BRIDGE_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BRIDGE_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BRIDGE_ENn_obuf_preio (
            .PADOEN(N__12278),
            .PADOUT(N__12277),
            .PADIN(N__12276),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6580),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__12269),
            .DIN(N__12268),
            .DOUT(N__12267),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__12269),
            .PADOUT(N__12268),
            .PADIN(N__12267),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__12260),
            .DIN(N__12259),
            .DOUT(N__12258),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__12260),
            .PADOUT(N__12259),
            .PADIN(N__12258),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__12251),
            .DIN(N__12250),
            .DOUT(N__12249),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__12251),
            .PADOUT(N__12250),
            .PADIN(N__12249),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__12242),
            .DIN(N__12241),
            .DOUT(N__12240),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__12242),
            .PADOUT(N__12241),
            .PADIN(N__12240),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS0n_obuf_iopad (
            .OE(N__12233),
            .DIN(N__12232),
            .DOUT(N__12231),
            .PACKAGEPIN(CIACS0n));
    defparam CIACS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS0n_obuf_preio (
            .PADOEN(N__12233),
            .PADOUT(N__12232),
            .PADIN(N__12231),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9199),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__12224),
            .DIN(N__12223),
            .DOUT(N__12222),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__12224),
            .PADOUT(N__12223),
            .PADIN(N__12222),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10966),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__12215),
            .DIN(N__12214),
            .DOUT(N__12213),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__12215),
            .PADOUT(N__12214),
            .PADIN(N__12213),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_5_iopad (
            .OE(N__12206),
            .DIN(N__12205),
            .DOUT(N__12204),
            .PACKAGEPIN(D[5]));
    defparam D_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_5_preio (
            .PADOEN(N__12206),
            .PADOUT(N__12205),
            .PADIN(N__12204),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4856),
            .DIN0(D_in_5),
            .DOUT0(N__5050),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__12197),
            .DIN(N__12196),
            .DOUT(N__12195),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__12197),
            .PADOUT(N__12196),
            .PADIN(N__12195),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__12188),
            .DIN(N__12187),
            .DOUT(N__12186),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__12188),
            .PADOUT(N__12187),
            .PADIN(N__12186),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__12179),
            .DIN(N__12178),
            .DOUT(N__12177),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__12179),
            .PADOUT(N__12178),
            .PADIN(N__12177),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CONFIGENn_obuf_iopad (
            .OE(N__12170),
            .DIN(N__12169),
            .DOUT(N__12168),
            .PACKAGEPIN(CONFIGENn));
    defparam CONFIGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CONFIGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CONFIGENn_obuf_preio (
            .PADOEN(N__12170),
            .PADOUT(N__12169),
            .PADIN(N__12168),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6730),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__12161),
            .DIN(N__12160),
            .DOUT(N__12159),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__12161),
            .PADOUT(N__12160),
            .PADIN(N__12159),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10621),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__12152),
            .DIN(N__12151),
            .DOUT(N__12150),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__12152),
            .PADOUT(N__12151),
            .PADIN(N__12150),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_P0_obuf_iopad (
            .OE(N__12143),
            .DIN(N__12142),
            .DOUT(N__12141),
            .PACKAGEPIN(PIO_P0));
    defparam PIO_P0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_P0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_P0_obuf_preio (
            .PADOEN(N__12143),
            .PADOUT(N__12142),
            .PADIN(N__12141),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4465),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ATA_MODE_S_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ATA_MODE_S_ibuf_iopad (
            .OE(N__12134),
            .DIN(N__12133),
            .DOUT(N__12132),
            .PACKAGEPIN(ATA_MODE_S));
    defparam ATA_MODE_S_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ATA_MODE_S_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ATA_MODE_S_ibuf_preio (
            .PADOEN(N__12134),
            .PADOUT(N__12133),
            .PADIN(N__12132),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PIO_S0_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__12125),
            .DIN(N__12124),
            .DOUT(N__12123),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__12125),
            .PADOUT(N__12124),
            .PADIN(N__12123),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ATA_ENn_obuf_iopad (
            .OE(N__12116),
            .DIN(N__12115),
            .DOUT(N__12114),
            .PACKAGEPIN(ATA_ENn));
    defparam ATA_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ATA_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ATA_ENn_obuf_preio (
            .PADOEN(N__12116),
            .PADOUT(N__12115),
            .PADIN(N__12114),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9988),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__12107),
            .DIN(N__12106),
            .DOUT(N__12105),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__12107),
            .PADOUT(N__12106),
            .PADIN(N__12105),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS1n_obuf_iopad (
            .OE(N__12098),
            .DIN(N__12097),
            .DOUT(N__12096),
            .PACKAGEPIN(CIACS1n));
    defparam CIACS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS1n_obuf_preio (
            .PADOEN(N__12098),
            .PADOUT(N__12097),
            .PADIN(N__12096),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9154),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_obuf_iopad (
            .OE(N__12089),
            .DIN(N__12088),
            .DOUT(N__12087),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGSPACEn_obuf_preio (
            .PADOEN(N__12089),
            .PADOUT(N__12088),
            .PADIN(N__12087),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9238),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__12080),
            .DIN(N__12079),
            .DOUT(N__12078),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__12080),
            .PADOUT(N__12079),
            .PADIN(N__12078),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_CIA_obuf_iopad (
            .OE(N__12071),
            .DIN(N__12070),
            .DOUT(N__12069),
            .PACKAGEPIN(CLK_CIA));
    defparam CLK_CIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_CIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_CIA_obuf_preio (
            .PADOEN(N__12071),
            .PADOUT(N__12070),
            .PADIN(N__12069),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10441),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__12062),
            .DIN(N__12061),
            .DOUT(N__12060),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__12062),
            .PADOUT(N__12061),
            .PADIN(N__12060),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__12053),
            .DIN(N__12052),
            .DOUT(N__12051),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__12053),
            .PADOUT(N__12052),
            .PADIN(N__12051),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9873),
            .DIN0(TACKn_in),
            .DOUT0(N__9600),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__12044),
            .DIN(N__12043),
            .DOUT(N__12042),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__12044),
            .PADOUT(N__12043),
            .PADIN(N__12042),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__12035),
            .DIN(N__12034),
            .DOUT(N__12033),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__12035),
            .PADOUT(N__12034),
            .PADIN(N__12033),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9340),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_S0_obuf_iopad (
            .OE(N__12026),
            .DIN(N__12025),
            .DOUT(N__12024),
            .PACKAGEPIN(PIO_S0));
    defparam PIO_S0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_S0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_S0_obuf_preio (
            .PADOEN(N__12026),
            .PADOUT(N__12025),
            .PADIN(N__12024),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4444),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__12017),
            .DIN(N__12016),
            .DOUT(N__12015),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__12017),
            .PADOUT(N__12016),
            .PADIN(N__12015),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_S2_obuf_iopad (
            .OE(N__12008),
            .DIN(N__12007),
            .DOUT(N__12006),
            .PACKAGEPIN(PIO_S2));
    defparam PIO_S2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_S2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_S2_obuf_preio (
            .PADOEN(N__12008),
            .PADOUT(N__12007),
            .PADIN(N__12006),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9799),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_6_iopad (
            .OE(N__11999),
            .DIN(N__11998),
            .DOUT(N__11997),
            .PACKAGEPIN(D[6]));
    defparam D_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_6_preio (
            .PADOEN(N__11999),
            .PADOUT(N__11998),
            .PADIN(N__11997),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4857),
            .DIN0(D_in_6),
            .DOUT0(N__5872),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11990),
            .DIN(N__11989),
            .DOUT(N__11988),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11990),
            .PADOUT(N__11989),
            .PADIN(N__11988),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__11981),
            .DIN(N__11980),
            .DOUT(N__11979),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__11981),
            .PADOUT(N__11980),
            .PADIN(N__11979),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_S1_obuf_iopad (
            .OE(N__11972),
            .DIN(N__11971),
            .DOUT(N__11970),
            .PACKAGEPIN(PIO_S1));
    defparam PIO_S1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_S1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_S1_obuf_preio (
            .PADOEN(N__11972),
            .PADOUT(N__11971),
            .PADIN(N__11970),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9798),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_0_iopad (
            .OE(N__11963),
            .DIN(N__11962),
            .DOUT(N__11961),
            .PACKAGEPIN(TM[0]));
    defparam TM_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_0_preio (
            .PADOEN(N__11963),
            .PADOUT(N__11962),
            .PADIN(N__11961),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11954),
            .DIN(N__11953),
            .DOUT(N__11952),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11954),
            .PADOUT(N__11953),
            .PADIN(N__11952),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11945),
            .DIN(N__11944),
            .DOUT(N__11943),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11945),
            .PADOUT(N__11944),
            .PADIN(N__11943),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11936),
            .DIN(N__11935),
            .DOUT(N__11934),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11936),
            .PADOUT(N__11935),
            .PADIN(N__11934),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__11927),
            .DIN(N__11926),
            .DOUT(N__11925),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__11927),
            .PADOUT(N__11926),
            .PADIN(N__11925),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__11918),
            .DIN(N__11917),
            .DOUT(N__11916),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__11918),
            .PADOUT(N__11917),
            .PADIN(N__11916),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__11909),
            .DIN(N__11908),
            .DOUT(N__11907),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__11909),
            .PADOUT(N__11908),
            .PADIN(N__11907),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9823),
            .DIN0(),
            .DOUT0(N__9613),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2885 (
            .O(N__11890),
            .I(N__11886));
    InMux I__2884 (
            .O(N__11889),
            .I(N__11883));
    LocalMux I__2883 (
            .O(N__11886),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__2882 (
            .O(N__11883),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    InMux I__2881 (
            .O(N__11878),
            .I(N__11875));
    LocalMux I__2880 (
            .O(N__11875),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__2879 (
            .O(N__11872),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__2878 (
            .O(N__11869),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__2877 (
            .O(N__11866),
            .I(N__11862));
    InMux I__2876 (
            .O(N__11865),
            .I(N__11859));
    LocalMux I__2875 (
            .O(N__11862),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__2874 (
            .O(N__11859),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    ClkMux I__2873 (
            .O(N__11854),
            .I(N__11827));
    ClkMux I__2872 (
            .O(N__11853),
            .I(N__11827));
    ClkMux I__2871 (
            .O(N__11852),
            .I(N__11827));
    ClkMux I__2870 (
            .O(N__11851),
            .I(N__11827));
    ClkMux I__2869 (
            .O(N__11850),
            .I(N__11827));
    ClkMux I__2868 (
            .O(N__11849),
            .I(N__11827));
    ClkMux I__2867 (
            .O(N__11848),
            .I(N__11827));
    ClkMux I__2866 (
            .O(N__11847),
            .I(N__11827));
    ClkMux I__2865 (
            .O(N__11846),
            .I(N__11827));
    GlobalMux I__2864 (
            .O(N__11827),
            .I(N__11824));
    gio2CtrlBuf I__2863 (
            .O(N__11824),
            .I(CLK6_c_g));
    InMux I__2862 (
            .O(N__11821),
            .I(N__11817));
    InMux I__2861 (
            .O(N__11820),
            .I(N__11814));
    LocalMux I__2860 (
            .O(N__11817),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__2859 (
            .O(N__11814),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    InMux I__2858 (
            .O(N__11809),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__2857 (
            .O(N__11806),
            .I(N__11802));
    InMux I__2856 (
            .O(N__11805),
            .I(N__11799));
    LocalMux I__2855 (
            .O(N__11802),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__2854 (
            .O(N__11799),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__2853 (
            .O(N__11794),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__2852 (
            .O(N__11791),
            .I(N__11787));
    InMux I__2851 (
            .O(N__11790),
            .I(N__11784));
    LocalMux I__2850 (
            .O(N__11787),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__2849 (
            .O(N__11784),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    InMux I__2848 (
            .O(N__11779),
            .I(N__11776));
    LocalMux I__2847 (
            .O(N__11776),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__2846 (
            .O(N__11773),
            .I(bfn_14_8_0_));
    InMux I__2845 (
            .O(N__11770),
            .I(N__11766));
    InMux I__2844 (
            .O(N__11769),
            .I(N__11763));
    LocalMux I__2843 (
            .O(N__11766),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__2842 (
            .O(N__11763),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    InMux I__2841 (
            .O(N__11758),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    CascadeMux I__2840 (
            .O(N__11755),
            .I(N__11752));
    InMux I__2839 (
            .O(N__11752),
            .I(N__11748));
    InMux I__2838 (
            .O(N__11751),
            .I(N__11745));
    LocalMux I__2837 (
            .O(N__11748),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__2836 (
            .O(N__11745),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__2835 (
            .O(N__11740),
            .I(N__11737));
    LocalMux I__2834 (
            .O(N__11737),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__2833 (
            .O(N__11734),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__2832 (
            .O(N__11731),
            .I(N__11727));
    InMux I__2831 (
            .O(N__11730),
            .I(N__11724));
    LocalMux I__2830 (
            .O(N__11727),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__2829 (
            .O(N__11724),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    InMux I__2828 (
            .O(N__11719),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__2827 (
            .O(N__11716),
            .I(N__11712));
    InMux I__2826 (
            .O(N__11715),
            .I(N__11709));
    LocalMux I__2825 (
            .O(N__11712),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__2824 (
            .O(N__11709),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__2823 (
            .O(N__11704),
            .I(N__11701));
    LocalMux I__2822 (
            .O(N__11701),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__2821 (
            .O(N__11698),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__2820 (
            .O(N__11695),
            .I(N__11691));
    InMux I__2819 (
            .O(N__11694),
            .I(N__11688));
    LocalMux I__2818 (
            .O(N__11691),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__2817 (
            .O(N__11688),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    InMux I__2816 (
            .O(N__11683),
            .I(N__11680));
    LocalMux I__2815 (
            .O(N__11680),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__2814 (
            .O(N__11677),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__2813 (
            .O(N__11674),
            .I(N__11670));
    InMux I__2812 (
            .O(N__11673),
            .I(N__11667));
    LocalMux I__2811 (
            .O(N__11670),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__2810 (
            .O(N__11667),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__2809 (
            .O(N__11662),
            .I(N__11659));
    LocalMux I__2808 (
            .O(N__11659),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__2807 (
            .O(N__11656),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__2806 (
            .O(N__11653),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__2805 (
            .O(N__11650),
            .I(N__11646));
    InMux I__2804 (
            .O(N__11649),
            .I(N__11643));
    LocalMux I__2803 (
            .O(N__11646),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__2802 (
            .O(N__11643),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    CascadeMux I__2801 (
            .O(N__11638),
            .I(N__11634));
    InMux I__2800 (
            .O(N__11637),
            .I(N__11628));
    InMux I__2799 (
            .O(N__11634),
            .I(N__11628));
    InMux I__2798 (
            .O(N__11633),
            .I(N__11625));
    LocalMux I__2797 (
            .O(N__11628),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__2796 (
            .O(N__11625),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    CascadeMux I__2795 (
            .O(N__11620),
            .I(N__11614));
    InMux I__2794 (
            .O(N__11619),
            .I(N__11611));
    InMux I__2793 (
            .O(N__11618),
            .I(N__11606));
    InMux I__2792 (
            .O(N__11617),
            .I(N__11606));
    InMux I__2791 (
            .O(N__11614),
            .I(N__11603));
    LocalMux I__2790 (
            .O(N__11611),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2789 (
            .O(N__11606),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2788 (
            .O(N__11603),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__2787 (
            .O(N__11596),
            .I(N__11592));
    InMux I__2786 (
            .O(N__11595),
            .I(N__11589));
    LocalMux I__2785 (
            .O(N__11592),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__2784 (
            .O(N__11589),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__2783 (
            .O(N__11584),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__2782 (
            .O(N__11581),
            .I(N__11577));
    InMux I__2781 (
            .O(N__11580),
            .I(N__11574));
    LocalMux I__2780 (
            .O(N__11577),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__2779 (
            .O(N__11574),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__2778 (
            .O(N__11569),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    InMux I__2777 (
            .O(N__11566),
            .I(N__11562));
    InMux I__2776 (
            .O(N__11565),
            .I(N__11559));
    LocalMux I__2775 (
            .O(N__11562),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__2774 (
            .O(N__11559),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    InMux I__2773 (
            .O(N__11554),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    CascadeMux I__2772 (
            .O(N__11551),
            .I(N__11548));
    InMux I__2771 (
            .O(N__11548),
            .I(N__11544));
    InMux I__2770 (
            .O(N__11547),
            .I(N__11541));
    LocalMux I__2769 (
            .O(N__11544),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__2768 (
            .O(N__11541),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    CascadeMux I__2767 (
            .O(N__11536),
            .I(N__11533));
    InMux I__2766 (
            .O(N__11533),
            .I(N__11530));
    LocalMux I__2765 (
            .O(N__11530),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__2764 (
            .O(N__11527),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    InMux I__2763 (
            .O(N__11524),
            .I(N__11521));
    LocalMux I__2762 (
            .O(N__11521),
            .I(N__11517));
    InMux I__2761 (
            .O(N__11520),
            .I(N__11514));
    Odrv4 I__2760 (
            .O(N__11517),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__2759 (
            .O(N__11514),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    CascadeMux I__2758 (
            .O(N__11509),
            .I(N__11506));
    InMux I__2757 (
            .O(N__11506),
            .I(N__11503));
    LocalMux I__2756 (
            .O(N__11503),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__2755 (
            .O(N__11500),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__2754 (
            .O(N__11497),
            .I(N__11494));
    LocalMux I__2753 (
            .O(N__11494),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__2752 (
            .O(N__11491),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__2751 (
            .O(N__11488),
            .I(N__11484));
    InMux I__2750 (
            .O(N__11487),
            .I(N__11481));
    LocalMux I__2749 (
            .O(N__11484),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__2748 (
            .O(N__11481),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__2747 (
            .O(N__11476),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__2746 (
            .O(N__11473),
            .I(N__11469));
    InMux I__2745 (
            .O(N__11472),
            .I(N__11466));
    LocalMux I__2744 (
            .O(N__11469),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__2743 (
            .O(N__11466),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    CascadeMux I__2742 (
            .O(N__11461),
            .I(N__11458));
    InMux I__2741 (
            .O(N__11458),
            .I(N__11455));
    LocalMux I__2740 (
            .O(N__11455),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__2739 (
            .O(N__11452),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__2738 (
            .O(N__11449),
            .I(N__11445));
    InMux I__2737 (
            .O(N__11448),
            .I(N__11442));
    LocalMux I__2736 (
            .O(N__11445),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__2735 (
            .O(N__11442),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    CascadeMux I__2734 (
            .O(N__11437),
            .I(N__11434));
    InMux I__2733 (
            .O(N__11434),
            .I(N__11431));
    LocalMux I__2732 (
            .O(N__11431),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__2731 (
            .O(N__11428),
            .I(bfn_14_6_0_));
    InMux I__2730 (
            .O(N__11425),
            .I(N__11421));
    InMux I__2729 (
            .O(N__11424),
            .I(N__11418));
    LocalMux I__2728 (
            .O(N__11421),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__2727 (
            .O(N__11418),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    InMux I__2726 (
            .O(N__11413),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__2725 (
            .O(N__11410),
            .I(N__11406));
    InMux I__2724 (
            .O(N__11409),
            .I(N__11403));
    LocalMux I__2723 (
            .O(N__11406),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__2722 (
            .O(N__11403),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    InMux I__2721 (
            .O(N__11398),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__2720 (
            .O(N__11395),
            .I(N__11391));
    InMux I__2719 (
            .O(N__11394),
            .I(N__11388));
    LocalMux I__2718 (
            .O(N__11391),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__2717 (
            .O(N__11388),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__2716 (
            .O(N__11383),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__2715 (
            .O(N__11380),
            .I(N__11376));
    InMux I__2714 (
            .O(N__11379),
            .I(N__11373));
    LocalMux I__2713 (
            .O(N__11376),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__2712 (
            .O(N__11373),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__2711 (
            .O(N__11368),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    CascadeMux I__2710 (
            .O(N__11365),
            .I(N__11362));
    InMux I__2709 (
            .O(N__11362),
            .I(N__11358));
    InMux I__2708 (
            .O(N__11361),
            .I(N__11355));
    LocalMux I__2707 (
            .O(N__11358),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__2706 (
            .O(N__11355),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    InMux I__2705 (
            .O(N__11350),
            .I(N__11347));
    LocalMux I__2704 (
            .O(N__11347),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__2703 (
            .O(N__11344),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__2702 (
            .O(N__11341),
            .I(N__11338));
    LocalMux I__2701 (
            .O(N__11338),
            .I(\U409_TICK.TICK503_11 ));
    CascadeMux I__2700 (
            .O(N__11335),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    CascadeMux I__2699 (
            .O(N__11332),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    CascadeMux I__2698 (
            .O(N__11329),
            .I(N__11325));
    InMux I__2697 (
            .O(N__11328),
            .I(N__11316));
    InMux I__2696 (
            .O(N__11325),
            .I(N__11307));
    InMux I__2695 (
            .O(N__11324),
            .I(N__11307));
    InMux I__2694 (
            .O(N__11323),
            .I(N__11307));
    InMux I__2693 (
            .O(N__11322),
            .I(N__11307));
    InMux I__2692 (
            .O(N__11321),
            .I(N__11300));
    InMux I__2691 (
            .O(N__11320),
            .I(N__11300));
    InMux I__2690 (
            .O(N__11319),
            .I(N__11300));
    LocalMux I__2689 (
            .O(N__11316),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__2688 (
            .O(N__11307),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__2687 (
            .O(N__11300),
            .I(\U409_TICK.TICK503_10 ));
    InMux I__2686 (
            .O(N__11293),
            .I(N__11283));
    InMux I__2685 (
            .O(N__11292),
            .I(N__11274));
    InMux I__2684 (
            .O(N__11291),
            .I(N__11274));
    InMux I__2683 (
            .O(N__11290),
            .I(N__11274));
    InMux I__2682 (
            .O(N__11289),
            .I(N__11274));
    InMux I__2681 (
            .O(N__11288),
            .I(N__11267));
    InMux I__2680 (
            .O(N__11287),
            .I(N__11267));
    InMux I__2679 (
            .O(N__11286),
            .I(N__11267));
    LocalMux I__2678 (
            .O(N__11283),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__2677 (
            .O(N__11274),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__2676 (
            .O(N__11267),
            .I(\U409_TICK.TICK503_14 ));
    CascadeMux I__2675 (
            .O(N__11260),
            .I(N__11254));
    CascadeMux I__2674 (
            .O(N__11259),
            .I(N__11250));
    CascadeMux I__2673 (
            .O(N__11258),
            .I(N__11244));
    InMux I__2672 (
            .O(N__11257),
            .I(N__11241));
    InMux I__2671 (
            .O(N__11254),
            .I(N__11236));
    InMux I__2670 (
            .O(N__11253),
            .I(N__11236));
    InMux I__2669 (
            .O(N__11250),
            .I(N__11233));
    InMux I__2668 (
            .O(N__11249),
            .I(N__11224));
    InMux I__2667 (
            .O(N__11248),
            .I(N__11224));
    InMux I__2666 (
            .O(N__11247),
            .I(N__11224));
    InMux I__2665 (
            .O(N__11244),
            .I(N__11224));
    LocalMux I__2664 (
            .O(N__11241),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__2663 (
            .O(N__11236),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__2662 (
            .O(N__11233),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__2661 (
            .O(N__11224),
            .I(\U409_TICK.TICK503_9 ));
    InMux I__2660 (
            .O(N__11215),
            .I(N__11211));
    InMux I__2659 (
            .O(N__11214),
            .I(N__11207));
    LocalMux I__2658 (
            .O(N__11211),
            .I(N__11204));
    InMux I__2657 (
            .O(N__11210),
            .I(N__11201));
    LocalMux I__2656 (
            .O(N__11207),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    Odrv4 I__2655 (
            .O(N__11204),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__2654 (
            .O(N__11201),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    CascadeMux I__2653 (
            .O(N__11194),
            .I(N__11188));
    InMux I__2652 (
            .O(N__11193),
            .I(N__11185));
    InMux I__2651 (
            .O(N__11192),
            .I(N__11180));
    InMux I__2650 (
            .O(N__11191),
            .I(N__11180));
    InMux I__2649 (
            .O(N__11188),
            .I(N__11177));
    LocalMux I__2648 (
            .O(N__11185),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__2647 (
            .O(N__11180),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__2646 (
            .O(N__11177),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    CascadeMux I__2645 (
            .O(N__11170),
            .I(N__11167));
    InMux I__2644 (
            .O(N__11167),
            .I(N__11163));
    InMux I__2643 (
            .O(N__11166),
            .I(N__11160));
    LocalMux I__2642 (
            .O(N__11163),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__2641 (
            .O(N__11160),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    InMux I__2640 (
            .O(N__11155),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__2639 (
            .O(N__11152),
            .I(N__11148));
    InMux I__2638 (
            .O(N__11151),
            .I(N__11145));
    LocalMux I__2637 (
            .O(N__11148),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__2636 (
            .O(N__11145),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    InMux I__2635 (
            .O(N__11140),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__2634 (
            .O(N__11137),
            .I(N__11133));
    InMux I__2633 (
            .O(N__11136),
            .I(N__11130));
    LocalMux I__2632 (
            .O(N__11133),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__2631 (
            .O(N__11130),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__2630 (
            .O(N__11125),
            .I(N__11122));
    LocalMux I__2629 (
            .O(N__11122),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__2628 (
            .O(N__11119),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    CascadeMux I__2627 (
            .O(N__11116),
            .I(N__11113));
    InMux I__2626 (
            .O(N__11113),
            .I(N__11109));
    InMux I__2625 (
            .O(N__11112),
            .I(N__11106));
    LocalMux I__2624 (
            .O(N__11109),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__2623 (
            .O(N__11106),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__2622 (
            .O(N__11101),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    InMux I__2621 (
            .O(N__11098),
            .I(N__11094));
    InMux I__2620 (
            .O(N__11097),
            .I(N__11091));
    LocalMux I__2619 (
            .O(N__11094),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__2618 (
            .O(N__11091),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    CascadeMux I__2617 (
            .O(N__11086),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    CascadeMux I__2616 (
            .O(N__11083),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    CascadeMux I__2615 (
            .O(N__11080),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    CascadeMux I__2614 (
            .O(N__11077),
            .I(N__11070));
    InMux I__2613 (
            .O(N__11076),
            .I(N__11059));
    InMux I__2612 (
            .O(N__11075),
            .I(N__11059));
    InMux I__2611 (
            .O(N__11074),
            .I(N__11059));
    InMux I__2610 (
            .O(N__11073),
            .I(N__11059));
    InMux I__2609 (
            .O(N__11070),
            .I(N__11052));
    InMux I__2608 (
            .O(N__11069),
            .I(N__11052));
    InMux I__2607 (
            .O(N__11068),
            .I(N__11052));
    LocalMux I__2606 (
            .O(N__11059),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__2605 (
            .O(N__11052),
            .I(\U409_TICK.TICK603_10 ));
    CascadeMux I__2604 (
            .O(N__11047),
            .I(N__11038));
    CascadeMux I__2603 (
            .O(N__11046),
            .I(N__11035));
    InMux I__2602 (
            .O(N__11045),
            .I(N__11032));
    InMux I__2601 (
            .O(N__11044),
            .I(N__11025));
    InMux I__2600 (
            .O(N__11043),
            .I(N__11025));
    InMux I__2599 (
            .O(N__11042),
            .I(N__11025));
    InMux I__2598 (
            .O(N__11041),
            .I(N__11018));
    InMux I__2597 (
            .O(N__11038),
            .I(N__11018));
    InMux I__2596 (
            .O(N__11035),
            .I(N__11018));
    LocalMux I__2595 (
            .O(N__11032),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__2594 (
            .O(N__11025),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__2593 (
            .O(N__11018),
            .I(\U409_TICK.TICK603_9 ));
    CascadeMux I__2592 (
            .O(N__11011),
            .I(\U409_TICK.TICK603_8_cascade_ ));
    InMux I__2591 (
            .O(N__11008),
            .I(N__11005));
    LocalMux I__2590 (
            .O(N__11005),
            .I(\U409_TICK.TICK603_11 ));
    CascadeMux I__2589 (
            .O(N__11002),
            .I(N__10999));
    InMux I__2588 (
            .O(N__10999),
            .I(N__10989));
    InMux I__2587 (
            .O(N__10998),
            .I(N__10982));
    InMux I__2586 (
            .O(N__10997),
            .I(N__10982));
    InMux I__2585 (
            .O(N__10996),
            .I(N__10982));
    InMux I__2584 (
            .O(N__10995),
            .I(N__10973));
    InMux I__2583 (
            .O(N__10994),
            .I(N__10973));
    InMux I__2582 (
            .O(N__10993),
            .I(N__10973));
    InMux I__2581 (
            .O(N__10992),
            .I(N__10973));
    LocalMux I__2580 (
            .O(N__10989),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__2579 (
            .O(N__10982),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__2578 (
            .O(N__10973),
            .I(\U409_TICK.TICK603_14 ));
    IoInMux I__2577 (
            .O(N__10966),
            .I(N__10963));
    LocalMux I__2576 (
            .O(N__10963),
            .I(N__10960));
    Span12Mux_s0_v I__2575 (
            .O(N__10960),
            .I(N__10957));
    Span12Mux_v I__2574 (
            .O(N__10957),
            .I(N__10953));
    InMux I__2573 (
            .O(N__10956),
            .I(N__10950));
    Odrv12 I__2572 (
            .O(N__10953),
            .I(TICK50_c));
    LocalMux I__2571 (
            .O(N__10950),
            .I(TICK50_c));
    InMux I__2570 (
            .O(N__10945),
            .I(N__10937));
    InMux I__2569 (
            .O(N__10944),
            .I(N__10937));
    InMux I__2568 (
            .O(N__10943),
            .I(N__10932));
    InMux I__2567 (
            .O(N__10942),
            .I(N__10932));
    LocalMux I__2566 (
            .O(N__10937),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__2565 (
            .O(N__10932),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    InMux I__2564 (
            .O(N__10927),
            .I(N__10919));
    InMux I__2563 (
            .O(N__10926),
            .I(N__10919));
    InMux I__2562 (
            .O(N__10925),
            .I(N__10914));
    InMux I__2561 (
            .O(N__10924),
            .I(N__10914));
    LocalMux I__2560 (
            .O(N__10919),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__2559 (
            .O(N__10914),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    CascadeMux I__2558 (
            .O(N__10909),
            .I(N__10904));
    CascadeMux I__2557 (
            .O(N__10908),
            .I(N__10900));
    InMux I__2556 (
            .O(N__10907),
            .I(N__10895));
    InMux I__2555 (
            .O(N__10904),
            .I(N__10895));
    InMux I__2554 (
            .O(N__10903),
            .I(N__10890));
    InMux I__2553 (
            .O(N__10900),
            .I(N__10890));
    LocalMux I__2552 (
            .O(N__10895),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__2551 (
            .O(N__10890),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    CascadeMux I__2550 (
            .O(N__10885),
            .I(N__10877));
    InMux I__2549 (
            .O(N__10884),
            .I(N__10874));
    InMux I__2548 (
            .O(N__10883),
            .I(N__10871));
    InMux I__2547 (
            .O(N__10882),
            .I(N__10866));
    InMux I__2546 (
            .O(N__10881),
            .I(N__10866));
    InMux I__2545 (
            .O(N__10880),
            .I(N__10861));
    InMux I__2544 (
            .O(N__10877),
            .I(N__10861));
    LocalMux I__2543 (
            .O(N__10874),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__2542 (
            .O(N__10871),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__2541 (
            .O(N__10866),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__2540 (
            .O(N__10861),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    InMux I__2539 (
            .O(N__10852),
            .I(N__10848));
    InMux I__2538 (
            .O(N__10851),
            .I(N__10845));
    LocalMux I__2537 (
            .O(N__10848),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0 ));
    LocalMux I__2536 (
            .O(N__10845),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0 ));
    InMux I__2535 (
            .O(N__10840),
            .I(N__10837));
    LocalMux I__2534 (
            .O(N__10837),
            .I(N__10829));
    InMux I__2533 (
            .O(N__10836),
            .I(N__10826));
    CascadeMux I__2532 (
            .O(N__10835),
            .I(N__10819));
    CascadeMux I__2531 (
            .O(N__10834),
            .I(N__10816));
    InMux I__2530 (
            .O(N__10833),
            .I(N__10813));
    InMux I__2529 (
            .O(N__10832),
            .I(N__10810));
    Span4Mux_v I__2528 (
            .O(N__10829),
            .I(N__10803));
    LocalMux I__2527 (
            .O(N__10826),
            .I(N__10803));
    InMux I__2526 (
            .O(N__10825),
            .I(N__10796));
    InMux I__2525 (
            .O(N__10824),
            .I(N__10796));
    InMux I__2524 (
            .O(N__10823),
            .I(N__10796));
    InMux I__2523 (
            .O(N__10822),
            .I(N__10793));
    InMux I__2522 (
            .O(N__10819),
            .I(N__10788));
    InMux I__2521 (
            .O(N__10816),
            .I(N__10788));
    LocalMux I__2520 (
            .O(N__10813),
            .I(N__10783));
    LocalMux I__2519 (
            .O(N__10810),
            .I(N__10783));
    InMux I__2518 (
            .O(N__10809),
            .I(N__10780));
    CascadeMux I__2517 (
            .O(N__10808),
            .I(N__10777));
    Span4Mux_v I__2516 (
            .O(N__10803),
            .I(N__10773));
    LocalMux I__2515 (
            .O(N__10796),
            .I(N__10768));
    LocalMux I__2514 (
            .O(N__10793),
            .I(N__10768));
    LocalMux I__2513 (
            .O(N__10788),
            .I(N__10764));
    Span4Mux_v I__2512 (
            .O(N__10783),
            .I(N__10759));
    LocalMux I__2511 (
            .O(N__10780),
            .I(N__10759));
    InMux I__2510 (
            .O(N__10777),
            .I(N__10756));
    InMux I__2509 (
            .O(N__10776),
            .I(N__10753));
    Span4Mux_v I__2508 (
            .O(N__10773),
            .I(N__10746));
    Span4Mux_v I__2507 (
            .O(N__10768),
            .I(N__10746));
    InMux I__2506 (
            .O(N__10767),
            .I(N__10742));
    Span4Mux_v I__2505 (
            .O(N__10764),
            .I(N__10730));
    Span4Mux_h I__2504 (
            .O(N__10759),
            .I(N__10730));
    LocalMux I__2503 (
            .O(N__10756),
            .I(N__10730));
    LocalMux I__2502 (
            .O(N__10753),
            .I(N__10730));
    InMux I__2501 (
            .O(N__10752),
            .I(N__10725));
    InMux I__2500 (
            .O(N__10751),
            .I(N__10725));
    Span4Mux_h I__2499 (
            .O(N__10746),
            .I(N__10721));
    InMux I__2498 (
            .O(N__10745),
            .I(N__10718));
    LocalMux I__2497 (
            .O(N__10742),
            .I(N__10715));
    InMux I__2496 (
            .O(N__10741),
            .I(N__10711));
    InMux I__2495 (
            .O(N__10740),
            .I(N__10708));
    InMux I__2494 (
            .O(N__10739),
            .I(N__10705));
    Span4Mux_v I__2493 (
            .O(N__10730),
            .I(N__10702));
    LocalMux I__2492 (
            .O(N__10725),
            .I(N__10699));
    InMux I__2491 (
            .O(N__10724),
            .I(N__10696));
    Span4Mux_h I__2490 (
            .O(N__10721),
            .I(N__10692));
    LocalMux I__2489 (
            .O(N__10718),
            .I(N__10689));
    Span4Mux_h I__2488 (
            .O(N__10715),
            .I(N__10686));
    InMux I__2487 (
            .O(N__10714),
            .I(N__10683));
    LocalMux I__2486 (
            .O(N__10711),
            .I(N__10676));
    LocalMux I__2485 (
            .O(N__10708),
            .I(N__10676));
    LocalMux I__2484 (
            .O(N__10705),
            .I(N__10676));
    Span4Mux_h I__2483 (
            .O(N__10702),
            .I(N__10669));
    Span4Mux_h I__2482 (
            .O(N__10699),
            .I(N__10669));
    LocalMux I__2481 (
            .O(N__10696),
            .I(N__10669));
    InMux I__2480 (
            .O(N__10695),
            .I(N__10666));
    Span4Mux_v I__2479 (
            .O(N__10692),
            .I(N__10663));
    Span12Mux_s11_v I__2478 (
            .O(N__10689),
            .I(N__10656));
    Sp12to4 I__2477 (
            .O(N__10686),
            .I(N__10656));
    LocalMux I__2476 (
            .O(N__10683),
            .I(N__10656));
    Span4Mux_v I__2475 (
            .O(N__10676),
            .I(N__10649));
    Span4Mux_v I__2474 (
            .O(N__10669),
            .I(N__10649));
    LocalMux I__2473 (
            .O(N__10666),
            .I(N__10649));
    Sp12to4 I__2472 (
            .O(N__10663),
            .I(N__10642));
    Span12Mux_v I__2471 (
            .O(N__10656),
            .I(N__10642));
    Sp12to4 I__2470 (
            .O(N__10649),
            .I(N__10642));
    Span12Mux_h I__2469 (
            .O(N__10642),
            .I(N__10639));
    Odrv12 I__2468 (
            .O(N__10639),
            .I(RESETn_c));
    IoInMux I__2467 (
            .O(N__10636),
            .I(N__10633));
    LocalMux I__2466 (
            .O(N__10633),
            .I(N__10630));
    Span12Mux_s2_v I__2465 (
            .O(N__10630),
            .I(N__10627));
    Odrv12 I__2464 (
            .O(N__10627),
            .I(RESETn_c_i));
    CascadeMux I__2463 (
            .O(N__10624),
            .I(\U409_TICK.TICK603_10_cascade_ ));
    IoInMux I__2462 (
            .O(N__10621),
            .I(N__10618));
    LocalMux I__2461 (
            .O(N__10618),
            .I(N__10615));
    Span4Mux_s3_v I__2460 (
            .O(N__10615),
            .I(N__10612));
    Span4Mux_v I__2459 (
            .O(N__10612),
            .I(N__10609));
    Span4Mux_h I__2458 (
            .O(N__10609),
            .I(N__10605));
    InMux I__2457 (
            .O(N__10608),
            .I(N__10602));
    Odrv4 I__2456 (
            .O(N__10605),
            .I(TICK60_c));
    LocalMux I__2455 (
            .O(N__10602),
            .I(TICK60_c));
    InMux I__2454 (
            .O(N__10597),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ));
    InMux I__2453 (
            .O(N__10594),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ));
    InMux I__2452 (
            .O(N__10591),
            .I(N__10588));
    LocalMux I__2451 (
            .O(N__10588),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_3_2 ));
    InMux I__2450 (
            .O(N__10585),
            .I(N__10582));
    LocalMux I__2449 (
            .O(N__10582),
            .I(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5 ));
    InMux I__2448 (
            .O(N__10579),
            .I(N__10574));
    InMux I__2447 (
            .O(N__10578),
            .I(N__10571));
    InMux I__2446 (
            .O(N__10577),
            .I(N__10568));
    LocalMux I__2445 (
            .O(N__10574),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__2444 (
            .O(N__10571),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__2443 (
            .O(N__10568),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    CascadeMux I__2442 (
            .O(N__10561),
            .I(N__10557));
    InMux I__2441 (
            .O(N__10560),
            .I(N__10553));
    InMux I__2440 (
            .O(N__10557),
            .I(N__10550));
    InMux I__2439 (
            .O(N__10556),
            .I(N__10547));
    LocalMux I__2438 (
            .O(N__10553),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__2437 (
            .O(N__10550),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__2436 (
            .O(N__10547),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    CascadeMux I__2435 (
            .O(N__10540),
            .I(\U409_CIA.CLK_CIA6_3_cascade_ ));
    InMux I__2434 (
            .O(N__10537),
            .I(N__10529));
    InMux I__2433 (
            .O(N__10536),
            .I(N__10524));
    InMux I__2432 (
            .O(N__10535),
            .I(N__10524));
    InMux I__2431 (
            .O(N__10534),
            .I(N__10519));
    InMux I__2430 (
            .O(N__10533),
            .I(N__10519));
    InMux I__2429 (
            .O(N__10532),
            .I(N__10516));
    LocalMux I__2428 (
            .O(N__10529),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__2427 (
            .O(N__10524),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__2426 (
            .O(N__10519),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__2425 (
            .O(N__10516),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    InMux I__2424 (
            .O(N__10507),
            .I(N__10504));
    LocalMux I__2423 (
            .O(N__10504),
            .I(\U409_CIA.CIA_CLK_COUNT11_2 ));
    CascadeMux I__2422 (
            .O(N__10501),
            .I(N__10498));
    InMux I__2421 (
            .O(N__10498),
            .I(N__10492));
    InMux I__2420 (
            .O(N__10497),
            .I(N__10492));
    LocalMux I__2419 (
            .O(N__10492),
            .I(\U409_CIA.CLK_CIA6_4 ));
    CascadeMux I__2418 (
            .O(N__10489),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_cascade_ ));
    InMux I__2417 (
            .O(N__10486),
            .I(N__10483));
    LocalMux I__2416 (
            .O(N__10483),
            .I(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3 ));
    ClkMux I__2415 (
            .O(N__10480),
            .I(N__10468));
    ClkMux I__2414 (
            .O(N__10479),
            .I(N__10468));
    ClkMux I__2413 (
            .O(N__10478),
            .I(N__10468));
    ClkMux I__2412 (
            .O(N__10477),
            .I(N__10468));
    GlobalMux I__2411 (
            .O(N__10468),
            .I(N__10465));
    gio2CtrlBuf I__2410 (
            .O(N__10465),
            .I(CLK28_IN_c_g));
    InMux I__2409 (
            .O(N__10462),
            .I(N__10456));
    InMux I__2408 (
            .O(N__10461),
            .I(N__10451));
    InMux I__2407 (
            .O(N__10460),
            .I(N__10451));
    InMux I__2406 (
            .O(N__10459),
            .I(N__10448));
    LocalMux I__2405 (
            .O(N__10456),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__2404 (
            .O(N__10451),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__2403 (
            .O(N__10448),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    IoInMux I__2402 (
            .O(N__10441),
            .I(N__10438));
    LocalMux I__2401 (
            .O(N__10438),
            .I(N__10435));
    Span4Mux_s2_v I__2400 (
            .O(N__10435),
            .I(N__10432));
    Span4Mux_h I__2399 (
            .O(N__10432),
            .I(N__10428));
    InMux I__2398 (
            .O(N__10431),
            .I(N__10425));
    Span4Mux_v I__2397 (
            .O(N__10428),
            .I(N__10421));
    LocalMux I__2396 (
            .O(N__10425),
            .I(N__10418));
    CascadeMux I__2395 (
            .O(N__10424),
            .I(N__10414));
    Sp12to4 I__2394 (
            .O(N__10421),
            .I(N__10409));
    Span12Mux_h I__2393 (
            .O(N__10418),
            .I(N__10409));
    InMux I__2392 (
            .O(N__10417),
            .I(N__10404));
    InMux I__2391 (
            .O(N__10414),
            .I(N__10404));
    Odrv12 I__2390 (
            .O(N__10409),
            .I(CLK_CIA_c));
    LocalMux I__2389 (
            .O(N__10404),
            .I(CLK_CIA_c));
    InMux I__2388 (
            .O(N__10399),
            .I(N__10396));
    LocalMux I__2387 (
            .O(N__10396),
            .I(\U409_CIA.CLK_CIA_r_1_0 ));
    CascadeMux I__2386 (
            .O(N__10393),
            .I(N__10384));
    InMux I__2385 (
            .O(N__10392),
            .I(N__10381));
    InMux I__2384 (
            .O(N__10391),
            .I(N__10376));
    InMux I__2383 (
            .O(N__10390),
            .I(N__10376));
    InMux I__2382 (
            .O(N__10389),
            .I(N__10373));
    InMux I__2381 (
            .O(N__10388),
            .I(N__10370));
    InMux I__2380 (
            .O(N__10387),
            .I(N__10367));
    InMux I__2379 (
            .O(N__10384),
            .I(N__10364));
    LocalMux I__2378 (
            .O(N__10381),
            .I(N__10360));
    LocalMux I__2377 (
            .O(N__10376),
            .I(N__10353));
    LocalMux I__2376 (
            .O(N__10373),
            .I(N__10345));
    LocalMux I__2375 (
            .O(N__10370),
            .I(N__10342));
    LocalMux I__2374 (
            .O(N__10367),
            .I(N__10339));
    LocalMux I__2373 (
            .O(N__10364),
            .I(N__10336));
    ClkMux I__2372 (
            .O(N__10363),
            .I(N__10303));
    Glb2LocalMux I__2371 (
            .O(N__10360),
            .I(N__10303));
    ClkMux I__2370 (
            .O(N__10359),
            .I(N__10303));
    ClkMux I__2369 (
            .O(N__10358),
            .I(N__10303));
    ClkMux I__2368 (
            .O(N__10357),
            .I(N__10303));
    ClkMux I__2367 (
            .O(N__10356),
            .I(N__10303));
    Glb2LocalMux I__2366 (
            .O(N__10353),
            .I(N__10303));
    ClkMux I__2365 (
            .O(N__10352),
            .I(N__10303));
    ClkMux I__2364 (
            .O(N__10351),
            .I(N__10303));
    ClkMux I__2363 (
            .O(N__10350),
            .I(N__10303));
    ClkMux I__2362 (
            .O(N__10349),
            .I(N__10303));
    ClkMux I__2361 (
            .O(N__10348),
            .I(N__10303));
    Glb2LocalMux I__2360 (
            .O(N__10345),
            .I(N__10303));
    Glb2LocalMux I__2359 (
            .O(N__10342),
            .I(N__10303));
    Glb2LocalMux I__2358 (
            .O(N__10339),
            .I(N__10303));
    Glb2LocalMux I__2357 (
            .O(N__10336),
            .I(N__10303));
    GlobalMux I__2356 (
            .O(N__10303),
            .I(N__10300));
    gio2CtrlBuf I__2355 (
            .O(N__10300),
            .I(CLK40_IN_c_g));
    IoInMux I__2354 (
            .O(N__10297),
            .I(N__10294));
    LocalMux I__2353 (
            .O(N__10294),
            .I(N__10291));
    Span12Mux_s6_v I__2352 (
            .O(N__10291),
            .I(N__10288));
    Odrv12 I__2351 (
            .O(N__10288),
            .I(GB_BUFFER_CLK40_IN_c_g_THRU_CO));
    InMux I__2350 (
            .O(N__10285),
            .I(N__10280));
    InMux I__2349 (
            .O(N__10284),
            .I(N__10275));
    InMux I__2348 (
            .O(N__10283),
            .I(N__10275));
    LocalMux I__2347 (
            .O(N__10280),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    LocalMux I__2346 (
            .O(N__10275),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    InMux I__2345 (
            .O(N__10270),
            .I(N__10264));
    InMux I__2344 (
            .O(N__10269),
            .I(N__10261));
    InMux I__2343 (
            .O(N__10268),
            .I(N__10256));
    InMux I__2342 (
            .O(N__10267),
            .I(N__10256));
    LocalMux I__2341 (
            .O(N__10264),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__2340 (
            .O(N__10261),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__2339 (
            .O(N__10256),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    InMux I__2338 (
            .O(N__10249),
            .I(N__10245));
    InMux I__2337 (
            .O(N__10248),
            .I(N__10242));
    LocalMux I__2336 (
            .O(N__10245),
            .I(\U409_TRANSFER_ACK.N_3_0 ));
    LocalMux I__2335 (
            .O(N__10242),
            .I(\U409_TRANSFER_ACK.N_3_0 ));
    CascadeMux I__2334 (
            .O(N__10237),
            .I(N__10234));
    InMux I__2333 (
            .O(N__10234),
            .I(N__10231));
    LocalMux I__2332 (
            .O(N__10231),
            .I(N__10226));
    InMux I__2331 (
            .O(N__10230),
            .I(N__10223));
    InMux I__2330 (
            .O(N__10229),
            .I(N__10220));
    Span4Mux_v I__2329 (
            .O(N__10226),
            .I(N__10217));
    LocalMux I__2328 (
            .O(N__10223),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__2327 (
            .O(N__10220),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    Odrv4 I__2326 (
            .O(N__10217),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    CascadeMux I__2325 (
            .O(N__10210),
            .I(\U409_TRANSFER_ACK.N_6_0_cascade_ ));
    InMux I__2324 (
            .O(N__10207),
            .I(N__10204));
    LocalMux I__2323 (
            .O(N__10204),
            .I(N__10198));
    CascadeMux I__2322 (
            .O(N__10203),
            .I(N__10195));
    CascadeMux I__2321 (
            .O(N__10202),
            .I(N__10192));
    CascadeMux I__2320 (
            .O(N__10201),
            .I(N__10188));
    Span4Mux_h I__2319 (
            .O(N__10198),
            .I(N__10185));
    InMux I__2318 (
            .O(N__10195),
            .I(N__10180));
    InMux I__2317 (
            .O(N__10192),
            .I(N__10180));
    InMux I__2316 (
            .O(N__10191),
            .I(N__10175));
    InMux I__2315 (
            .O(N__10188),
            .I(N__10175));
    Odrv4 I__2314 (
            .O(N__10185),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__2313 (
            .O(N__10180),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__2312 (
            .O(N__10175),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    InMux I__2311 (
            .O(N__10168),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__2310 (
            .O(N__10165),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__2309 (
            .O(N__10162),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__2308 (
            .O(N__10159),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    CascadeMux I__2307 (
            .O(N__10156),
            .I(N__10152));
    InMux I__2306 (
            .O(N__10155),
            .I(N__10149));
    InMux I__2305 (
            .O(N__10152),
            .I(N__10146));
    LocalMux I__2304 (
            .O(N__10149),
            .I(N__10143));
    LocalMux I__2303 (
            .O(N__10146),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ));
    Odrv4 I__2302 (
            .O(N__10143),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ));
    CascadeMux I__2301 (
            .O(N__10138),
            .I(N__10135));
    InMux I__2300 (
            .O(N__10135),
            .I(N__10126));
    InMux I__2299 (
            .O(N__10134),
            .I(N__10126));
    InMux I__2298 (
            .O(N__10133),
            .I(N__10123));
    InMux I__2297 (
            .O(N__10132),
            .I(N__10118));
    InMux I__2296 (
            .O(N__10131),
            .I(N__10118));
    LocalMux I__2295 (
            .O(N__10126),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__2294 (
            .O(N__10123),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__2293 (
            .O(N__10118),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    InMux I__2292 (
            .O(N__10111),
            .I(N__10107));
    InMux I__2291 (
            .O(N__10110),
            .I(N__10101));
    LocalMux I__2290 (
            .O(N__10107),
            .I(N__10098));
    InMux I__2289 (
            .O(N__10106),
            .I(N__10093));
    InMux I__2288 (
            .O(N__10105),
            .I(N__10093));
    InMux I__2287 (
            .O(N__10104),
            .I(N__10090));
    LocalMux I__2286 (
            .O(N__10101),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    Odrv4 I__2285 (
            .O(N__10098),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__2284 (
            .O(N__10093),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__2283 (
            .O(N__10090),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    SRMux I__2282 (
            .O(N__10081),
            .I(N__10077));
    SRMux I__2281 (
            .O(N__10080),
            .I(N__10073));
    LocalMux I__2280 (
            .O(N__10077),
            .I(N__10070));
    SRMux I__2279 (
            .O(N__10076),
            .I(N__10067));
    LocalMux I__2278 (
            .O(N__10073),
            .I(N__10064));
    Span4Mux_v I__2277 (
            .O(N__10070),
            .I(N__10059));
    LocalMux I__2276 (
            .O(N__10067),
            .I(N__10059));
    Span4Mux_v I__2275 (
            .O(N__10064),
            .I(N__10056));
    Span4Mux_v I__2274 (
            .O(N__10059),
            .I(N__10053));
    Odrv4 I__2273 (
            .O(N__10056),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv4 I__2272 (
            .O(N__10053),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__2271 (
            .O(N__10048),
            .I(N__10045));
    LocalMux I__2270 (
            .O(N__10045),
            .I(N__10042));
    Span4Mux_v I__2269 (
            .O(N__10042),
            .I(N__10039));
    Odrv4 I__2268 (
            .O(N__10039),
            .I(\U409_ADDRESS_DECODE.un1_Z2_SPACEZ0 ));
    InMux I__2267 (
            .O(N__10036),
            .I(N__10031));
    InMux I__2266 (
            .O(N__10035),
            .I(N__10028));
    CascadeMux I__2265 (
            .O(N__10034),
            .I(N__10025));
    LocalMux I__2264 (
            .O(N__10031),
            .I(N__10022));
    LocalMux I__2263 (
            .O(N__10028),
            .I(N__10019));
    InMux I__2262 (
            .O(N__10025),
            .I(N__10016));
    Span4Mux_h I__2261 (
            .O(N__10022),
            .I(N__10011));
    Span4Mux_v I__2260 (
            .O(N__10019),
            .I(N__10008));
    LocalMux I__2259 (
            .O(N__10016),
            .I(N__10005));
    InMux I__2258 (
            .O(N__10015),
            .I(N__10002));
    InMux I__2257 (
            .O(N__10014),
            .I(N__9999));
    Odrv4 I__2256 (
            .O(N__10011),
            .I(U409_ADDRESS_DECODE_ATA_ROM_EN));
    Odrv4 I__2255 (
            .O(N__10008),
            .I(U409_ADDRESS_DECODE_ATA_ROM_EN));
    Odrv4 I__2254 (
            .O(N__10005),
            .I(U409_ADDRESS_DECODE_ATA_ROM_EN));
    LocalMux I__2253 (
            .O(N__10002),
            .I(U409_ADDRESS_DECODE_ATA_ROM_EN));
    LocalMux I__2252 (
            .O(N__9999),
            .I(U409_ADDRESS_DECODE_ATA_ROM_EN));
    IoInMux I__2251 (
            .O(N__9988),
            .I(N__9985));
    LocalMux I__2250 (
            .O(N__9985),
            .I(N__9982));
    Span12Mux_s10_h I__2249 (
            .O(N__9982),
            .I(N__9979));
    Odrv12 I__2248 (
            .O(N__9979),
            .I(U409_ADDRESS_DECODE_un1_ATA_ENn_i));
    CascadeMux I__2247 (
            .O(N__9976),
            .I(\U409_CIA.CLK_CIA6_4_cascade_ ));
    CascadeMux I__2246 (
            .O(N__9973),
            .I(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ));
    InMux I__2245 (
            .O(N__9970),
            .I(N__9966));
    InMux I__2244 (
            .O(N__9969),
            .I(N__9963));
    LocalMux I__2243 (
            .O(N__9966),
            .I(N__9957));
    LocalMux I__2242 (
            .O(N__9963),
            .I(N__9957));
    InMux I__2241 (
            .O(N__9962),
            .I(N__9954));
    Odrv12 I__2240 (
            .O(N__9957),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__2239 (
            .O(N__9954),
            .I(\U409_CIA.VMAZ0 ));
    InMux I__2238 (
            .O(N__9949),
            .I(N__9944));
    InMux I__2237 (
            .O(N__9948),
            .I(N__9941));
    InMux I__2236 (
            .O(N__9947),
            .I(N__9938));
    LocalMux I__2235 (
            .O(N__9944),
            .I(N__9935));
    LocalMux I__2234 (
            .O(N__9941),
            .I(N__9930));
    LocalMux I__2233 (
            .O(N__9938),
            .I(N__9930));
    Span4Mux_v I__2232 (
            .O(N__9935),
            .I(N__9926));
    Span4Mux_v I__2231 (
            .O(N__9930),
            .I(N__9923));
    InMux I__2230 (
            .O(N__9929),
            .I(N__9920));
    Span4Mux_h I__2229 (
            .O(N__9926),
            .I(N__9916));
    Span4Mux_h I__2228 (
            .O(N__9923),
            .I(N__9911));
    LocalMux I__2227 (
            .O(N__9920),
            .I(N__9911));
    InMux I__2226 (
            .O(N__9919),
            .I(N__9908));
    Odrv4 I__2225 (
            .O(N__9916),
            .I(AUTOCONFIG_SPACE));
    Odrv4 I__2224 (
            .O(N__9911),
            .I(AUTOCONFIG_SPACE));
    LocalMux I__2223 (
            .O(N__9908),
            .I(AUTOCONFIG_SPACE));
    InMux I__2222 (
            .O(N__9901),
            .I(N__9898));
    LocalMux I__2221 (
            .O(N__9898),
            .I(N__9893));
    InMux I__2220 (
            .O(N__9897),
            .I(N__9890));
    InMux I__2219 (
            .O(N__9896),
            .I(N__9887));
    Span4Mux_v I__2218 (
            .O(N__9893),
            .I(N__9884));
    LocalMux I__2217 (
            .O(N__9890),
            .I(N__9879));
    LocalMux I__2216 (
            .O(N__9887),
            .I(N__9879));
    Odrv4 I__2215 (
            .O(N__9884),
            .I(CIA_SPACE));
    Odrv12 I__2214 (
            .O(N__9879),
            .I(CIA_SPACE));
    IoInMux I__2213 (
            .O(N__9874),
            .I(N__9870));
    IoInMux I__2212 (
            .O(N__9873),
            .I(N__9867));
    LocalMux I__2211 (
            .O(N__9870),
            .I(N__9862));
    LocalMux I__2210 (
            .O(N__9867),
            .I(N__9862));
    IoSpan4Mux I__2209 (
            .O(N__9862),
            .I(N__9859));
    Span4Mux_s2_v I__2208 (
            .O(N__9859),
            .I(N__9856));
    Span4Mux_v I__2207 (
            .O(N__9856),
            .I(N__9852));
    InMux I__2206 (
            .O(N__9855),
            .I(N__9849));
    Sp12to4 I__2205 (
            .O(N__9852),
            .I(N__9845));
    LocalMux I__2204 (
            .O(N__9849),
            .I(N__9842));
    CascadeMux I__2203 (
            .O(N__9848),
            .I(N__9839));
    Span12Mux_v I__2202 (
            .O(N__9845),
            .I(N__9836));
    Span4Mux_v I__2201 (
            .O(N__9842),
            .I(N__9833));
    InMux I__2200 (
            .O(N__9839),
            .I(N__9830));
    Odrv12 I__2199 (
            .O(N__9836),
            .I(TACK_EN));
    Odrv4 I__2198 (
            .O(N__9833),
            .I(TACK_EN));
    LocalMux I__2197 (
            .O(N__9830),
            .I(TACK_EN));
    IoInMux I__2196 (
            .O(N__9823),
            .I(N__9820));
    LocalMux I__2195 (
            .O(N__9820),
            .I(N__9817));
    Span4Mux_s3_v I__2194 (
            .O(N__9817),
            .I(N__9814));
    Span4Mux_h I__2193 (
            .O(N__9814),
            .I(N__9811));
    Span4Mux_h I__2192 (
            .O(N__9811),
            .I(N__9808));
    Sp12to4 I__2191 (
            .O(N__9808),
            .I(N__9805));
    Span12Mux_v I__2190 (
            .O(N__9805),
            .I(N__9802));
    Odrv12 I__2189 (
            .O(N__9802),
            .I(TCIn_1_i));
    IoInMux I__2188 (
            .O(N__9799),
            .I(N__9795));
    IoInMux I__2187 (
            .O(N__9798),
            .I(N__9792));
    LocalMux I__2186 (
            .O(N__9795),
            .I(N__9787));
    LocalMux I__2185 (
            .O(N__9792),
            .I(N__9787));
    IoSpan4Mux I__2184 (
            .O(N__9787),
            .I(N__9782));
    IoInMux I__2183 (
            .O(N__9786),
            .I(N__9779));
    IoInMux I__2182 (
            .O(N__9785),
            .I(N__9776));
    IoSpan4Mux I__2181 (
            .O(N__9782),
            .I(N__9773));
    LocalMux I__2180 (
            .O(N__9779),
            .I(N__9768));
    LocalMux I__2179 (
            .O(N__9776),
            .I(N__9768));
    IoSpan4Mux I__2178 (
            .O(N__9773),
            .I(N__9763));
    IoSpan4Mux I__2177 (
            .O(N__9768),
            .I(N__9763));
    Span4Mux_s0_h I__2176 (
            .O(N__9763),
            .I(N__9760));
    Span4Mux_h I__2175 (
            .O(N__9760),
            .I(N__9756));
    IoInMux I__2174 (
            .O(N__9759),
            .I(N__9753));
    Span4Mux_h I__2173 (
            .O(N__9756),
            .I(N__9750));
    LocalMux I__2172 (
            .O(N__9753),
            .I(N__9747));
    Span4Mux_h I__2171 (
            .O(N__9750),
            .I(N__9742));
    Span4Mux_s2_v I__2170 (
            .O(N__9747),
            .I(N__9742));
    Span4Mux_v I__2169 (
            .O(N__9742),
            .I(N__9739));
    Odrv4 I__2168 (
            .O(N__9739),
            .I(CONSTANT_ONE_NET));
    SRMux I__2167 (
            .O(N__9736),
            .I(N__9703));
    SRMux I__2166 (
            .O(N__9735),
            .I(N__9703));
    SRMux I__2165 (
            .O(N__9734),
            .I(N__9703));
    SRMux I__2164 (
            .O(N__9733),
            .I(N__9703));
    SRMux I__2163 (
            .O(N__9732),
            .I(N__9703));
    SRMux I__2162 (
            .O(N__9731),
            .I(N__9703));
    SRMux I__2161 (
            .O(N__9730),
            .I(N__9703));
    SRMux I__2160 (
            .O(N__9729),
            .I(N__9703));
    SRMux I__2159 (
            .O(N__9728),
            .I(N__9703));
    SRMux I__2158 (
            .O(N__9727),
            .I(N__9703));
    SRMux I__2157 (
            .O(N__9726),
            .I(N__9703));
    GlobalMux I__2156 (
            .O(N__9703),
            .I(N__9700));
    gio2CtrlBuf I__2155 (
            .O(N__9700),
            .I(RESETn_c_i_g));
    CascadeMux I__2154 (
            .O(N__9697),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_ ));
    InMux I__2153 (
            .O(N__9694),
            .I(N__9691));
    LocalMux I__2152 (
            .O(N__9691),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ));
    InMux I__2151 (
            .O(N__9688),
            .I(N__9684));
    InMux I__2150 (
            .O(N__9687),
            .I(N__9681));
    LocalMux I__2149 (
            .O(N__9684),
            .I(\U409_TRANSFER_ACK.N_17_mux ));
    LocalMux I__2148 (
            .O(N__9681),
            .I(\U409_TRANSFER_ACK.N_17_mux ));
    InMux I__2147 (
            .O(N__9676),
            .I(N__9670));
    InMux I__2146 (
            .O(N__9675),
            .I(N__9665));
    InMux I__2145 (
            .O(N__9674),
            .I(N__9665));
    InMux I__2144 (
            .O(N__9673),
            .I(N__9662));
    LocalMux I__2143 (
            .O(N__9670),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__2142 (
            .O(N__9665),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__2141 (
            .O(N__9662),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    InMux I__2140 (
            .O(N__9655),
            .I(N__9649));
    CascadeMux I__2139 (
            .O(N__9654),
            .I(N__9646));
    InMux I__2138 (
            .O(N__9653),
            .I(N__9641));
    InMux I__2137 (
            .O(N__9652),
            .I(N__9641));
    LocalMux I__2136 (
            .O(N__9649),
            .I(N__9638));
    InMux I__2135 (
            .O(N__9646),
            .I(N__9635));
    LocalMux I__2134 (
            .O(N__9641),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    Odrv4 I__2133 (
            .O(N__9638),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__2132 (
            .O(N__9635),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    InMux I__2131 (
            .O(N__9628),
            .I(N__9624));
    InMux I__2130 (
            .O(N__9627),
            .I(N__9621));
    LocalMux I__2129 (
            .O(N__9624),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    LocalMux I__2128 (
            .O(N__9621),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    CascadeMux I__2127 (
            .O(N__9616),
            .I(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ));
    IoInMux I__2126 (
            .O(N__9613),
            .I(N__9609));
    IoInMux I__2125 (
            .O(N__9612),
            .I(N__9606));
    LocalMux I__2124 (
            .O(N__9609),
            .I(N__9601));
    LocalMux I__2123 (
            .O(N__9606),
            .I(N__9601));
    IoSpan4Mux I__2122 (
            .O(N__9601),
            .I(N__9597));
    IoInMux I__2121 (
            .O(N__9600),
            .I(N__9594));
    Span4Mux_s3_v I__2120 (
            .O(N__9597),
            .I(N__9591));
    LocalMux I__2119 (
            .O(N__9594),
            .I(N__9588));
    Span4Mux_v I__2118 (
            .O(N__9591),
            .I(N__9583));
    Span4Mux_s3_v I__2117 (
            .O(N__9588),
            .I(N__9583));
    Sp12to4 I__2116 (
            .O(N__9583),
            .I(N__9580));
    Span12Mux_h I__2115 (
            .O(N__9580),
            .I(N__9577));
    Span12Mux_v I__2114 (
            .O(N__9577),
            .I(N__9572));
    InMux I__2113 (
            .O(N__9576),
            .I(N__9567));
    InMux I__2112 (
            .O(N__9575),
            .I(N__9567));
    Odrv12 I__2111 (
            .O(N__9572),
            .I(TACK_OUTn));
    LocalMux I__2110 (
            .O(N__9567),
            .I(TACK_OUTn));
    InMux I__2109 (
            .O(N__9562),
            .I(N__9558));
    InMux I__2108 (
            .O(N__9561),
            .I(N__9555));
    LocalMux I__2107 (
            .O(N__9558),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    LocalMux I__2106 (
            .O(N__9555),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    InMux I__2105 (
            .O(N__9550),
            .I(N__9545));
    InMux I__2104 (
            .O(N__9549),
            .I(N__9540));
    InMux I__2103 (
            .O(N__9548),
            .I(N__9540));
    LocalMux I__2102 (
            .O(N__9545),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__2101 (
            .O(N__9540),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__2100 (
            .O(N__9535),
            .I(N__9532));
    LocalMux I__2099 (
            .O(N__9532),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    InMux I__2098 (
            .O(N__9529),
            .I(N__9524));
    InMux I__2097 (
            .O(N__9528),
            .I(N__9521));
    InMux I__2096 (
            .O(N__9527),
            .I(N__9518));
    LocalMux I__2095 (
            .O(N__9524),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    LocalMux I__2094 (
            .O(N__9521),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    LocalMux I__2093 (
            .O(N__9518),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    InMux I__2092 (
            .O(N__9511),
            .I(N__9507));
    InMux I__2091 (
            .O(N__9510),
            .I(N__9504));
    LocalMux I__2090 (
            .O(N__9507),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    LocalMux I__2089 (
            .O(N__9504),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    InMux I__2088 (
            .O(N__9499),
            .I(N__9494));
    InMux I__2087 (
            .O(N__9498),
            .I(N__9489));
    InMux I__2086 (
            .O(N__9497),
            .I(N__9485));
    LocalMux I__2085 (
            .O(N__9494),
            .I(N__9482));
    InMux I__2084 (
            .O(N__9493),
            .I(N__9479));
    InMux I__2083 (
            .O(N__9492),
            .I(N__9476));
    LocalMux I__2082 (
            .O(N__9489),
            .I(N__9472));
    InMux I__2081 (
            .O(N__9488),
            .I(N__9469));
    LocalMux I__2080 (
            .O(N__9485),
            .I(N__9466));
    Span4Mux_v I__2079 (
            .O(N__9482),
            .I(N__9461));
    LocalMux I__2078 (
            .O(N__9479),
            .I(N__9461));
    LocalMux I__2077 (
            .O(N__9476),
            .I(N__9458));
    InMux I__2076 (
            .O(N__9475),
            .I(N__9455));
    Span4Mux_v I__2075 (
            .O(N__9472),
            .I(N__9450));
    LocalMux I__2074 (
            .O(N__9469),
            .I(N__9450));
    Span4Mux_v I__2073 (
            .O(N__9466),
            .I(N__9447));
    Span4Mux_h I__2072 (
            .O(N__9461),
            .I(N__9440));
    Span4Mux_v I__2071 (
            .O(N__9458),
            .I(N__9440));
    LocalMux I__2070 (
            .O(N__9455),
            .I(N__9440));
    Span4Mux_v I__2069 (
            .O(N__9450),
            .I(N__9437));
    Span4Mux_h I__2068 (
            .O(N__9447),
            .I(N__9432));
    Span4Mux_v I__2067 (
            .O(N__9440),
            .I(N__9432));
    Sp12to4 I__2066 (
            .O(N__9437),
            .I(N__9427));
    Sp12to4 I__2065 (
            .O(N__9432),
            .I(N__9427));
    Span12Mux_h I__2064 (
            .O(N__9427),
            .I(N__9424));
    Span12Mux_v I__2063 (
            .O(N__9424),
            .I(N__9421));
    Odrv12 I__2062 (
            .O(N__9421),
            .I(TSn_c));
    InMux I__2061 (
            .O(N__9418),
            .I(N__9401));
    InMux I__2060 (
            .O(N__9417),
            .I(N__9401));
    InMux I__2059 (
            .O(N__9416),
            .I(N__9401));
    InMux I__2058 (
            .O(N__9415),
            .I(N__9401));
    InMux I__2057 (
            .O(N__9414),
            .I(N__9401));
    InMux I__2056 (
            .O(N__9413),
            .I(N__9396));
    InMux I__2055 (
            .O(N__9412),
            .I(N__9396));
    LocalMux I__2054 (
            .O(N__9401),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__2053 (
            .O(N__9396),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    InMux I__2052 (
            .O(N__9391),
            .I(N__9388));
    LocalMux I__2051 (
            .O(N__9388),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    CascadeMux I__2050 (
            .O(N__9385),
            .I(N__9382));
    InMux I__2049 (
            .O(N__9382),
            .I(N__9379));
    LocalMux I__2048 (
            .O(N__9379),
            .I(N__9376));
    Span4Mux_h I__2047 (
            .O(N__9376),
            .I(N__9373));
    Sp12to4 I__2046 (
            .O(N__9373),
            .I(N__9370));
    Span12Mux_h I__2045 (
            .O(N__9370),
            .I(N__9367));
    Span12Mux_v I__2044 (
            .O(N__9367),
            .I(N__9364));
    Odrv12 I__2043 (
            .O(N__9364),
            .I(TACKn_in));
    CascadeMux I__2042 (
            .O(N__9361),
            .I(N__9358));
    InMux I__2041 (
            .O(N__9358),
            .I(N__9355));
    LocalMux I__2040 (
            .O(N__9355),
            .I(N__9351));
    InMux I__2039 (
            .O(N__9354),
            .I(N__9348));
    Span4Mux_v I__2038 (
            .O(N__9351),
            .I(N__9343));
    LocalMux I__2037 (
            .O(N__9348),
            .I(N__9343));
    Odrv4 I__2036 (
            .O(N__9343),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn));
    IoInMux I__2035 (
            .O(N__9340),
            .I(N__9337));
    LocalMux I__2034 (
            .O(N__9337),
            .I(N__9334));
    Span12Mux_s1_v I__2033 (
            .O(N__9334),
            .I(N__9331));
    Span12Mux_h I__2032 (
            .O(N__9331),
            .I(N__9328));
    Odrv12 I__2031 (
            .O(N__9328),
            .I(BUFENn_c));
    InMux I__2030 (
            .O(N__9325),
            .I(N__9319));
    InMux I__2029 (
            .O(N__9324),
            .I(N__9319));
    LocalMux I__2028 (
            .O(N__9319),
            .I(N__9316));
    Span4Mux_v I__2027 (
            .O(N__9316),
            .I(N__9312));
    InMux I__2026 (
            .O(N__9315),
            .I(N__9309));
    Odrv4 I__2025 (
            .O(N__9312),
            .I(U409_ADDRESS_DECODE_un2_REGSPACEn_0));
    LocalMux I__2024 (
            .O(N__9309),
            .I(U409_ADDRESS_DECODE_un2_REGSPACEn_0));
    InMux I__2023 (
            .O(N__9304),
            .I(N__9298));
    InMux I__2022 (
            .O(N__9303),
            .I(N__9298));
    LocalMux I__2021 (
            .O(N__9298),
            .I(N__9292));
    InMux I__2020 (
            .O(N__9297),
            .I(N__9286));
    InMux I__2019 (
            .O(N__9296),
            .I(N__9286));
    InMux I__2018 (
            .O(N__9295),
            .I(N__9283));
    Span4Mux_h I__2017 (
            .O(N__9292),
            .I(N__9280));
    InMux I__2016 (
            .O(N__9291),
            .I(N__9277));
    LocalMux I__2015 (
            .O(N__9286),
            .I(N__9271));
    LocalMux I__2014 (
            .O(N__9283),
            .I(N__9271));
    Span4Mux_v I__2013 (
            .O(N__9280),
            .I(N__9266));
    LocalMux I__2012 (
            .O(N__9277),
            .I(N__9266));
    InMux I__2011 (
            .O(N__9276),
            .I(N__9263));
    Span4Mux_v I__2010 (
            .O(N__9271),
            .I(N__9260));
    Span4Mux_h I__2009 (
            .O(N__9266),
            .I(N__9257));
    LocalMux I__2008 (
            .O(N__9263),
            .I(N__9254));
    Sp12to4 I__2007 (
            .O(N__9260),
            .I(N__9251));
    Span4Mux_v I__2006 (
            .O(N__9257),
            .I(N__9248));
    Span4Mux_v I__2005 (
            .O(N__9254),
            .I(N__9245));
    Odrv12 I__2004 (
            .O(N__9251),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    Odrv4 I__2003 (
            .O(N__9248),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    Odrv4 I__2002 (
            .O(N__9245),
            .I(U409_ADDRESS_DECODE_Z2_SPACE));
    IoInMux I__2001 (
            .O(N__9238),
            .I(N__9235));
    LocalMux I__2000 (
            .O(N__9235),
            .I(N__9232));
    IoSpan4Mux I__1999 (
            .O(N__9232),
            .I(N__9229));
    Sp12to4 I__1998 (
            .O(N__9229),
            .I(N__9226));
    Span12Mux_v I__1997 (
            .O(N__9226),
            .I(N__9223));
    Odrv12 I__1996 (
            .O(N__9223),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn_i));
    CascadeMux I__1995 (
            .O(N__9220),
            .I(CIA_ENABLE_cascade_));
    InMux I__1994 (
            .O(N__9217),
            .I(N__9214));
    LocalMux I__1993 (
            .O(N__9214),
            .I(N__9211));
    Span4Mux_v I__1992 (
            .O(N__9211),
            .I(N__9208));
    Sp12to4 I__1991 (
            .O(N__9208),
            .I(N__9205));
    Span12Mux_h I__1990 (
            .O(N__9205),
            .I(N__9202));
    Odrv12 I__1989 (
            .O(N__9202),
            .I(A_c_12));
    IoInMux I__1988 (
            .O(N__9199),
            .I(N__9196));
    LocalMux I__1987 (
            .O(N__9196),
            .I(N__9193));
    Span4Mux_s1_h I__1986 (
            .O(N__9193),
            .I(N__9190));
    Sp12to4 I__1985 (
            .O(N__9190),
            .I(N__9187));
    Span12Mux_s8_v I__1984 (
            .O(N__9187),
            .I(N__9184));
    Span12Mux_h I__1983 (
            .O(N__9184),
            .I(N__9181));
    Odrv12 I__1982 (
            .O(N__9181),
            .I(U409_ADDRESS_DECODE_un1_CIACS0n_i));
    InMux I__1981 (
            .O(N__9178),
            .I(N__9175));
    LocalMux I__1980 (
            .O(N__9175),
            .I(CIA_ENABLE));
    InMux I__1979 (
            .O(N__9172),
            .I(N__9169));
    LocalMux I__1978 (
            .O(N__9169),
            .I(N__9166));
    Span4Mux_v I__1977 (
            .O(N__9166),
            .I(N__9163));
    Sp12to4 I__1976 (
            .O(N__9163),
            .I(N__9160));
    Span12Mux_h I__1975 (
            .O(N__9160),
            .I(N__9157));
    Odrv12 I__1974 (
            .O(N__9157),
            .I(A_c_13));
    IoInMux I__1973 (
            .O(N__9154),
            .I(N__9151));
    LocalMux I__1972 (
            .O(N__9151),
            .I(N__9148));
    IoSpan4Mux I__1971 (
            .O(N__9148),
            .I(N__9145));
    IoSpan4Mux I__1970 (
            .O(N__9145),
            .I(N__9142));
    Sp12to4 I__1969 (
            .O(N__9142),
            .I(N__9139));
    Span12Mux_s7_h I__1968 (
            .O(N__9139),
            .I(N__9136));
    Odrv12 I__1967 (
            .O(N__9136),
            .I(U409_ADDRESS_DECODE_un1_CIACS1n_i));
    CascadeMux I__1966 (
            .O(N__9133),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ));
    CascadeMux I__1965 (
            .O(N__9130),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    CascadeMux I__1964 (
            .O(N__9127),
            .I(N__9121));
    InMux I__1963 (
            .O(N__9126),
            .I(N__9116));
    InMux I__1962 (
            .O(N__9125),
            .I(N__9116));
    InMux I__1961 (
            .O(N__9124),
            .I(N__9111));
    InMux I__1960 (
            .O(N__9121),
            .I(N__9111));
    LocalMux I__1959 (
            .O(N__9116),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__1958 (
            .O(N__9111),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    InMux I__1957 (
            .O(N__9106),
            .I(N__9100));
    InMux I__1956 (
            .O(N__9105),
            .I(N__9100));
    LocalMux I__1955 (
            .O(N__9100),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    CascadeMux I__1954 (
            .O(N__9097),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ));
    InMux I__1953 (
            .O(N__9094),
            .I(N__9079));
    InMux I__1952 (
            .O(N__9093),
            .I(N__9079));
    InMux I__1951 (
            .O(N__9092),
            .I(N__9079));
    InMux I__1950 (
            .O(N__9091),
            .I(N__9079));
    InMux I__1949 (
            .O(N__9090),
            .I(N__9079));
    LocalMux I__1948 (
            .O(N__9079),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    CascadeMux I__1947 (
            .O(N__9076),
            .I(N__9071));
    CascadeMux I__1946 (
            .O(N__9075),
            .I(N__9068));
    CascadeMux I__1945 (
            .O(N__9074),
            .I(N__9065));
    InMux I__1944 (
            .O(N__9071),
            .I(N__9055));
    InMux I__1943 (
            .O(N__9068),
            .I(N__9055));
    InMux I__1942 (
            .O(N__9065),
            .I(N__9055));
    InMux I__1941 (
            .O(N__9064),
            .I(N__9055));
    LocalMux I__1940 (
            .O(N__9055),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    CascadeMux I__1939 (
            .O(N__9052),
            .I(N__9047));
    InMux I__1938 (
            .O(N__9051),
            .I(N__9041));
    InMux I__1937 (
            .O(N__9050),
            .I(N__9041));
    InMux I__1936 (
            .O(N__9047),
            .I(N__9038));
    InMux I__1935 (
            .O(N__9046),
            .I(N__9035));
    LocalMux I__1934 (
            .O(N__9041),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1933 (
            .O(N__9038),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1932 (
            .O(N__9035),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__1931 (
            .O(N__9028),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_ ));
    InMux I__1930 (
            .O(N__9025),
            .I(N__9019));
    InMux I__1929 (
            .O(N__9024),
            .I(N__9016));
    InMux I__1928 (
            .O(N__9023),
            .I(N__9011));
    InMux I__1927 (
            .O(N__9022),
            .I(N__9011));
    LocalMux I__1926 (
            .O(N__9019),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__1925 (
            .O(N__9016),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__1924 (
            .O(N__9011),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    InMux I__1923 (
            .O(N__9004),
            .I(N__8998));
    InMux I__1922 (
            .O(N__9003),
            .I(N__8998));
    LocalMux I__1921 (
            .O(N__8998),
            .I(N__8995));
    Odrv4 I__1920 (
            .O(N__8995),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    CascadeMux I__1919 (
            .O(N__8992),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ));
    InMux I__1918 (
            .O(N__8989),
            .I(N__8982));
    InMux I__1917 (
            .O(N__8988),
            .I(N__8982));
    InMux I__1916 (
            .O(N__8987),
            .I(N__8979));
    LocalMux I__1915 (
            .O(N__8982),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__1914 (
            .O(N__8979),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    CascadeMux I__1913 (
            .O(N__8974),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_ ));
    InMux I__1912 (
            .O(N__8971),
            .I(N__8968));
    LocalMux I__1911 (
            .O(N__8968),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_2 ));
    InMux I__1910 (
            .O(N__8965),
            .I(N__8959));
    InMux I__1909 (
            .O(N__8964),
            .I(N__8959));
    LocalMux I__1908 (
            .O(N__8959),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    InMux I__1907 (
            .O(N__8956),
            .I(N__8953));
    LocalMux I__1906 (
            .O(N__8953),
            .I(N__8949));
    InMux I__1905 (
            .O(N__8952),
            .I(N__8946));
    Span4Mux_v I__1904 (
            .O(N__8949),
            .I(N__8941));
    LocalMux I__1903 (
            .O(N__8946),
            .I(N__8941));
    Span4Mux_v I__1902 (
            .O(N__8941),
            .I(N__8937));
    InMux I__1901 (
            .O(N__8940),
            .I(N__8934));
    Odrv4 I__1900 (
            .O(N__8937),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn));
    LocalMux I__1899 (
            .O(N__8934),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn));
    CascadeMux I__1898 (
            .O(N__8929),
            .I(N__8926));
    InMux I__1897 (
            .O(N__8926),
            .I(N__8922));
    InMux I__1896 (
            .O(N__8925),
            .I(N__8919));
    LocalMux I__1895 (
            .O(N__8922),
            .I(N__8914));
    LocalMux I__1894 (
            .O(N__8919),
            .I(N__8914));
    Span4Mux_h I__1893 (
            .O(N__8914),
            .I(N__8911));
    Span4Mux_v I__1892 (
            .O(N__8911),
            .I(N__8908));
    Span4Mux_v I__1891 (
            .O(N__8908),
            .I(N__8905));
    Odrv4 I__1890 (
            .O(N__8905),
            .I(AUTOVECTOR));
    InMux I__1889 (
            .O(N__8902),
            .I(N__8899));
    LocalMux I__1888 (
            .O(N__8899),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0 ));
    InMux I__1887 (
            .O(N__8896),
            .I(N__8893));
    LocalMux I__1886 (
            .O(N__8893),
            .I(N__8890));
    Span4Mux_h I__1885 (
            .O(N__8890),
            .I(N__8887));
    Span4Mux_h I__1884 (
            .O(N__8887),
            .I(N__8884));
    Odrv4 I__1883 (
            .O(N__8884),
            .I(AC_TACK));
    CascadeMux I__1882 (
            .O(N__8881),
            .I(N__8878));
    InMux I__1881 (
            .O(N__8878),
            .I(N__8874));
    InMux I__1880 (
            .O(N__8877),
            .I(N__8871));
    LocalMux I__1879 (
            .O(N__8874),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    LocalMux I__1878 (
            .O(N__8871),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    CascadeMux I__1877 (
            .O(N__8866),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ));
    CascadeMux I__1876 (
            .O(N__8863),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ));
    CascadeMux I__1875 (
            .O(N__8860),
            .I(N__8856));
    InMux I__1874 (
            .O(N__8859),
            .I(N__8853));
    InMux I__1873 (
            .O(N__8856),
            .I(N__8850));
    LocalMux I__1872 (
            .O(N__8853),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__1871 (
            .O(N__8850),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    InMux I__1870 (
            .O(N__8845),
            .I(N__8842));
    LocalMux I__1869 (
            .O(N__8842),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3 ));
    InMux I__1868 (
            .O(N__8839),
            .I(N__8836));
    LocalMux I__1867 (
            .O(N__8836),
            .I(\U409_TRANSFER_ACK.ROMENn_1_sqmuxa_d ));
    IoInMux I__1866 (
            .O(N__8833),
            .I(N__8830));
    LocalMux I__1865 (
            .O(N__8830),
            .I(N__8827));
    IoSpan4Mux I__1864 (
            .O(N__8827),
            .I(N__8824));
    Sp12to4 I__1863 (
            .O(N__8824),
            .I(N__8821));
    Span12Mux_s6_v I__1862 (
            .O(N__8821),
            .I(N__8818));
    Span12Mux_v I__1861 (
            .O(N__8818),
            .I(N__8814));
    InMux I__1860 (
            .O(N__8817),
            .I(N__8811));
    Odrv12 I__1859 (
            .O(N__8814),
            .I(ROMENn_c));
    LocalMux I__1858 (
            .O(N__8811),
            .I(ROMENn_c));
    CascadeMux I__1857 (
            .O(N__8806),
            .I(N__8803));
    InMux I__1856 (
            .O(N__8803),
            .I(N__8799));
    InMux I__1855 (
            .O(N__8802),
            .I(N__8796));
    LocalMux I__1854 (
            .O(N__8799),
            .I(N__8790));
    LocalMux I__1853 (
            .O(N__8796),
            .I(N__8790));
    InMux I__1852 (
            .O(N__8795),
            .I(N__8783));
    Span4Mux_h I__1851 (
            .O(N__8790),
            .I(N__8780));
    InMux I__1850 (
            .O(N__8789),
            .I(N__8777));
    InMux I__1849 (
            .O(N__8788),
            .I(N__8770));
    InMux I__1848 (
            .O(N__8787),
            .I(N__8770));
    InMux I__1847 (
            .O(N__8786),
            .I(N__8770));
    LocalMux I__1846 (
            .O(N__8783),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    Odrv4 I__1845 (
            .O(N__8780),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1844 (
            .O(N__8777),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1843 (
            .O(N__8770),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    InMux I__1842 (
            .O(N__8761),
            .I(N__8758));
    LocalMux I__1841 (
            .O(N__8758),
            .I(N__8755));
    Span4Mux_h I__1840 (
            .O(N__8755),
            .I(N__8746));
    InMux I__1839 (
            .O(N__8754),
            .I(N__8743));
    InMux I__1838 (
            .O(N__8753),
            .I(N__8740));
    InMux I__1837 (
            .O(N__8752),
            .I(N__8737));
    InMux I__1836 (
            .O(N__8751),
            .I(N__8730));
    InMux I__1835 (
            .O(N__8750),
            .I(N__8730));
    InMux I__1834 (
            .O(N__8749),
            .I(N__8730));
    Odrv4 I__1833 (
            .O(N__8746),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1832 (
            .O(N__8743),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1831 (
            .O(N__8740),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1830 (
            .O(N__8737),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1829 (
            .O(N__8730),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    CascadeMux I__1828 (
            .O(N__8719),
            .I(N__8716));
    InMux I__1827 (
            .O(N__8716),
            .I(N__8713));
    LocalMux I__1826 (
            .O(N__8713),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20_2 ));
    InMux I__1825 (
            .O(N__8710),
            .I(N__8706));
    InMux I__1824 (
            .O(N__8709),
            .I(N__8703));
    LocalMux I__1823 (
            .O(N__8706),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__1822 (
            .O(N__8703),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__1821 (
            .O(N__8698),
            .I(N__8695));
    LocalMux I__1820 (
            .O(N__8695),
            .I(N__8692));
    Odrv4 I__1819 (
            .O(N__8692),
            .I(\U409_TRANSFER_ACK.G_14_0_o7_6 ));
    CascadeMux I__1818 (
            .O(N__8689),
            .I(\U409_TRANSFER_ACK.G_14_0_4_cascade_ ));
    InMux I__1817 (
            .O(N__8686),
            .I(N__8683));
    LocalMux I__1816 (
            .O(N__8683),
            .I(\U409_TRANSFER_ACK.g0_0_0_o6_4 ));
    CascadeMux I__1815 (
            .O(N__8680),
            .I(N__8677));
    InMux I__1814 (
            .O(N__8677),
            .I(N__8671));
    InMux I__1813 (
            .O(N__8676),
            .I(N__8671));
    LocalMux I__1812 (
            .O(N__8671),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER15_out ));
    CascadeMux I__1811 (
            .O(N__8668),
            .I(N__8664));
    CascadeMux I__1810 (
            .O(N__8667),
            .I(N__8658));
    InMux I__1809 (
            .O(N__8664),
            .I(N__8653));
    InMux I__1808 (
            .O(N__8663),
            .I(N__8650));
    InMux I__1807 (
            .O(N__8662),
            .I(N__8641));
    InMux I__1806 (
            .O(N__8661),
            .I(N__8641));
    InMux I__1805 (
            .O(N__8658),
            .I(N__8641));
    InMux I__1804 (
            .O(N__8657),
            .I(N__8641));
    InMux I__1803 (
            .O(N__8656),
            .I(N__8638));
    LocalMux I__1802 (
            .O(N__8653),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1801 (
            .O(N__8650),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1800 (
            .O(N__8641),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1799 (
            .O(N__8638),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    CascadeMux I__1798 (
            .O(N__8629),
            .I(N__8620));
    CascadeMux I__1797 (
            .O(N__8628),
            .I(N__8617));
    InMux I__1796 (
            .O(N__8627),
            .I(N__8614));
    InMux I__1795 (
            .O(N__8626),
            .I(N__8611));
    InMux I__1794 (
            .O(N__8625),
            .I(N__8602));
    InMux I__1793 (
            .O(N__8624),
            .I(N__8602));
    InMux I__1792 (
            .O(N__8623),
            .I(N__8602));
    InMux I__1791 (
            .O(N__8620),
            .I(N__8602));
    InMux I__1790 (
            .O(N__8617),
            .I(N__8599));
    LocalMux I__1789 (
            .O(N__8614),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1788 (
            .O(N__8611),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1787 (
            .O(N__8602),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1786 (
            .O(N__8599),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__1785 (
            .O(N__8590),
            .I(N__8585));
    InMux I__1784 (
            .O(N__8589),
            .I(N__8580));
    InMux I__1783 (
            .O(N__8588),
            .I(N__8580));
    LocalMux I__1782 (
            .O(N__8585),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ));
    LocalMux I__1781 (
            .O(N__8580),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ));
    CascadeMux I__1780 (
            .O(N__8575),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0_cascade_ ));
    InMux I__1779 (
            .O(N__8572),
            .I(N__8567));
    InMux I__1778 (
            .O(N__8571),
            .I(N__8564));
    InMux I__1777 (
            .O(N__8570),
            .I(N__8561));
    LocalMux I__1776 (
            .O(N__8567),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ));
    LocalMux I__1775 (
            .O(N__8564),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ));
    LocalMux I__1774 (
            .O(N__8561),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ));
    InMux I__1773 (
            .O(N__8554),
            .I(N__8551));
    LocalMux I__1772 (
            .O(N__8551),
            .I(\U409_TRANSFER_ACK.ROMENn_1_sqmuxa_0_c ));
    InMux I__1771 (
            .O(N__8548),
            .I(N__8539));
    InMux I__1770 (
            .O(N__8547),
            .I(N__8533));
    InMux I__1769 (
            .O(N__8546),
            .I(N__8528));
    InMux I__1768 (
            .O(N__8545),
            .I(N__8523));
    InMux I__1767 (
            .O(N__8544),
            .I(N__8523));
    InMux I__1766 (
            .O(N__8543),
            .I(N__8517));
    InMux I__1765 (
            .O(N__8542),
            .I(N__8517));
    LocalMux I__1764 (
            .O(N__8539),
            .I(N__8514));
    InMux I__1763 (
            .O(N__8538),
            .I(N__8509));
    InMux I__1762 (
            .O(N__8537),
            .I(N__8509));
    InMux I__1761 (
            .O(N__8536),
            .I(N__8506));
    LocalMux I__1760 (
            .O(N__8533),
            .I(N__8502));
    InMux I__1759 (
            .O(N__8532),
            .I(N__8497));
    InMux I__1758 (
            .O(N__8531),
            .I(N__8497));
    LocalMux I__1757 (
            .O(N__8528),
            .I(N__8492));
    LocalMux I__1756 (
            .O(N__8523),
            .I(N__8492));
    InMux I__1755 (
            .O(N__8522),
            .I(N__8489));
    LocalMux I__1754 (
            .O(N__8517),
            .I(N__8485));
    Span4Mux_h I__1753 (
            .O(N__8514),
            .I(N__8478));
    LocalMux I__1752 (
            .O(N__8509),
            .I(N__8478));
    LocalMux I__1751 (
            .O(N__8506),
            .I(N__8478));
    InMux I__1750 (
            .O(N__8505),
            .I(N__8475));
    Span4Mux_v I__1749 (
            .O(N__8502),
            .I(N__8466));
    LocalMux I__1748 (
            .O(N__8497),
            .I(N__8466));
    Span4Mux_v I__1747 (
            .O(N__8492),
            .I(N__8466));
    LocalMux I__1746 (
            .O(N__8489),
            .I(N__8466));
    InMux I__1745 (
            .O(N__8488),
            .I(N__8463));
    Span4Mux_v I__1744 (
            .O(N__8485),
            .I(N__8460));
    Span4Mux_v I__1743 (
            .O(N__8478),
            .I(N__8455));
    LocalMux I__1742 (
            .O(N__8475),
            .I(N__8455));
    Span4Mux_h I__1741 (
            .O(N__8466),
            .I(N__8450));
    LocalMux I__1740 (
            .O(N__8463),
            .I(N__8450));
    Span4Mux_v I__1739 (
            .O(N__8460),
            .I(N__8445));
    Span4Mux_v I__1738 (
            .O(N__8455),
            .I(N__8445));
    Span4Mux_v I__1737 (
            .O(N__8450),
            .I(N__8442));
    Sp12to4 I__1736 (
            .O(N__8445),
            .I(N__8437));
    Sp12to4 I__1735 (
            .O(N__8442),
            .I(N__8437));
    Odrv12 I__1734 (
            .O(N__8437),
            .I(A_c_21));
    InMux I__1733 (
            .O(N__8434),
            .I(N__8430));
    InMux I__1732 (
            .O(N__8433),
            .I(N__8427));
    LocalMux I__1731 (
            .O(N__8430),
            .I(N__8424));
    LocalMux I__1730 (
            .O(N__8427),
            .I(N__8421));
    Span4Mux_v I__1729 (
            .O(N__8424),
            .I(N__8413));
    Span4Mux_v I__1728 (
            .O(N__8421),
            .I(N__8413));
    InMux I__1727 (
            .O(N__8420),
            .I(N__8410));
    InMux I__1726 (
            .O(N__8419),
            .I(N__8407));
    InMux I__1725 (
            .O(N__8418),
            .I(N__8404));
    Sp12to4 I__1724 (
            .O(N__8413),
            .I(N__8399));
    LocalMux I__1723 (
            .O(N__8410),
            .I(N__8399));
    LocalMux I__1722 (
            .O(N__8407),
            .I(N__8394));
    LocalMux I__1721 (
            .O(N__8404),
            .I(N__8394));
    Odrv12 I__1720 (
            .O(N__8399),
            .I(U409_ADDRESS_DECODE_ROMEN_1));
    Odrv4 I__1719 (
            .O(N__8394),
            .I(U409_ADDRESS_DECODE_ROMEN_1));
    InMux I__1718 (
            .O(N__8389),
            .I(N__8384));
    InMux I__1717 (
            .O(N__8388),
            .I(N__8381));
    CascadeMux I__1716 (
            .O(N__8387),
            .I(N__8378));
    LocalMux I__1715 (
            .O(N__8384),
            .I(N__8374));
    LocalMux I__1714 (
            .O(N__8381),
            .I(N__8371));
    InMux I__1713 (
            .O(N__8378),
            .I(N__8368));
    CascadeMux I__1712 (
            .O(N__8377),
            .I(N__8365));
    Span4Mux_v I__1711 (
            .O(N__8374),
            .I(N__8362));
    Span4Mux_h I__1710 (
            .O(N__8371),
            .I(N__8359));
    LocalMux I__1709 (
            .O(N__8368),
            .I(N__8356));
    InMux I__1708 (
            .O(N__8365),
            .I(N__8353));
    Span4Mux_h I__1707 (
            .O(N__8362),
            .I(N__8350));
    Span4Mux_h I__1706 (
            .O(N__8359),
            .I(N__8347));
    Span4Mux_h I__1705 (
            .O(N__8356),
            .I(N__8344));
    LocalMux I__1704 (
            .O(N__8353),
            .I(N__8341));
    Sp12to4 I__1703 (
            .O(N__8350),
            .I(N__8338));
    Sp12to4 I__1702 (
            .O(N__8347),
            .I(N__8333));
    Sp12to4 I__1701 (
            .O(N__8344),
            .I(N__8333));
    Span12Mux_h I__1700 (
            .O(N__8341),
            .I(N__8330));
    Span12Mux_h I__1699 (
            .O(N__8338),
            .I(N__8327));
    Span12Mux_v I__1698 (
            .O(N__8333),
            .I(N__8324));
    Span12Mux_v I__1697 (
            .O(N__8330),
            .I(N__8321));
    Span12Mux_v I__1696 (
            .O(N__8327),
            .I(N__8316));
    Span12Mux_h I__1695 (
            .O(N__8324),
            .I(N__8316));
    Odrv12 I__1694 (
            .O(N__8321),
            .I(OVL_c));
    Odrv12 I__1693 (
            .O(N__8316),
            .I(OVL_c));
    InMux I__1692 (
            .O(N__8311),
            .I(N__8308));
    LocalMux I__1691 (
            .O(N__8308),
            .I(N__8305));
    Span12Mux_v I__1690 (
            .O(N__8305),
            .I(N__8301));
    InMux I__1689 (
            .O(N__8304),
            .I(N__8298));
    Odrv12 I__1688 (
            .O(N__8301),
            .I(\U409_ADDRESS_DECODE.LOWROMZ0Z_3 ));
    LocalMux I__1687 (
            .O(N__8298),
            .I(\U409_ADDRESS_DECODE.LOWROMZ0Z_3 ));
    CascadeMux I__1686 (
            .O(N__8293),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn_cascade_));
    IoInMux I__1685 (
            .O(N__8290),
            .I(N__8287));
    LocalMux I__1684 (
            .O(N__8287),
            .I(N__8284));
    IoSpan4Mux I__1683 (
            .O(N__8284),
            .I(N__8281));
    IoSpan4Mux I__1682 (
            .O(N__8281),
            .I(N__8278));
    Span4Mux_s1_v I__1681 (
            .O(N__8278),
            .I(N__8275));
    Sp12to4 I__1680 (
            .O(N__8275),
            .I(N__8272));
    Odrv12 I__1679 (
            .O(N__8272),
            .I(PORTSIZE_0_i));
    CascadeMux I__1678 (
            .O(N__8269),
            .I(\U409_TRANSFER_ACK.G_14_0_o7_2_cascade_ ));
    InMux I__1677 (
            .O(N__8266),
            .I(N__8263));
    LocalMux I__1676 (
            .O(N__8263),
            .I(N__8260));
    Span4Mux_h I__1675 (
            .O(N__8260),
            .I(N__8257));
    Odrv4 I__1674 (
            .O(N__8257),
            .I(\U409_TRANSFER_ACK.G_14_0_o7_4 ));
    InMux I__1673 (
            .O(N__8254),
            .I(N__8248));
    CascadeMux I__1672 (
            .O(N__8253),
            .I(N__8245));
    CascadeMux I__1671 (
            .O(N__8252),
            .I(N__8242));
    InMux I__1670 (
            .O(N__8251),
            .I(N__8238));
    LocalMux I__1669 (
            .O(N__8248),
            .I(N__8233));
    InMux I__1668 (
            .O(N__8245),
            .I(N__8230));
    InMux I__1667 (
            .O(N__8242),
            .I(N__8227));
    CascadeMux I__1666 (
            .O(N__8241),
            .I(N__8224));
    LocalMux I__1665 (
            .O(N__8238),
            .I(N__8218));
    CascadeMux I__1664 (
            .O(N__8237),
            .I(N__8212));
    CascadeMux I__1663 (
            .O(N__8236),
            .I(N__8209));
    Span4Mux_h I__1662 (
            .O(N__8233),
            .I(N__8202));
    LocalMux I__1661 (
            .O(N__8230),
            .I(N__8202));
    LocalMux I__1660 (
            .O(N__8227),
            .I(N__8202));
    InMux I__1659 (
            .O(N__8224),
            .I(N__8199));
    InMux I__1658 (
            .O(N__8223),
            .I(N__8194));
    InMux I__1657 (
            .O(N__8222),
            .I(N__8194));
    InMux I__1656 (
            .O(N__8221),
            .I(N__8191));
    Span4Mux_v I__1655 (
            .O(N__8218),
            .I(N__8188));
    InMux I__1654 (
            .O(N__8217),
            .I(N__8183));
    InMux I__1653 (
            .O(N__8216),
            .I(N__8183));
    InMux I__1652 (
            .O(N__8215),
            .I(N__8180));
    InMux I__1651 (
            .O(N__8212),
            .I(N__8177));
    InMux I__1650 (
            .O(N__8209),
            .I(N__8174));
    Span4Mux_v I__1649 (
            .O(N__8202),
            .I(N__8167));
    LocalMux I__1648 (
            .O(N__8199),
            .I(N__8167));
    LocalMux I__1647 (
            .O(N__8194),
            .I(N__8167));
    LocalMux I__1646 (
            .O(N__8191),
            .I(N__8164));
    Span4Mux_v I__1645 (
            .O(N__8188),
            .I(N__8159));
    LocalMux I__1644 (
            .O(N__8183),
            .I(N__8159));
    LocalMux I__1643 (
            .O(N__8180),
            .I(N__8156));
    LocalMux I__1642 (
            .O(N__8177),
            .I(N__8153));
    LocalMux I__1641 (
            .O(N__8174),
            .I(N__8150));
    Span4Mux_v I__1640 (
            .O(N__8167),
            .I(N__8145));
    Span4Mux_v I__1639 (
            .O(N__8164),
            .I(N__8145));
    Span4Mux_h I__1638 (
            .O(N__8159),
            .I(N__8138));
    Span4Mux_v I__1637 (
            .O(N__8156),
            .I(N__8138));
    Span4Mux_v I__1636 (
            .O(N__8153),
            .I(N__8138));
    Span12Mux_v I__1635 (
            .O(N__8150),
            .I(N__8131));
    Sp12to4 I__1634 (
            .O(N__8145),
            .I(N__8131));
    Sp12to4 I__1633 (
            .O(N__8138),
            .I(N__8131));
    Odrv12 I__1632 (
            .O(N__8131),
            .I(A_c_20));
    CascadeMux I__1631 (
            .O(N__8128),
            .I(N__8123));
    CascadeMux I__1630 (
            .O(N__8127),
            .I(N__8120));
    InMux I__1629 (
            .O(N__8126),
            .I(N__8116));
    InMux I__1628 (
            .O(N__8123),
            .I(N__8113));
    InMux I__1627 (
            .O(N__8120),
            .I(N__8110));
    InMux I__1626 (
            .O(N__8119),
            .I(N__8107));
    LocalMux I__1625 (
            .O(N__8116),
            .I(ATA_BASE_7));
    LocalMux I__1624 (
            .O(N__8113),
            .I(ATA_BASE_7));
    LocalMux I__1623 (
            .O(N__8110),
            .I(ATA_BASE_7));
    LocalMux I__1622 (
            .O(N__8107),
            .I(ATA_BASE_7));
    InMux I__1621 (
            .O(N__8098),
            .I(N__8093));
    InMux I__1620 (
            .O(N__8097),
            .I(N__8089));
    InMux I__1619 (
            .O(N__8096),
            .I(N__8086));
    LocalMux I__1618 (
            .O(N__8093),
            .I(N__8083));
    InMux I__1617 (
            .O(N__8092),
            .I(N__8080));
    LocalMux I__1616 (
            .O(N__8089),
            .I(N__8077));
    LocalMux I__1615 (
            .O(N__8086),
            .I(ATA_BASE_4));
    Odrv4 I__1614 (
            .O(N__8083),
            .I(ATA_BASE_4));
    LocalMux I__1613 (
            .O(N__8080),
            .I(ATA_BASE_4));
    Odrv4 I__1612 (
            .O(N__8077),
            .I(ATA_BASE_4));
    InMux I__1611 (
            .O(N__8068),
            .I(N__8065));
    LocalMux I__1610 (
            .O(N__8065),
            .I(\U409_TRANSFER_ACK.G_14_0_o7_3 ));
    InMux I__1609 (
            .O(N__8062),
            .I(N__8059));
    LocalMux I__1608 (
            .O(N__8059),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_1_0 ));
    InMux I__1607 (
            .O(N__8056),
            .I(N__8052));
    InMux I__1606 (
            .O(N__8055),
            .I(N__8049));
    LocalMux I__1605 (
            .O(N__8052),
            .I(\U409_TRANSFER_ACK.N_13 ));
    LocalMux I__1604 (
            .O(N__8049),
            .I(\U409_TRANSFER_ACK.N_13 ));
    CascadeMux I__1603 (
            .O(N__8044),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20_cascade_ ));
    InMux I__1602 (
            .O(N__8041),
            .I(N__8037));
    CascadeMux I__1601 (
            .O(N__8040),
            .I(N__8034));
    LocalMux I__1600 (
            .O(N__8037),
            .I(N__8025));
    InMux I__1599 (
            .O(N__8034),
            .I(N__8022));
    InMux I__1598 (
            .O(N__8033),
            .I(N__8019));
    InMux I__1597 (
            .O(N__8032),
            .I(N__8014));
    InMux I__1596 (
            .O(N__8031),
            .I(N__8011));
    InMux I__1595 (
            .O(N__8030),
            .I(N__8005));
    InMux I__1594 (
            .O(N__8029),
            .I(N__8005));
    CascadeMux I__1593 (
            .O(N__8028),
            .I(N__8001));
    Span4Mux_h I__1592 (
            .O(N__8025),
            .I(N__7994));
    LocalMux I__1591 (
            .O(N__8022),
            .I(N__7994));
    LocalMux I__1590 (
            .O(N__8019),
            .I(N__7994));
    InMux I__1589 (
            .O(N__8018),
            .I(N__7991));
    InMux I__1588 (
            .O(N__8017),
            .I(N__7988));
    LocalMux I__1587 (
            .O(N__8014),
            .I(N__7983));
    LocalMux I__1586 (
            .O(N__8011),
            .I(N__7983));
    InMux I__1585 (
            .O(N__8010),
            .I(N__7980));
    LocalMux I__1584 (
            .O(N__8005),
            .I(N__7977));
    InMux I__1583 (
            .O(N__8004),
            .I(N__7974));
    InMux I__1582 (
            .O(N__8001),
            .I(N__7970));
    Span4Mux_v I__1581 (
            .O(N__7994),
            .I(N__7964));
    LocalMux I__1580 (
            .O(N__7991),
            .I(N__7964));
    LocalMux I__1579 (
            .O(N__7988),
            .I(N__7961));
    Span4Mux_v I__1578 (
            .O(N__7983),
            .I(N__7952));
    LocalMux I__1577 (
            .O(N__7980),
            .I(N__7952));
    Span4Mux_v I__1576 (
            .O(N__7977),
            .I(N__7952));
    LocalMux I__1575 (
            .O(N__7974),
            .I(N__7952));
    InMux I__1574 (
            .O(N__7973),
            .I(N__7949));
    LocalMux I__1573 (
            .O(N__7970),
            .I(N__7946));
    InMux I__1572 (
            .O(N__7969),
            .I(N__7943));
    Span4Mux_v I__1571 (
            .O(N__7964),
            .I(N__7940));
    Span4Mux_v I__1570 (
            .O(N__7961),
            .I(N__7933));
    Span4Mux_h I__1569 (
            .O(N__7952),
            .I(N__7933));
    LocalMux I__1568 (
            .O(N__7949),
            .I(N__7933));
    Sp12to4 I__1567 (
            .O(N__7946),
            .I(N__7928));
    LocalMux I__1566 (
            .O(N__7943),
            .I(N__7928));
    Span4Mux_h I__1565 (
            .O(N__7940),
            .I(N__7925));
    Span4Mux_v I__1564 (
            .O(N__7933),
            .I(N__7922));
    Span12Mux_v I__1563 (
            .O(N__7928),
            .I(N__7919));
    Sp12to4 I__1562 (
            .O(N__7925),
            .I(N__7914));
    Sp12to4 I__1561 (
            .O(N__7922),
            .I(N__7914));
    Odrv12 I__1560 (
            .O(N__7919),
            .I(A_c_23));
    Odrv12 I__1559 (
            .O(N__7914),
            .I(A_c_23));
    InMux I__1558 (
            .O(N__7909),
            .I(N__7906));
    LocalMux I__1557 (
            .O(N__7906),
            .I(N__7903));
    Odrv4 I__1556 (
            .O(N__7903),
            .I(\U409_TRANSFER_ACK.N_24 ));
    CascadeMux I__1555 (
            .O(N__7900),
            .I(N__7897));
    InMux I__1554 (
            .O(N__7897),
            .I(N__7894));
    LocalMux I__1553 (
            .O(N__7894),
            .I(N__7891));
    Span12Mux_h I__1552 (
            .O(N__7891),
            .I(N__7888));
    Odrv12 I__1551 (
            .O(N__7888),
            .I(\U409_TRANSFER_ACK.G_14_0_1_1 ));
    CascadeMux I__1550 (
            .O(N__7885),
            .I(\U409_TRANSFER_ACK.G_14_0_1_cascade_ ));
    CascadeMux I__1549 (
            .O(N__7882),
            .I(\U409_ADDRESS_DECODE.un2_REGSPACEn_0_0_cascade_ ));
    InMux I__1548 (
            .O(N__7879),
            .I(N__7871));
    InMux I__1547 (
            .O(N__7878),
            .I(N__7871));
    CascadeMux I__1546 (
            .O(N__7877),
            .I(N__7866));
    InMux I__1545 (
            .O(N__7876),
            .I(N__7863));
    LocalMux I__1544 (
            .O(N__7871),
            .I(N__7859));
    CascadeMux I__1543 (
            .O(N__7870),
            .I(N__7856));
    InMux I__1542 (
            .O(N__7869),
            .I(N__7851));
    InMux I__1541 (
            .O(N__7866),
            .I(N__7851));
    LocalMux I__1540 (
            .O(N__7863),
            .I(N__7848));
    InMux I__1539 (
            .O(N__7862),
            .I(N__7845));
    Span4Mux_v I__1538 (
            .O(N__7859),
            .I(N__7842));
    InMux I__1537 (
            .O(N__7856),
            .I(N__7839));
    LocalMux I__1536 (
            .O(N__7851),
            .I(N__7835));
    Span4Mux_v I__1535 (
            .O(N__7848),
            .I(N__7830));
    LocalMux I__1534 (
            .O(N__7845),
            .I(N__7830));
    Span4Mux_v I__1533 (
            .O(N__7842),
            .I(N__7825));
    LocalMux I__1532 (
            .O(N__7839),
            .I(N__7825));
    InMux I__1531 (
            .O(N__7838),
            .I(N__7819));
    Span4Mux_v I__1530 (
            .O(N__7835),
            .I(N__7816));
    Span4Mux_v I__1529 (
            .O(N__7830),
            .I(N__7813));
    Span4Mux_v I__1528 (
            .O(N__7825),
            .I(N__7810));
    InMux I__1527 (
            .O(N__7824),
            .I(N__7805));
    InMux I__1526 (
            .O(N__7823),
            .I(N__7805));
    InMux I__1525 (
            .O(N__7822),
            .I(N__7802));
    LocalMux I__1524 (
            .O(N__7819),
            .I(N__7789));
    Sp12to4 I__1523 (
            .O(N__7816),
            .I(N__7789));
    Sp12to4 I__1522 (
            .O(N__7813),
            .I(N__7789));
    Sp12to4 I__1521 (
            .O(N__7810),
            .I(N__7789));
    LocalMux I__1520 (
            .O(N__7805),
            .I(N__7789));
    LocalMux I__1519 (
            .O(N__7802),
            .I(N__7789));
    Span12Mux_h I__1518 (
            .O(N__7789),
            .I(N__7786));
    Span12Mux_v I__1517 (
            .O(N__7786),
            .I(N__7783));
    Odrv12 I__1516 (
            .O(N__7783),
            .I(A_c_19));
    CascadeMux I__1515 (
            .O(N__7780),
            .I(N__7774));
    CascadeMux I__1514 (
            .O(N__7779),
            .I(N__7771));
    CascadeMux I__1513 (
            .O(N__7778),
            .I(N__7767));
    CascadeMux I__1512 (
            .O(N__7777),
            .I(N__7764));
    InMux I__1511 (
            .O(N__7774),
            .I(N__7761));
    InMux I__1510 (
            .O(N__7771),
            .I(N__7758));
    InMux I__1509 (
            .O(N__7770),
            .I(N__7755));
    InMux I__1508 (
            .O(N__7767),
            .I(N__7750));
    InMux I__1507 (
            .O(N__7764),
            .I(N__7750));
    LocalMux I__1506 (
            .O(N__7761),
            .I(N__7747));
    LocalMux I__1505 (
            .O(N__7758),
            .I(N__7742));
    LocalMux I__1504 (
            .O(N__7755),
            .I(N__7742));
    LocalMux I__1503 (
            .O(N__7750),
            .I(N__7739));
    Span4Mux_v I__1502 (
            .O(N__7747),
            .I(N__7736));
    Span4Mux_v I__1501 (
            .O(N__7742),
            .I(N__7731));
    Span12Mux_v I__1500 (
            .O(N__7739),
            .I(N__7726));
    Sp12to4 I__1499 (
            .O(N__7736),
            .I(N__7726));
    InMux I__1498 (
            .O(N__7735),
            .I(N__7723));
    InMux I__1497 (
            .O(N__7734),
            .I(N__7720));
    Span4Mux_v I__1496 (
            .O(N__7731),
            .I(N__7717));
    Span12Mux_s11_h I__1495 (
            .O(N__7726),
            .I(N__7710));
    LocalMux I__1494 (
            .O(N__7723),
            .I(N__7710));
    LocalMux I__1493 (
            .O(N__7720),
            .I(N__7710));
    Span4Mux_v I__1492 (
            .O(N__7717),
            .I(N__7707));
    Span12Mux_v I__1491 (
            .O(N__7710),
            .I(N__7702));
    Sp12to4 I__1490 (
            .O(N__7707),
            .I(N__7702));
    Odrv12 I__1489 (
            .O(N__7702),
            .I(A_c_18));
    InMux I__1488 (
            .O(N__7699),
            .I(N__7696));
    LocalMux I__1487 (
            .O(N__7696),
            .I(\U409_ADDRESS_DECODE.REG_SPACEZ0Z_2 ));
    InMux I__1486 (
            .O(N__7693),
            .I(N__7690));
    LocalMux I__1485 (
            .O(N__7690),
            .I(\U409_ADDRESS_DECODE.REG_SPACE_3 ));
    InMux I__1484 (
            .O(N__7687),
            .I(N__7684));
    LocalMux I__1483 (
            .O(N__7684),
            .I(\U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0 ));
    IoInMux I__1482 (
            .O(N__7681),
            .I(N__7678));
    LocalMux I__1481 (
            .O(N__7678),
            .I(N__7675));
    Span12Mux_s0_v I__1480 (
            .O(N__7675),
            .I(N__7672));
    Span12Mux_v I__1479 (
            .O(N__7672),
            .I(N__7669));
    Odrv12 I__1478 (
            .O(N__7669),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn_i));
    InMux I__1477 (
            .O(N__7666),
            .I(N__7662));
    CascadeMux I__1476 (
            .O(N__7665),
            .I(N__7655));
    LocalMux I__1475 (
            .O(N__7662),
            .I(N__7651));
    InMux I__1474 (
            .O(N__7661),
            .I(N__7648));
    InMux I__1473 (
            .O(N__7660),
            .I(N__7645));
    InMux I__1472 (
            .O(N__7659),
            .I(N__7640));
    InMux I__1471 (
            .O(N__7658),
            .I(N__7640));
    InMux I__1470 (
            .O(N__7655),
            .I(N__7635));
    InMux I__1469 (
            .O(N__7654),
            .I(N__7635));
    Span4Mux_h I__1468 (
            .O(N__7651),
            .I(N__7630));
    LocalMux I__1467 (
            .O(N__7648),
            .I(N__7630));
    LocalMux I__1466 (
            .O(N__7645),
            .I(N__7625));
    LocalMux I__1465 (
            .O(N__7640),
            .I(N__7625));
    LocalMux I__1464 (
            .O(N__7635),
            .I(N__7622));
    Span4Mux_v I__1463 (
            .O(N__7630),
            .I(N__7616));
    Span4Mux_h I__1462 (
            .O(N__7625),
            .I(N__7616));
    Span4Mux_h I__1461 (
            .O(N__7622),
            .I(N__7613));
    InMux I__1460 (
            .O(N__7621),
            .I(N__7610));
    Sp12to4 I__1459 (
            .O(N__7616),
            .I(N__7603));
    Sp12to4 I__1458 (
            .O(N__7613),
            .I(N__7603));
    LocalMux I__1457 (
            .O(N__7610),
            .I(N__7603));
    Span12Mux_v I__1456 (
            .O(N__7603),
            .I(N__7600));
    Odrv12 I__1455 (
            .O(N__7600),
            .I(A_c_17));
    CascadeMux I__1454 (
            .O(N__7597),
            .I(N__7592));
    CascadeMux I__1453 (
            .O(N__7596),
            .I(N__7589));
    InMux I__1452 (
            .O(N__7595),
            .I(N__7585));
    InMux I__1451 (
            .O(N__7592),
            .I(N__7582));
    InMux I__1450 (
            .O(N__7589),
            .I(N__7577));
    InMux I__1449 (
            .O(N__7588),
            .I(N__7577));
    LocalMux I__1448 (
            .O(N__7585),
            .I(ATA_BASE_1));
    LocalMux I__1447 (
            .O(N__7582),
            .I(ATA_BASE_1));
    LocalMux I__1446 (
            .O(N__7577),
            .I(ATA_BASE_1));
    InMux I__1445 (
            .O(N__7570),
            .I(N__7566));
    InMux I__1444 (
            .O(N__7569),
            .I(N__7563));
    LocalMux I__1443 (
            .O(N__7566),
            .I(U409_ADDRESS_DECODE_un1_Z2_SPACE_7_2));
    LocalMux I__1442 (
            .O(N__7563),
            .I(U409_ADDRESS_DECODE_un1_Z2_SPACE_7_2));
    CascadeMux I__1441 (
            .O(N__7558),
            .I(N__7553));
    InMux I__1440 (
            .O(N__7557),
            .I(N__7549));
    InMux I__1439 (
            .O(N__7556),
            .I(N__7546));
    InMux I__1438 (
            .O(N__7553),
            .I(N__7541));
    InMux I__1437 (
            .O(N__7552),
            .I(N__7541));
    LocalMux I__1436 (
            .O(N__7549),
            .I(N__7537));
    LocalMux I__1435 (
            .O(N__7546),
            .I(N__7534));
    LocalMux I__1434 (
            .O(N__7541),
            .I(N__7531));
    InMux I__1433 (
            .O(N__7540),
            .I(N__7528));
    Span4Mux_v I__1432 (
            .O(N__7537),
            .I(N__7525));
    Span4Mux_v I__1431 (
            .O(N__7534),
            .I(N__7522));
    Span4Mux_v I__1430 (
            .O(N__7531),
            .I(N__7517));
    LocalMux I__1429 (
            .O(N__7528),
            .I(N__7517));
    Sp12to4 I__1428 (
            .O(N__7525),
            .I(N__7512));
    Sp12to4 I__1427 (
            .O(N__7522),
            .I(N__7512));
    Span4Mux_v I__1426 (
            .O(N__7517),
            .I(N__7509));
    Span12Mux_h I__1425 (
            .O(N__7512),
            .I(N__7506));
    Span4Mux_v I__1424 (
            .O(N__7509),
            .I(N__7503));
    Span12Mux_v I__1423 (
            .O(N__7506),
            .I(N__7500));
    Sp12to4 I__1422 (
            .O(N__7503),
            .I(N__7497));
    Odrv12 I__1421 (
            .O(N__7500),
            .I(A_c_16));
    Odrv12 I__1420 (
            .O(N__7497),
            .I(A_c_16));
    InMux I__1419 (
            .O(N__7492),
            .I(N__7483));
    InMux I__1418 (
            .O(N__7491),
            .I(N__7478));
    InMux I__1417 (
            .O(N__7490),
            .I(N__7475));
    InMux I__1416 (
            .O(N__7489),
            .I(N__7472));
    InMux I__1415 (
            .O(N__7488),
            .I(N__7469));
    InMux I__1414 (
            .O(N__7487),
            .I(N__7466));
    CascadeMux I__1413 (
            .O(N__7486),
            .I(N__7463));
    LocalMux I__1412 (
            .O(N__7483),
            .I(N__7458));
    InMux I__1411 (
            .O(N__7482),
            .I(N__7455));
    InMux I__1410 (
            .O(N__7481),
            .I(N__7452));
    LocalMux I__1409 (
            .O(N__7478),
            .I(N__7445));
    LocalMux I__1408 (
            .O(N__7475),
            .I(N__7445));
    LocalMux I__1407 (
            .O(N__7472),
            .I(N__7442));
    LocalMux I__1406 (
            .O(N__7469),
            .I(N__7439));
    LocalMux I__1405 (
            .O(N__7466),
            .I(N__7436));
    InMux I__1404 (
            .O(N__7463),
            .I(N__7433));
    InMux I__1403 (
            .O(N__7462),
            .I(N__7428));
    InMux I__1402 (
            .O(N__7461),
            .I(N__7428));
    Span4Mux_v I__1401 (
            .O(N__7458),
            .I(N__7421));
    LocalMux I__1400 (
            .O(N__7455),
            .I(N__7421));
    LocalMux I__1399 (
            .O(N__7452),
            .I(N__7421));
    InMux I__1398 (
            .O(N__7451),
            .I(N__7418));
    InMux I__1397 (
            .O(N__7450),
            .I(N__7415));
    Span4Mux_v I__1396 (
            .O(N__7445),
            .I(N__7411));
    Span4Mux_v I__1395 (
            .O(N__7442),
            .I(N__7406));
    Span4Mux_v I__1394 (
            .O(N__7439),
            .I(N__7406));
    Span4Mux_v I__1393 (
            .O(N__7436),
            .I(N__7403));
    LocalMux I__1392 (
            .O(N__7433),
            .I(N__7400));
    LocalMux I__1391 (
            .O(N__7428),
            .I(N__7397));
    Span4Mux_h I__1390 (
            .O(N__7421),
            .I(N__7390));
    LocalMux I__1389 (
            .O(N__7418),
            .I(N__7390));
    LocalMux I__1388 (
            .O(N__7415),
            .I(N__7390));
    InMux I__1387 (
            .O(N__7414),
            .I(N__7387));
    Sp12to4 I__1386 (
            .O(N__7411),
            .I(N__7382));
    Sp12to4 I__1385 (
            .O(N__7406),
            .I(N__7382));
    Span4Mux_v I__1384 (
            .O(N__7403),
            .I(N__7379));
    Span4Mux_v I__1383 (
            .O(N__7400),
            .I(N__7370));
    Span4Mux_h I__1382 (
            .O(N__7397),
            .I(N__7370));
    Span4Mux_v I__1381 (
            .O(N__7390),
            .I(N__7370));
    LocalMux I__1380 (
            .O(N__7387),
            .I(N__7370));
    Span12Mux_h I__1379 (
            .O(N__7382),
            .I(N__7367));
    Span4Mux_v I__1378 (
            .O(N__7379),
            .I(N__7364));
    Sp12to4 I__1377 (
            .O(N__7370),
            .I(N__7361));
    Span12Mux_v I__1376 (
            .O(N__7367),
            .I(N__7358));
    Sp12to4 I__1375 (
            .O(N__7364),
            .I(N__7353));
    Span12Mux_v I__1374 (
            .O(N__7361),
            .I(N__7353));
    Odrv12 I__1373 (
            .O(N__7358),
            .I(A_c_22));
    Odrv12 I__1372 (
            .O(N__7353),
            .I(A_c_22));
    CascadeMux I__1371 (
            .O(N__7348),
            .I(N__7345));
    InMux I__1370 (
            .O(N__7345),
            .I(N__7339));
    InMux I__1369 (
            .O(N__7344),
            .I(N__7336));
    InMux I__1368 (
            .O(N__7343),
            .I(N__7331));
    InMux I__1367 (
            .O(N__7342),
            .I(N__7331));
    LocalMux I__1366 (
            .O(N__7339),
            .I(ATA_BASE_0));
    LocalMux I__1365 (
            .O(N__7336),
            .I(ATA_BASE_0));
    LocalMux I__1364 (
            .O(N__7331),
            .I(ATA_BASE_0));
    CascadeMux I__1363 (
            .O(N__7324),
            .I(N__7319));
    InMux I__1362 (
            .O(N__7323),
            .I(N__7315));
    InMux I__1361 (
            .O(N__7322),
            .I(N__7312));
    InMux I__1360 (
            .O(N__7319),
            .I(N__7309));
    InMux I__1359 (
            .O(N__7318),
            .I(N__7306));
    LocalMux I__1358 (
            .O(N__7315),
            .I(ATA_BASE_6));
    LocalMux I__1357 (
            .O(N__7312),
            .I(ATA_BASE_6));
    LocalMux I__1356 (
            .O(N__7309),
            .I(ATA_BASE_6));
    LocalMux I__1355 (
            .O(N__7306),
            .I(ATA_BASE_6));
    InMux I__1354 (
            .O(N__7297),
            .I(N__7279));
    InMux I__1353 (
            .O(N__7296),
            .I(N__7279));
    InMux I__1352 (
            .O(N__7295),
            .I(N__7279));
    InMux I__1351 (
            .O(N__7294),
            .I(N__7279));
    InMux I__1350 (
            .O(N__7293),
            .I(N__7279));
    InMux I__1349 (
            .O(N__7292),
            .I(N__7279));
    LocalMux I__1348 (
            .O(N__7279),
            .I(N__7274));
    InMux I__1347 (
            .O(N__7278),
            .I(N__7271));
    CascadeMux I__1346 (
            .O(N__7277),
            .I(N__7268));
    Span4Mux_v I__1345 (
            .O(N__7274),
            .I(N__7261));
    LocalMux I__1344 (
            .O(N__7271),
            .I(N__7258));
    InMux I__1343 (
            .O(N__7268),
            .I(N__7247));
    InMux I__1342 (
            .O(N__7267),
            .I(N__7247));
    InMux I__1341 (
            .O(N__7266),
            .I(N__7247));
    InMux I__1340 (
            .O(N__7265),
            .I(N__7247));
    InMux I__1339 (
            .O(N__7264),
            .I(N__7247));
    Odrv4 I__1338 (
            .O(N__7261),
            .I(un1_AUTOCONFIG_SPACE));
    Odrv4 I__1337 (
            .O(N__7258),
            .I(un1_AUTOCONFIG_SPACE));
    LocalMux I__1336 (
            .O(N__7247),
            .I(un1_AUTOCONFIG_SPACE));
    InMux I__1335 (
            .O(N__7240),
            .I(N__7237));
    LocalMux I__1334 (
            .O(N__7237),
            .I(N__7231));
    InMux I__1333 (
            .O(N__7236),
            .I(N__7224));
    InMux I__1332 (
            .O(N__7235),
            .I(N__7224));
    InMux I__1331 (
            .O(N__7234),
            .I(N__7224));
    Odrv4 I__1330 (
            .O(N__7231),
            .I(\U409_AUTOCONFIG.STATE_RNI0FVT2Z0Z_0 ));
    LocalMux I__1329 (
            .O(N__7224),
            .I(\U409_AUTOCONFIG.STATE_RNI0FVT2Z0Z_0 ));
    CascadeMux I__1328 (
            .O(N__7219),
            .I(N__7214));
    InMux I__1327 (
            .O(N__7218),
            .I(N__7209));
    InMux I__1326 (
            .O(N__7217),
            .I(N__7209));
    InMux I__1325 (
            .O(N__7214),
            .I(N__7206));
    LocalMux I__1324 (
            .O(N__7209),
            .I(N__7203));
    LocalMux I__1323 (
            .O(N__7206),
            .I(N__7200));
    Span4Mux_v I__1322 (
            .O(N__7203),
            .I(N__7195));
    Span4Mux_v I__1321 (
            .O(N__7200),
            .I(N__7195));
    Sp12to4 I__1320 (
            .O(N__7195),
            .I(N__7192));
    Span12Mux_h I__1319 (
            .O(N__7192),
            .I(N__7189));
    Odrv12 I__1318 (
            .O(N__7189),
            .I(D_in_7));
    CascadeMux I__1317 (
            .O(N__7186),
            .I(N__7181));
    InMux I__1316 (
            .O(N__7185),
            .I(N__7178));
    InMux I__1315 (
            .O(N__7184),
            .I(N__7175));
    InMux I__1314 (
            .O(N__7181),
            .I(N__7172));
    LocalMux I__1313 (
            .O(N__7178),
            .I(ATA_BASE_3));
    LocalMux I__1312 (
            .O(N__7175),
            .I(ATA_BASE_3));
    LocalMux I__1311 (
            .O(N__7172),
            .I(ATA_BASE_3));
    CascadeMux I__1310 (
            .O(N__7165),
            .I(N__7162));
    InMux I__1309 (
            .O(N__7162),
            .I(N__7159));
    LocalMux I__1308 (
            .O(N__7159),
            .I(U409_ADDRESS_DECODE_ATA_ROM_d));
    InMux I__1307 (
            .O(N__7156),
            .I(N__7153));
    LocalMux I__1306 (
            .O(N__7153),
            .I(N__7150));
    Odrv4 I__1305 (
            .O(N__7150),
            .I(\U409_ADDRESS_DECODE.g0_i_0Z0Z_0 ));
    InMux I__1304 (
            .O(N__7147),
            .I(N__7144));
    LocalMux I__1303 (
            .O(N__7144),
            .I(N__7141));
    Odrv4 I__1302 (
            .O(N__7141),
            .I(\U409_ADDRESS_DECODE.g0_i_o4Z0Z_1 ));
    InMux I__1301 (
            .O(N__7138),
            .I(N__7135));
    LocalMux I__1300 (
            .O(N__7135),
            .I(\U409_ADDRESS_DECODE.g0_i_o4Z0Z_0 ));
    InMux I__1299 (
            .O(N__7132),
            .I(N__7129));
    LocalMux I__1298 (
            .O(N__7129),
            .I(U409_ADDRESS_DECODE_ATA_ROM_0_1));
    CascadeMux I__1297 (
            .O(N__7126),
            .I(N__7122));
    InMux I__1296 (
            .O(N__7125),
            .I(N__7117));
    InMux I__1295 (
            .O(N__7122),
            .I(N__7117));
    LocalMux I__1294 (
            .O(N__7117),
            .I(N__7114));
    Odrv4 I__1293 (
            .O(N__7114),
            .I(\U409_TRANSFER_ACK.CO1 ));
    InMux I__1292 (
            .O(N__7111),
            .I(N__7106));
    InMux I__1291 (
            .O(N__7110),
            .I(N__7103));
    InMux I__1290 (
            .O(N__7109),
            .I(N__7100));
    LocalMux I__1289 (
            .O(N__7106),
            .I(N__7096));
    LocalMux I__1288 (
            .O(N__7103),
            .I(N__7093));
    LocalMux I__1287 (
            .O(N__7100),
            .I(N__7090));
    InMux I__1286 (
            .O(N__7099),
            .I(N__7087));
    Span4Mux_h I__1285 (
            .O(N__7096),
            .I(N__7076));
    Span4Mux_v I__1284 (
            .O(N__7093),
            .I(N__7076));
    Span4Mux_v I__1283 (
            .O(N__7090),
            .I(N__7076));
    LocalMux I__1282 (
            .O(N__7087),
            .I(N__7076));
    InMux I__1281 (
            .O(N__7086),
            .I(N__7073));
    CascadeMux I__1280 (
            .O(N__7085),
            .I(N__7070));
    Span4Mux_v I__1279 (
            .O(N__7076),
            .I(N__7065));
    LocalMux I__1278 (
            .O(N__7073),
            .I(N__7065));
    InMux I__1277 (
            .O(N__7070),
            .I(N__7062));
    Span4Mux_v I__1276 (
            .O(N__7065),
            .I(N__7059));
    LocalMux I__1275 (
            .O(N__7062),
            .I(N__7056));
    Span4Mux_v I__1274 (
            .O(N__7059),
            .I(N__7053));
    Span12Mux_h I__1273 (
            .O(N__7056),
            .I(N__7050));
    IoSpan4Mux I__1272 (
            .O(N__7053),
            .I(N__7047));
    Odrv12 I__1271 (
            .O(N__7050),
            .I(TM_c_1));
    Odrv4 I__1270 (
            .O(N__7047),
            .I(TM_c_1));
    CascadeMux I__1269 (
            .O(N__7042),
            .I(N__7037));
    InMux I__1268 (
            .O(N__7041),
            .I(N__7034));
    InMux I__1267 (
            .O(N__7040),
            .I(N__7031));
    InMux I__1266 (
            .O(N__7037),
            .I(N__7026));
    LocalMux I__1265 (
            .O(N__7034),
            .I(N__7023));
    LocalMux I__1264 (
            .O(N__7031),
            .I(N__7020));
    InMux I__1263 (
            .O(N__7030),
            .I(N__7017));
    InMux I__1262 (
            .O(N__7029),
            .I(N__7014));
    LocalMux I__1261 (
            .O(N__7026),
            .I(N__7010));
    Span4Mux_v I__1260 (
            .O(N__7023),
            .I(N__7001));
    Span4Mux_v I__1259 (
            .O(N__7020),
            .I(N__7001));
    LocalMux I__1258 (
            .O(N__7017),
            .I(N__7001));
    LocalMux I__1257 (
            .O(N__7014),
            .I(N__7001));
    InMux I__1256 (
            .O(N__7013),
            .I(N__6998));
    Span4Mux_v I__1255 (
            .O(N__7010),
            .I(N__6995));
    Span4Mux_v I__1254 (
            .O(N__7001),
            .I(N__6990));
    LocalMux I__1253 (
            .O(N__6998),
            .I(N__6990));
    Sp12to4 I__1252 (
            .O(N__6995),
            .I(N__6987));
    Span4Mux_h I__1251 (
            .O(N__6990),
            .I(N__6984));
    Span12Mux_h I__1250 (
            .O(N__6987),
            .I(N__6981));
    Span4Mux_v I__1249 (
            .O(N__6984),
            .I(N__6978));
    Span12Mux_v I__1248 (
            .O(N__6981),
            .I(N__6975));
    Span4Mux_v I__1247 (
            .O(N__6978),
            .I(N__6972));
    Odrv12 I__1246 (
            .O(N__6975),
            .I(TM_c_0));
    Odrv4 I__1245 (
            .O(N__6972),
            .I(TM_c_0));
    InMux I__1244 (
            .O(N__6967),
            .I(N__6961));
    InMux I__1243 (
            .O(N__6966),
            .I(N__6961));
    LocalMux I__1242 (
            .O(N__6961),
            .I(N__6958));
    Odrv12 I__1241 (
            .O(N__6958),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2 ));
    InMux I__1240 (
            .O(N__6955),
            .I(N__6952));
    LocalMux I__1239 (
            .O(N__6952),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3 ));
    CascadeMux I__1238 (
            .O(N__6949),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3_cascade_ ));
    InMux I__1237 (
            .O(N__6946),
            .I(N__6941));
    InMux I__1236 (
            .O(N__6945),
            .I(N__6936));
    InMux I__1235 (
            .O(N__6944),
            .I(N__6936));
    LocalMux I__1234 (
            .O(N__6941),
            .I(ATA_BASE_2));
    LocalMux I__1233 (
            .O(N__6936),
            .I(ATA_BASE_2));
    CascadeMux I__1232 (
            .O(N__6931),
            .I(N__6927));
    CascadeMux I__1231 (
            .O(N__6930),
            .I(N__6923));
    InMux I__1230 (
            .O(N__6927),
            .I(N__6920));
    InMux I__1229 (
            .O(N__6926),
            .I(N__6915));
    InMux I__1228 (
            .O(N__6923),
            .I(N__6915));
    LocalMux I__1227 (
            .O(N__6920),
            .I(N__6912));
    LocalMux I__1226 (
            .O(N__6915),
            .I(N__6909));
    Span4Mux_v I__1225 (
            .O(N__6912),
            .I(N__6906));
    Span4Mux_v I__1224 (
            .O(N__6909),
            .I(N__6903));
    Sp12to4 I__1223 (
            .O(N__6906),
            .I(N__6900));
    Sp12to4 I__1222 (
            .O(N__6903),
            .I(N__6895));
    Span12Mux_h I__1221 (
            .O(N__6900),
            .I(N__6895));
    Odrv12 I__1220 (
            .O(N__6895),
            .I(D_in_4));
    CascadeMux I__1219 (
            .O(N__6892),
            .I(N__6888));
    CascadeMux I__1218 (
            .O(N__6891),
            .I(N__6885));
    InMux I__1217 (
            .O(N__6888),
            .I(N__6880));
    InMux I__1216 (
            .O(N__6885),
            .I(N__6880));
    LocalMux I__1215 (
            .O(N__6880),
            .I(N__6877));
    Span4Mux_h I__1214 (
            .O(N__6877),
            .I(N__6874));
    Span4Mux_v I__1213 (
            .O(N__6874),
            .I(N__6870));
    InMux I__1212 (
            .O(N__6873),
            .I(N__6867));
    Span4Mux_v I__1211 (
            .O(N__6870),
            .I(N__6864));
    LocalMux I__1210 (
            .O(N__6867),
            .I(N__6861));
    Span4Mux_v I__1209 (
            .O(N__6864),
            .I(N__6858));
    Span12Mux_v I__1208 (
            .O(N__6861),
            .I(N__6855));
    Odrv4 I__1207 (
            .O(N__6858),
            .I(D_in_5));
    Odrv12 I__1206 (
            .O(N__6855),
            .I(D_in_5));
    InMux I__1205 (
            .O(N__6850),
            .I(N__6847));
    LocalMux I__1204 (
            .O(N__6847),
            .I(N__6843));
    CascadeMux I__1203 (
            .O(N__6846),
            .I(N__6840));
    Span4Mux_v I__1202 (
            .O(N__6843),
            .I(N__6837));
    InMux I__1201 (
            .O(N__6840),
            .I(N__6833));
    Span4Mux_v I__1200 (
            .O(N__6837),
            .I(N__6830));
    InMux I__1199 (
            .O(N__6836),
            .I(N__6827));
    LocalMux I__1198 (
            .O(N__6833),
            .I(N__6824));
    Sp12to4 I__1197 (
            .O(N__6830),
            .I(N__6821));
    LocalMux I__1196 (
            .O(N__6827),
            .I(N__6818));
    Span4Mux_v I__1195 (
            .O(N__6824),
            .I(N__6815));
    Span12Mux_h I__1194 (
            .O(N__6821),
            .I(N__6808));
    Span12Mux_v I__1193 (
            .O(N__6818),
            .I(N__6808));
    Sp12to4 I__1192 (
            .O(N__6815),
            .I(N__6808));
    Odrv12 I__1191 (
            .O(N__6808),
            .I(D_in_6));
    InMux I__1190 (
            .O(N__6805),
            .I(N__6797));
    InMux I__1189 (
            .O(N__6804),
            .I(N__6797));
    InMux I__1188 (
            .O(N__6803),
            .I(N__6792));
    InMux I__1187 (
            .O(N__6802),
            .I(N__6792));
    LocalMux I__1186 (
            .O(N__6797),
            .I(\U409_AUTOCONFIG.LIDE_CONF_RNIHQ9AZ0Z3 ));
    LocalMux I__1185 (
            .O(N__6792),
            .I(\U409_AUTOCONFIG.LIDE_CONF_RNIHQ9AZ0Z3 ));
    InMux I__1184 (
            .O(N__6787),
            .I(N__6783));
    CascadeMux I__1183 (
            .O(N__6786),
            .I(N__6779));
    LocalMux I__1182 (
            .O(N__6783),
            .I(N__6773));
    InMux I__1181 (
            .O(N__6782),
            .I(N__6770));
    InMux I__1180 (
            .O(N__6779),
            .I(N__6765));
    InMux I__1179 (
            .O(N__6778),
            .I(N__6765));
    InMux I__1178 (
            .O(N__6777),
            .I(N__6760));
    InMux I__1177 (
            .O(N__6776),
            .I(N__6760));
    Span4Mux_h I__1176 (
            .O(N__6773),
            .I(N__6757));
    LocalMux I__1175 (
            .O(N__6770),
            .I(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ));
    LocalMux I__1174 (
            .O(N__6765),
            .I(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ));
    LocalMux I__1173 (
            .O(N__6760),
            .I(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ));
    Odrv4 I__1172 (
            .O(N__6757),
            .I(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ));
    InMux I__1171 (
            .O(N__6748),
            .I(N__6744));
    CascadeMux I__1170 (
            .O(N__6747),
            .I(N__6741));
    LocalMux I__1169 (
            .O(N__6744),
            .I(N__6738));
    InMux I__1168 (
            .O(N__6741),
            .I(N__6735));
    Odrv4 I__1167 (
            .O(N__6738),
            .I(BRIDGE_BASE_3));
    LocalMux I__1166 (
            .O(N__6735),
            .I(BRIDGE_BASE_3));
    IoInMux I__1165 (
            .O(N__6730),
            .I(N__6727));
    LocalMux I__1164 (
            .O(N__6727),
            .I(N__6724));
    Span4Mux_s1_v I__1163 (
            .O(N__6724),
            .I(N__6721));
    Sp12to4 I__1162 (
            .O(N__6721),
            .I(N__6718));
    Span12Mux_h I__1161 (
            .O(N__6718),
            .I(N__6711));
    InMux I__1160 (
            .O(N__6717),
            .I(N__6707));
    InMux I__1159 (
            .O(N__6716),
            .I(N__6704));
    InMux I__1158 (
            .O(N__6715),
            .I(N__6699));
    InMux I__1157 (
            .O(N__6714),
            .I(N__6699));
    Span12Mux_v I__1156 (
            .O(N__6711),
            .I(N__6695));
    InMux I__1155 (
            .O(N__6710),
            .I(N__6692));
    LocalMux I__1154 (
            .O(N__6707),
            .I(N__6687));
    LocalMux I__1153 (
            .O(N__6704),
            .I(N__6687));
    LocalMux I__1152 (
            .O(N__6699),
            .I(N__6684));
    InMux I__1151 (
            .O(N__6698),
            .I(N__6681));
    Odrv12 I__1150 (
            .O(N__6695),
            .I(CONFIGENn_c));
    LocalMux I__1149 (
            .O(N__6692),
            .I(CONFIGENn_c));
    Odrv12 I__1148 (
            .O(N__6687),
            .I(CONFIGENn_c));
    Odrv4 I__1147 (
            .O(N__6684),
            .I(CONFIGENn_c));
    LocalMux I__1146 (
            .O(N__6681),
            .I(CONFIGENn_c));
    CascadeMux I__1145 (
            .O(N__6670),
            .I(N__6666));
    InMux I__1144 (
            .O(N__6669),
            .I(N__6663));
    InMux I__1143 (
            .O(N__6666),
            .I(N__6660));
    LocalMux I__1142 (
            .O(N__6663),
            .I(N__6653));
    LocalMux I__1141 (
            .O(N__6660),
            .I(N__6653));
    InMux I__1140 (
            .O(N__6659),
            .I(N__6650));
    InMux I__1139 (
            .O(N__6658),
            .I(N__6647));
    Odrv4 I__1138 (
            .O(N__6653),
            .I(ATA_BASE_5));
    LocalMux I__1137 (
            .O(N__6650),
            .I(ATA_BASE_5));
    LocalMux I__1136 (
            .O(N__6647),
            .I(ATA_BASE_5));
    InMux I__1135 (
            .O(N__6640),
            .I(N__6637));
    LocalMux I__1134 (
            .O(N__6637),
            .I(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_0 ));
    CascadeMux I__1133 (
            .O(N__6634),
            .I(N__6631));
    InMux I__1132 (
            .O(N__6631),
            .I(N__6628));
    LocalMux I__1131 (
            .O(N__6628),
            .I(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_4 ));
    InMux I__1130 (
            .O(N__6625),
            .I(N__6622));
    LocalMux I__1129 (
            .O(N__6622),
            .I(N__6616));
    InMux I__1128 (
            .O(N__6621),
            .I(N__6611));
    InMux I__1127 (
            .O(N__6620),
            .I(N__6611));
    InMux I__1126 (
            .O(N__6619),
            .I(N__6608));
    Span4Mux_h I__1125 (
            .O(N__6616),
            .I(N__6604));
    LocalMux I__1124 (
            .O(N__6611),
            .I(N__6599));
    LocalMux I__1123 (
            .O(N__6608),
            .I(N__6599));
    InMux I__1122 (
            .O(N__6607),
            .I(N__6596));
    Span4Mux_v I__1121 (
            .O(N__6604),
            .I(N__6589));
    Span4Mux_h I__1120 (
            .O(N__6599),
            .I(N__6589));
    LocalMux I__1119 (
            .O(N__6596),
            .I(N__6589));
    Span4Mux_h I__1118 (
            .O(N__6589),
            .I(N__6586));
    Span4Mux_v I__1117 (
            .O(N__6586),
            .I(N__6583));
    Odrv4 I__1116 (
            .O(N__6583),
            .I(A_c_31));
    IoInMux I__1115 (
            .O(N__6580),
            .I(N__6577));
    LocalMux I__1114 (
            .O(N__6577),
            .I(N__6574));
    Span12Mux_s9_h I__1113 (
            .O(N__6574),
            .I(N__6571));
    Span12Mux_h I__1112 (
            .O(N__6571),
            .I(N__6568));
    Odrv12 I__1111 (
            .O(N__6568),
            .I(U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i));
    InMux I__1110 (
            .O(N__6565),
            .I(N__6561));
    InMux I__1109 (
            .O(N__6564),
            .I(N__6558));
    LocalMux I__1108 (
            .O(N__6561),
            .I(N__6555));
    LocalMux I__1107 (
            .O(N__6558),
            .I(N__6552));
    Span4Mux_v I__1106 (
            .O(N__6555),
            .I(N__6549));
    Odrv12 I__1105 (
            .O(N__6552),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6 ));
    Odrv4 I__1104 (
            .O(N__6549),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6 ));
    CascadeMux I__1103 (
            .O(N__6544),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0_cascade_ ));
    InMux I__1102 (
            .O(N__6541),
            .I(N__6538));
    LocalMux I__1101 (
            .O(N__6538),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ));
    InMux I__1100 (
            .O(N__6535),
            .I(N__6532));
    LocalMux I__1099 (
            .O(N__6532),
            .I(\U409_ADDRESS_DECODE.g2Z0Z_5 ));
    InMux I__1098 (
            .O(N__6529),
            .I(N__6524));
    InMux I__1097 (
            .O(N__6528),
            .I(N__6521));
    InMux I__1096 (
            .O(N__6527),
            .I(N__6518));
    LocalMux I__1095 (
            .O(N__6524),
            .I(N__6514));
    LocalMux I__1094 (
            .O(N__6521),
            .I(N__6511));
    LocalMux I__1093 (
            .O(N__6518),
            .I(N__6508));
    InMux I__1092 (
            .O(N__6517),
            .I(N__6504));
    Span4Mux_h I__1091 (
            .O(N__6514),
            .I(N__6499));
    Span4Mux_v I__1090 (
            .O(N__6511),
            .I(N__6499));
    Span4Mux_h I__1089 (
            .O(N__6508),
            .I(N__6496));
    InMux I__1088 (
            .O(N__6507),
            .I(N__6493));
    LocalMux I__1087 (
            .O(N__6504),
            .I(N__6490));
    Span4Mux_v I__1086 (
            .O(N__6499),
            .I(N__6487));
    Span4Mux_v I__1085 (
            .O(N__6496),
            .I(N__6482));
    LocalMux I__1084 (
            .O(N__6493),
            .I(N__6482));
    Sp12to4 I__1083 (
            .O(N__6490),
            .I(N__6479));
    Span4Mux_v I__1082 (
            .O(N__6487),
            .I(N__6476));
    Sp12to4 I__1081 (
            .O(N__6482),
            .I(N__6473));
    Span12Mux_v I__1080 (
            .O(N__6479),
            .I(N__6470));
    Sp12to4 I__1079 (
            .O(N__6476),
            .I(N__6465));
    Span12Mux_v I__1078 (
            .O(N__6473),
            .I(N__6465));
    Odrv12 I__1077 (
            .O(N__6470),
            .I(A_c_28));
    Odrv12 I__1076 (
            .O(N__6465),
            .I(A_c_28));
    InMux I__1075 (
            .O(N__6460),
            .I(N__6457));
    LocalMux I__1074 (
            .O(N__6457),
            .I(U409_ADDRESS_DECODE_g2_6));
    CascadeMux I__1073 (
            .O(N__6454),
            .I(U409_ADDRESS_DECODE_g2_7_cascade_));
    InMux I__1072 (
            .O(N__6451),
            .I(N__6448));
    LocalMux I__1071 (
            .O(N__6448),
            .I(N__6445));
    Odrv12 I__1070 (
            .O(N__6445),
            .I(\U409_TRANSFER_ACK.G_14_0_o7_0 ));
    IoInMux I__1069 (
            .O(N__6442),
            .I(N__6439));
    LocalMux I__1068 (
            .O(N__6439),
            .I(N__6436));
    Span4Mux_s0_h I__1067 (
            .O(N__6436),
            .I(N__6433));
    Sp12to4 I__1066 (
            .O(N__6433),
            .I(N__6430));
    Span12Mux_s11_v I__1065 (
            .O(N__6430),
            .I(N__6427));
    Span12Mux_h I__1064 (
            .O(N__6427),
            .I(N__6424));
    Odrv12 I__1063 (
            .O(N__6424),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn_i));
    InMux I__1062 (
            .O(N__6421),
            .I(N__6418));
    LocalMux I__1061 (
            .O(N__6418),
            .I(\U409_ADDRESS_DECODE.un1_Z2_SPACE_6Z0Z_1 ));
    InMux I__1060 (
            .O(N__6415),
            .I(N__6412));
    LocalMux I__1059 (
            .O(N__6412),
            .I(\U409_ADDRESS_DECODE.un1_Z2_SPACE_6Z0Z_0 ));
    CascadeMux I__1058 (
            .O(N__6409),
            .I(\U409_ADDRESS_DECODE.un1_Z2_SPACE_7Z0Z_3_cascade_ ));
    CascadeMux I__1057 (
            .O(N__6406),
            .I(N__6403));
    InMux I__1056 (
            .O(N__6403),
            .I(N__6397));
    InMux I__1055 (
            .O(N__6402),
            .I(N__6391));
    InMux I__1054 (
            .O(N__6401),
            .I(N__6391));
    InMux I__1053 (
            .O(N__6400),
            .I(N__6388));
    LocalMux I__1052 (
            .O(N__6397),
            .I(N__6384));
    InMux I__1051 (
            .O(N__6396),
            .I(N__6381));
    LocalMux I__1050 (
            .O(N__6391),
            .I(N__6376));
    LocalMux I__1049 (
            .O(N__6388),
            .I(N__6376));
    CascadeMux I__1048 (
            .O(N__6387),
            .I(N__6373));
    Span4Mux_v I__1047 (
            .O(N__6384),
            .I(N__6367));
    LocalMux I__1046 (
            .O(N__6381),
            .I(N__6367));
    Span4Mux_v I__1045 (
            .O(N__6376),
            .I(N__6364));
    InMux I__1044 (
            .O(N__6373),
            .I(N__6361));
    InMux I__1043 (
            .O(N__6372),
            .I(N__6358));
    Span4Mux_v I__1042 (
            .O(N__6367),
            .I(N__6355));
    Sp12to4 I__1041 (
            .O(N__6364),
            .I(N__6348));
    LocalMux I__1040 (
            .O(N__6361),
            .I(N__6348));
    LocalMux I__1039 (
            .O(N__6358),
            .I(N__6348));
    Sp12to4 I__1038 (
            .O(N__6355),
            .I(N__6345));
    Span12Mux_h I__1037 (
            .O(N__6348),
            .I(N__6342));
    Span12Mux_h I__1036 (
            .O(N__6345),
            .I(N__6339));
    Span12Mux_v I__1035 (
            .O(N__6342),
            .I(N__6336));
    Span12Mux_v I__1034 (
            .O(N__6339),
            .I(N__6333));
    Odrv12 I__1033 (
            .O(N__6336),
            .I(RnW_c));
    Odrv12 I__1032 (
            .O(N__6333),
            .I(RnW_c));
    CascadeMux I__1031 (
            .O(N__6328),
            .I(\U409_ADDRESS_DECODE.un1_Z2_SPACEZ0_cascade_ ));
    InMux I__1030 (
            .O(N__6325),
            .I(N__6322));
    LocalMux I__1029 (
            .O(N__6322),
            .I(N__6319));
    Odrv4 I__1028 (
            .O(N__6319),
            .I(\U409_ADDRESS_DECODE.g2Z0Z_10 ));
    CascadeMux I__1027 (
            .O(N__6316),
            .I(\U409_ADDRESS_DECODE.g2Z0Z_11_cascade_ ));
    InMux I__1026 (
            .O(N__6313),
            .I(N__6310));
    LocalMux I__1025 (
            .O(N__6310),
            .I(N__6307));
    Span4Mux_v I__1024 (
            .O(N__6307),
            .I(N__6304));
    Odrv4 I__1023 (
            .O(N__6304),
            .I(\U409_ADDRESS_DECODE.g2Z0Z_9 ));
    InMux I__1022 (
            .O(N__6301),
            .I(N__6289));
    InMux I__1021 (
            .O(N__6300),
            .I(N__6289));
    CascadeMux I__1020 (
            .O(N__6299),
            .I(N__6285));
    CascadeMux I__1019 (
            .O(N__6298),
            .I(N__6282));
    CascadeMux I__1018 (
            .O(N__6297),
            .I(N__6279));
    CascadeMux I__1017 (
            .O(N__6296),
            .I(N__6276));
    InMux I__1016 (
            .O(N__6295),
            .I(N__6271));
    InMux I__1015 (
            .O(N__6294),
            .I(N__6271));
    LocalMux I__1014 (
            .O(N__6289),
            .I(N__6267));
    InMux I__1013 (
            .O(N__6288),
            .I(N__6262));
    InMux I__1012 (
            .O(N__6285),
            .I(N__6262));
    InMux I__1011 (
            .O(N__6282),
            .I(N__6257));
    InMux I__1010 (
            .O(N__6279),
            .I(N__6257));
    InMux I__1009 (
            .O(N__6276),
            .I(N__6254));
    LocalMux I__1008 (
            .O(N__6271),
            .I(N__6251));
    InMux I__1007 (
            .O(N__6270),
            .I(N__6248));
    Span4Mux_h I__1006 (
            .O(N__6267),
            .I(N__6234));
    LocalMux I__1005 (
            .O(N__6262),
            .I(N__6234));
    LocalMux I__1004 (
            .O(N__6257),
            .I(N__6234));
    LocalMux I__1003 (
            .O(N__6254),
            .I(N__6234));
    Span4Mux_v I__1002 (
            .O(N__6251),
            .I(N__6228));
    LocalMux I__1001 (
            .O(N__6248),
            .I(N__6228));
    InMux I__1000 (
            .O(N__6247),
            .I(N__6221));
    InMux I__999 (
            .O(N__6246),
            .I(N__6221));
    InMux I__998 (
            .O(N__6245),
            .I(N__6221));
    InMux I__997 (
            .O(N__6244),
            .I(N__6216));
    InMux I__996 (
            .O(N__6243),
            .I(N__6216));
    Span4Mux_v I__995 (
            .O(N__6234),
            .I(N__6213));
    InMux I__994 (
            .O(N__6233),
            .I(N__6210));
    Span4Mux_h I__993 (
            .O(N__6228),
            .I(N__6203));
    LocalMux I__992 (
            .O(N__6221),
            .I(N__6203));
    LocalMux I__991 (
            .O(N__6216),
            .I(N__6203));
    Sp12to4 I__990 (
            .O(N__6213),
            .I(N__6198));
    LocalMux I__989 (
            .O(N__6210),
            .I(N__6198));
    Span4Mux_v I__988 (
            .O(N__6203),
            .I(N__6195));
    Span12Mux_h I__987 (
            .O(N__6198),
            .I(N__6192));
    Span4Mux_h I__986 (
            .O(N__6195),
            .I(N__6189));
    Span12Mux_v I__985 (
            .O(N__6192),
            .I(N__6186));
    Sp12to4 I__984 (
            .O(N__6189),
            .I(N__6183));
    Odrv12 I__983 (
            .O(N__6186),
            .I(A_c_1));
    Odrv12 I__982 (
            .O(N__6183),
            .I(A_c_1));
    InMux I__981 (
            .O(N__6178),
            .I(N__6171));
    InMux I__980 (
            .O(N__6177),
            .I(N__6171));
    InMux I__979 (
            .O(N__6176),
            .I(N__6167));
    LocalMux I__978 (
            .O(N__6171),
            .I(N__6164));
    CascadeMux I__977 (
            .O(N__6170),
            .I(N__6161));
    LocalMux I__976 (
            .O(N__6167),
            .I(N__6155));
    Span4Mux_v I__975 (
            .O(N__6164),
            .I(N__6151));
    InMux I__974 (
            .O(N__6161),
            .I(N__6148));
    InMux I__973 (
            .O(N__6160),
            .I(N__6145));
    InMux I__972 (
            .O(N__6159),
            .I(N__6140));
    InMux I__971 (
            .O(N__6158),
            .I(N__6140));
    Span4Mux_h I__970 (
            .O(N__6155),
            .I(N__6137));
    InMux I__969 (
            .O(N__6154),
            .I(N__6134));
    Odrv4 I__968 (
            .O(N__6151),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__967 (
            .O(N__6148),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__966 (
            .O(N__6145),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__965 (
            .O(N__6140),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    Odrv4 I__964 (
            .O(N__6137),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__963 (
            .O(N__6134),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    InMux I__962 (
            .O(N__6121),
            .I(N__6115));
    InMux I__961 (
            .O(N__6120),
            .I(N__6115));
    LocalMux I__960 (
            .O(N__6115),
            .I(N__6112));
    Odrv4 I__959 (
            .O(N__6112),
            .I(\U409_AUTOCONFIG.un1_STATE_1_0 ));
    InMux I__958 (
            .O(N__6109),
            .I(N__6105));
    InMux I__957 (
            .O(N__6108),
            .I(N__6102));
    LocalMux I__956 (
            .O(N__6105),
            .I(N__6099));
    LocalMux I__955 (
            .O(N__6102),
            .I(N__6096));
    Odrv4 I__954 (
            .O(N__6099),
            .I(BRIDGE_BASE_0));
    Odrv4 I__953 (
            .O(N__6096),
            .I(BRIDGE_BASE_0));
    CascadeMux I__952 (
            .O(N__6091),
            .I(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_2_cascade_ ));
    InMux I__951 (
            .O(N__6088),
            .I(N__6082));
    InMux I__950 (
            .O(N__6087),
            .I(N__6082));
    LocalMux I__949 (
            .O(N__6082),
            .I(N__6078));
    InMux I__948 (
            .O(N__6081),
            .I(N__6075));
    Span4Mux_v I__947 (
            .O(N__6078),
            .I(N__6071));
    LocalMux I__946 (
            .O(N__6075),
            .I(N__6068));
    InMux I__945 (
            .O(N__6074),
            .I(N__6065));
    Span4Mux_v I__944 (
            .O(N__6071),
            .I(N__6062));
    Span4Mux_v I__943 (
            .O(N__6068),
            .I(N__6059));
    LocalMux I__942 (
            .O(N__6065),
            .I(N__6056));
    Span4Mux_h I__941 (
            .O(N__6062),
            .I(N__6053));
    Span4Mux_v I__940 (
            .O(N__6059),
            .I(N__6050));
    Sp12to4 I__939 (
            .O(N__6056),
            .I(N__6047));
    Sp12to4 I__938 (
            .O(N__6053),
            .I(N__6040));
    Sp12to4 I__937 (
            .O(N__6050),
            .I(N__6040));
    Span12Mux_v I__936 (
            .O(N__6047),
            .I(N__6040));
    Odrv12 I__935 (
            .O(N__6040),
            .I(A_c_26));
    CascadeMux I__934 (
            .O(N__6037),
            .I(N__6033));
    InMux I__933 (
            .O(N__6036),
            .I(N__6027));
    InMux I__932 (
            .O(N__6033),
            .I(N__6027));
    InMux I__931 (
            .O(N__6032),
            .I(N__6023));
    LocalMux I__930 (
            .O(N__6027),
            .I(N__6020));
    InMux I__929 (
            .O(N__6026),
            .I(N__6017));
    LocalMux I__928 (
            .O(N__6023),
            .I(N__6014));
    Span4Mux_v I__927 (
            .O(N__6020),
            .I(N__6011));
    LocalMux I__926 (
            .O(N__6017),
            .I(N__6008));
    Span4Mux_v I__925 (
            .O(N__6014),
            .I(N__6005));
    Span4Mux_h I__924 (
            .O(N__6011),
            .I(N__6000));
    Span4Mux_v I__923 (
            .O(N__6008),
            .I(N__6000));
    Sp12to4 I__922 (
            .O(N__6005),
            .I(N__5995));
    Sp12to4 I__921 (
            .O(N__6000),
            .I(N__5995));
    Odrv12 I__920 (
            .O(N__5995),
            .I(A_c_25));
    CascadeMux I__919 (
            .O(N__5992),
            .I(N__5988));
    InMux I__918 (
            .O(N__5991),
            .I(N__5984));
    InMux I__917 (
            .O(N__5988),
            .I(N__5979));
    InMux I__916 (
            .O(N__5987),
            .I(N__5979));
    LocalMux I__915 (
            .O(N__5984),
            .I(N__5975));
    LocalMux I__914 (
            .O(N__5979),
            .I(N__5972));
    InMux I__913 (
            .O(N__5978),
            .I(N__5969));
    Span4Mux_v I__912 (
            .O(N__5975),
            .I(N__5966));
    Span4Mux_h I__911 (
            .O(N__5972),
            .I(N__5963));
    LocalMux I__910 (
            .O(N__5969),
            .I(N__5960));
    Span4Mux_v I__909 (
            .O(N__5966),
            .I(N__5957));
    Sp12to4 I__908 (
            .O(N__5963),
            .I(N__5952));
    Sp12to4 I__907 (
            .O(N__5960),
            .I(N__5952));
    Sp12to4 I__906 (
            .O(N__5957),
            .I(N__5947));
    Span12Mux_v I__905 (
            .O(N__5952),
            .I(N__5947));
    Odrv12 I__904 (
            .O(N__5947),
            .I(A_c_24));
    InMux I__903 (
            .O(N__5944),
            .I(N__5941));
    LocalMux I__902 (
            .O(N__5941),
            .I(\U409_ADDRESS_DECODE.g2Z0Z_4 ));
    CascadeMux I__901 (
            .O(N__5938),
            .I(\U409_ADDRESS_DECODE.un1_Z2_SPACE_7Z0Z_1_cascade_ ));
    CascadeMux I__900 (
            .O(N__5935),
            .I(N__5931));
    InMux I__899 (
            .O(N__5934),
            .I(N__5928));
    InMux I__898 (
            .O(N__5931),
            .I(N__5925));
    LocalMux I__897 (
            .O(N__5928),
            .I(N__5917));
    LocalMux I__896 (
            .O(N__5925),
            .I(N__5917));
    InMux I__895 (
            .O(N__5924),
            .I(N__5914));
    InMux I__894 (
            .O(N__5923),
            .I(N__5911));
    InMux I__893 (
            .O(N__5922),
            .I(N__5908));
    Odrv4 I__892 (
            .O(N__5917),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__891 (
            .O(N__5914),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__890 (
            .O(N__5911),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__889 (
            .O(N__5908),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    InMux I__888 (
            .O(N__5899),
            .I(N__5895));
    InMux I__887 (
            .O(N__5898),
            .I(N__5892));
    LocalMux I__886 (
            .O(N__5895),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ));
    LocalMux I__885 (
            .O(N__5892),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ));
    CascadeMux I__884 (
            .O(N__5887),
            .I(N__5884));
    InMux I__883 (
            .O(N__5884),
            .I(N__5880));
    InMux I__882 (
            .O(N__5883),
            .I(N__5877));
    LocalMux I__881 (
            .O(N__5880),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ));
    LocalMux I__880 (
            .O(N__5877),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ));
    IoInMux I__879 (
            .O(N__5872),
            .I(N__5869));
    LocalMux I__878 (
            .O(N__5869),
            .I(N__5866));
    IoSpan4Mux I__877 (
            .O(N__5866),
            .I(N__5863));
    Span4Mux_s2_v I__876 (
            .O(N__5863),
            .I(N__5860));
    Sp12to4 I__875 (
            .O(N__5860),
            .I(N__5857));
    Span12Mux_s11_v I__874 (
            .O(N__5857),
            .I(N__5854));
    Odrv12 I__873 (
            .O(N__5854),
            .I(U409_AUTOCONFIG_D_OUT_0_i_2));
    CascadeMux I__872 (
            .O(N__5851),
            .I(N__5848));
    InMux I__871 (
            .O(N__5848),
            .I(N__5845));
    LocalMux I__870 (
            .O(N__5845),
            .I(N__5841));
    InMux I__869 (
            .O(N__5844),
            .I(N__5838));
    Odrv12 I__868 (
            .O(N__5841),
            .I(BRIDGE_BASE_1));
    LocalMux I__867 (
            .O(N__5838),
            .I(BRIDGE_BASE_1));
    InMux I__866 (
            .O(N__5833),
            .I(N__5830));
    LocalMux I__865 (
            .O(N__5830),
            .I(N__5826));
    InMux I__864 (
            .O(N__5829),
            .I(N__5823));
    Odrv12 I__863 (
            .O(N__5826),
            .I(BRIDGE_BASE_2));
    LocalMux I__862 (
            .O(N__5823),
            .I(BRIDGE_BASE_2));
    InMux I__861 (
            .O(N__5818),
            .I(N__5811));
    InMux I__860 (
            .O(N__5817),
            .I(N__5803));
    InMux I__859 (
            .O(N__5816),
            .I(N__5803));
    InMux I__858 (
            .O(N__5815),
            .I(N__5803));
    InMux I__857 (
            .O(N__5814),
            .I(N__5799));
    LocalMux I__856 (
            .O(N__5811),
            .I(N__5796));
    InMux I__855 (
            .O(N__5810),
            .I(N__5793));
    LocalMux I__854 (
            .O(N__5803),
            .I(N__5790));
    CascadeMux I__853 (
            .O(N__5802),
            .I(N__5785));
    LocalMux I__852 (
            .O(N__5799),
            .I(N__5782));
    Sp12to4 I__851 (
            .O(N__5796),
            .I(N__5777));
    LocalMux I__850 (
            .O(N__5793),
            .I(N__5777));
    Span4Mux_v I__849 (
            .O(N__5790),
            .I(N__5774));
    InMux I__848 (
            .O(N__5789),
            .I(N__5771));
    InMux I__847 (
            .O(N__5788),
            .I(N__5768));
    InMux I__846 (
            .O(N__5785),
            .I(N__5765));
    Span12Mux_v I__845 (
            .O(N__5782),
            .I(N__5762));
    Span12Mux_v I__844 (
            .O(N__5777),
            .I(N__5751));
    Sp12to4 I__843 (
            .O(N__5774),
            .I(N__5751));
    LocalMux I__842 (
            .O(N__5771),
            .I(N__5751));
    LocalMux I__841 (
            .O(N__5768),
            .I(N__5751));
    LocalMux I__840 (
            .O(N__5765),
            .I(N__5751));
    Odrv12 I__839 (
            .O(N__5762),
            .I(A_c_5));
    Odrv12 I__838 (
            .O(N__5751),
            .I(A_c_5));
    CascadeMux I__837 (
            .O(N__5746),
            .I(N__5742));
    InMux I__836 (
            .O(N__5745),
            .I(N__5737));
    InMux I__835 (
            .O(N__5742),
            .I(N__5737));
    LocalMux I__834 (
            .O(N__5737),
            .I(\U409_AUTOCONFIG.N_68 ));
    CascadeMux I__833 (
            .O(N__5734),
            .I(N__5730));
    InMux I__832 (
            .O(N__5733),
            .I(N__5724));
    InMux I__831 (
            .O(N__5730),
            .I(N__5721));
    InMux I__830 (
            .O(N__5729),
            .I(N__5716));
    InMux I__829 (
            .O(N__5728),
            .I(N__5716));
    InMux I__828 (
            .O(N__5727),
            .I(N__5713));
    LocalMux I__827 (
            .O(N__5724),
            .I(N__5709));
    LocalMux I__826 (
            .O(N__5721),
            .I(N__5704));
    LocalMux I__825 (
            .O(N__5716),
            .I(N__5704));
    LocalMux I__824 (
            .O(N__5713),
            .I(N__5698));
    CascadeMux I__823 (
            .O(N__5712),
            .I(N__5690));
    Span4Mux_v I__822 (
            .O(N__5709),
            .I(N__5685));
    Span4Mux_v I__821 (
            .O(N__5704),
            .I(N__5685));
    InMux I__820 (
            .O(N__5703),
            .I(N__5680));
    InMux I__819 (
            .O(N__5702),
            .I(N__5680));
    InMux I__818 (
            .O(N__5701),
            .I(N__5677));
    Span4Mux_v I__817 (
            .O(N__5698),
            .I(N__5674));
    InMux I__816 (
            .O(N__5697),
            .I(N__5667));
    InMux I__815 (
            .O(N__5696),
            .I(N__5667));
    InMux I__814 (
            .O(N__5695),
            .I(N__5667));
    InMux I__813 (
            .O(N__5694),
            .I(N__5664));
    InMux I__812 (
            .O(N__5693),
            .I(N__5659));
    InMux I__811 (
            .O(N__5690),
            .I(N__5659));
    Sp12to4 I__810 (
            .O(N__5685),
            .I(N__5644));
    LocalMux I__809 (
            .O(N__5680),
            .I(N__5644));
    LocalMux I__808 (
            .O(N__5677),
            .I(N__5644));
    Sp12to4 I__807 (
            .O(N__5674),
            .I(N__5644));
    LocalMux I__806 (
            .O(N__5667),
            .I(N__5644));
    LocalMux I__805 (
            .O(N__5664),
            .I(N__5644));
    LocalMux I__804 (
            .O(N__5659),
            .I(N__5644));
    Odrv12 I__803 (
            .O(N__5644),
            .I(A_c_4));
    InMux I__802 (
            .O(N__5641),
            .I(N__5638));
    LocalMux I__801 (
            .O(N__5638),
            .I(\U409_AUTOCONFIG.N_47 ));
    InMux I__800 (
            .O(N__5635),
            .I(N__5632));
    LocalMux I__799 (
            .O(N__5632),
            .I(N__5629));
    Span4Mux_v I__798 (
            .O(N__5629),
            .I(N__5626));
    Sp12to4 I__797 (
            .O(N__5626),
            .I(N__5623));
    Span12Mux_h I__796 (
            .O(N__5623),
            .I(N__5620));
    Span12Mux_h I__795 (
            .O(N__5620),
            .I(N__5617));
    Span12Mux_v I__794 (
            .O(N__5617),
            .I(N__5614));
    Odrv12 I__793 (
            .O(N__5614),
            .I(AUTOBOOT_c));
    InMux I__792 (
            .O(N__5611),
            .I(N__5607));
    InMux I__791 (
            .O(N__5610),
            .I(N__5604));
    LocalMux I__790 (
            .O(N__5607),
            .I(N__5601));
    LocalMux I__789 (
            .O(N__5604),
            .I(N__5598));
    Span4Mux_v I__788 (
            .O(N__5601),
            .I(N__5594));
    Span4Mux_v I__787 (
            .O(N__5598),
            .I(N__5591));
    InMux I__786 (
            .O(N__5597),
            .I(N__5588));
    Odrv4 I__785 (
            .O(N__5594),
            .I(\U409_AUTOCONFIG.N_196_1 ));
    Odrv4 I__784 (
            .O(N__5591),
            .I(\U409_AUTOCONFIG.N_196_1 ));
    LocalMux I__783 (
            .O(N__5588),
            .I(\U409_AUTOCONFIG.N_196_1 ));
    InMux I__782 (
            .O(N__5581),
            .I(N__5570));
    InMux I__781 (
            .O(N__5580),
            .I(N__5570));
    InMux I__780 (
            .O(N__5579),
            .I(N__5565));
    InMux I__779 (
            .O(N__5578),
            .I(N__5565));
    InMux I__778 (
            .O(N__5577),
            .I(N__5561));
    CascadeMux I__777 (
            .O(N__5576),
            .I(N__5556));
    CascadeMux I__776 (
            .O(N__5575),
            .I(N__5552));
    LocalMux I__775 (
            .O(N__5570),
            .I(N__5547));
    LocalMux I__774 (
            .O(N__5565),
            .I(N__5547));
    InMux I__773 (
            .O(N__5564),
            .I(N__5544));
    LocalMux I__772 (
            .O(N__5561),
            .I(N__5537));
    InMux I__771 (
            .O(N__5560),
            .I(N__5534));
    InMux I__770 (
            .O(N__5559),
            .I(N__5531));
    InMux I__769 (
            .O(N__5556),
            .I(N__5526));
    InMux I__768 (
            .O(N__5555),
            .I(N__5526));
    InMux I__767 (
            .O(N__5552),
            .I(N__5523));
    Span4Mux_h I__766 (
            .O(N__5547),
            .I(N__5518));
    LocalMux I__765 (
            .O(N__5544),
            .I(N__5518));
    InMux I__764 (
            .O(N__5543),
            .I(N__5513));
    InMux I__763 (
            .O(N__5542),
            .I(N__5513));
    InMux I__762 (
            .O(N__5541),
            .I(N__5508));
    InMux I__761 (
            .O(N__5540),
            .I(N__5508));
    Span4Mux_v I__760 (
            .O(N__5537),
            .I(N__5501));
    LocalMux I__759 (
            .O(N__5534),
            .I(N__5501));
    LocalMux I__758 (
            .O(N__5531),
            .I(N__5501));
    LocalMux I__757 (
            .O(N__5526),
            .I(N__5498));
    LocalMux I__756 (
            .O(N__5523),
            .I(N__5495));
    Span4Mux_h I__755 (
            .O(N__5518),
            .I(N__5488));
    LocalMux I__754 (
            .O(N__5513),
            .I(N__5488));
    LocalMux I__753 (
            .O(N__5508),
            .I(N__5488));
    Span4Mux_v I__752 (
            .O(N__5501),
            .I(N__5485));
    Span4Mux_v I__751 (
            .O(N__5498),
            .I(N__5478));
    Span4Mux_v I__750 (
            .O(N__5495),
            .I(N__5478));
    Span4Mux_v I__749 (
            .O(N__5488),
            .I(N__5478));
    Sp12to4 I__748 (
            .O(N__5485),
            .I(N__5473));
    Sp12to4 I__747 (
            .O(N__5478),
            .I(N__5473));
    Span12Mux_h I__746 (
            .O(N__5473),
            .I(N__5470));
    Odrv12 I__745 (
            .O(N__5470),
            .I(A_c_2));
    InMux I__744 (
            .O(N__5467),
            .I(N__5459));
    InMux I__743 (
            .O(N__5466),
            .I(N__5459));
    InMux I__742 (
            .O(N__5465),
            .I(N__5456));
    CascadeMux I__741 (
            .O(N__5464),
            .I(N__5452));
    LocalMux I__740 (
            .O(N__5459),
            .I(N__5445));
    LocalMux I__739 (
            .O(N__5456),
            .I(N__5442));
    InMux I__738 (
            .O(N__5455),
            .I(N__5437));
    InMux I__737 (
            .O(N__5452),
            .I(N__5437));
    CascadeMux I__736 (
            .O(N__5451),
            .I(N__5434));
    InMux I__735 (
            .O(N__5450),
            .I(N__5428));
    InMux I__734 (
            .O(N__5449),
            .I(N__5425));
    InMux I__733 (
            .O(N__5448),
            .I(N__5422));
    Span4Mux_v I__732 (
            .O(N__5445),
            .I(N__5419));
    Span4Mux_v I__731 (
            .O(N__5442),
            .I(N__5414));
    LocalMux I__730 (
            .O(N__5437),
            .I(N__5414));
    InMux I__729 (
            .O(N__5434),
            .I(N__5409));
    InMux I__728 (
            .O(N__5433),
            .I(N__5409));
    InMux I__727 (
            .O(N__5432),
            .I(N__5406));
    InMux I__726 (
            .O(N__5431),
            .I(N__5403));
    LocalMux I__725 (
            .O(N__5428),
            .I(N__5400));
    LocalMux I__724 (
            .O(N__5425),
            .I(N__5387));
    LocalMux I__723 (
            .O(N__5422),
            .I(N__5387));
    Sp12to4 I__722 (
            .O(N__5419),
            .I(N__5387));
    Sp12to4 I__721 (
            .O(N__5414),
            .I(N__5387));
    LocalMux I__720 (
            .O(N__5409),
            .I(N__5387));
    LocalMux I__719 (
            .O(N__5406),
            .I(N__5387));
    LocalMux I__718 (
            .O(N__5403),
            .I(N__5384));
    Sp12to4 I__717 (
            .O(N__5400),
            .I(N__5381));
    Span12Mux_h I__716 (
            .O(N__5387),
            .I(N__5378));
    Span12Mux_v I__715 (
            .O(N__5384),
            .I(N__5375));
    Span12Mux_v I__714 (
            .O(N__5381),
            .I(N__5372));
    Span12Mux_v I__713 (
            .O(N__5378),
            .I(N__5369));
    Odrv12 I__712 (
            .O(N__5375),
            .I(A_c_3));
    Odrv12 I__711 (
            .O(N__5372),
            .I(A_c_3));
    Odrv12 I__710 (
            .O(N__5369),
            .I(A_c_3));
    CascadeMux I__709 (
            .O(N__5362),
            .I(N__5359));
    InMux I__708 (
            .O(N__5359),
            .I(N__5356));
    LocalMux I__707 (
            .O(N__5356),
            .I(N__5353));
    Odrv4 I__706 (
            .O(N__5353),
            .I(\U409_AUTOCONFIG.N_54 ));
    InMux I__705 (
            .O(N__5350),
            .I(N__5347));
    LocalMux I__704 (
            .O(N__5347),
            .I(\U409_ADDRESS_DECODE.g2_5_0 ));
    CascadeMux I__703 (
            .O(N__5344),
            .I(\U409_ADDRESS_DECODE.g2_6_0_cascade_ ));
    InMux I__702 (
            .O(N__5341),
            .I(N__5335));
    InMux I__701 (
            .O(N__5340),
            .I(N__5329));
    InMux I__700 (
            .O(N__5339),
            .I(N__5329));
    InMux I__699 (
            .O(N__5338),
            .I(N__5326));
    LocalMux I__698 (
            .O(N__5335),
            .I(N__5323));
    InMux I__697 (
            .O(N__5334),
            .I(N__5320));
    LocalMux I__696 (
            .O(N__5329),
            .I(N__5315));
    LocalMux I__695 (
            .O(N__5326),
            .I(N__5315));
    Span4Mux_v I__694 (
            .O(N__5323),
            .I(N__5312));
    LocalMux I__693 (
            .O(N__5320),
            .I(N__5307));
    Sp12to4 I__692 (
            .O(N__5315),
            .I(N__5307));
    Span4Mux_v I__691 (
            .O(N__5312),
            .I(N__5304));
    Span12Mux_v I__690 (
            .O(N__5307),
            .I(N__5301));
    Span4Mux_h I__689 (
            .O(N__5304),
            .I(N__5298));
    Odrv12 I__688 (
            .O(N__5301),
            .I(A_c_29));
    Odrv4 I__687 (
            .O(N__5298),
            .I(A_c_29));
    CascadeMux I__686 (
            .O(N__5293),
            .I(N__5288));
    InMux I__685 (
            .O(N__5292),
            .I(N__5283));
    InMux I__684 (
            .O(N__5291),
            .I(N__5283));
    InMux I__683 (
            .O(N__5288),
            .I(N__5280));
    LocalMux I__682 (
            .O(N__5283),
            .I(N__5275));
    LocalMux I__681 (
            .O(N__5280),
            .I(N__5272));
    InMux I__680 (
            .O(N__5279),
            .I(N__5269));
    InMux I__679 (
            .O(N__5278),
            .I(N__5266));
    Span4Mux_h I__678 (
            .O(N__5275),
            .I(N__5259));
    Span4Mux_h I__677 (
            .O(N__5272),
            .I(N__5259));
    LocalMux I__676 (
            .O(N__5269),
            .I(N__5259));
    LocalMux I__675 (
            .O(N__5266),
            .I(N__5256));
    Span4Mux_h I__674 (
            .O(N__5259),
            .I(N__5253));
    Span12Mux_v I__673 (
            .O(N__5256),
            .I(N__5250));
    Span4Mux_v I__672 (
            .O(N__5253),
            .I(N__5247));
    Odrv12 I__671 (
            .O(N__5250),
            .I(A_c_30));
    Odrv4 I__670 (
            .O(N__5247),
            .I(A_c_30));
    CascadeMux I__669 (
            .O(N__5242),
            .I(N__5236));
    InMux I__668 (
            .O(N__5241),
            .I(N__5231));
    InMux I__667 (
            .O(N__5240),
            .I(N__5231));
    InMux I__666 (
            .O(N__5239),
            .I(N__5228));
    InMux I__665 (
            .O(N__5236),
            .I(N__5225));
    LocalMux I__664 (
            .O(N__5231),
            .I(N__5222));
    LocalMux I__663 (
            .O(N__5228),
            .I(N__5219));
    LocalMux I__662 (
            .O(N__5225),
            .I(N__5216));
    Span4Mux_v I__661 (
            .O(N__5222),
            .I(N__5213));
    Span4Mux_v I__660 (
            .O(N__5219),
            .I(N__5210));
    Span4Mux_v I__659 (
            .O(N__5216),
            .I(N__5207));
    Sp12to4 I__658 (
            .O(N__5213),
            .I(N__5202));
    Sp12to4 I__657 (
            .O(N__5210),
            .I(N__5202));
    Sp12to4 I__656 (
            .O(N__5207),
            .I(N__5199));
    Odrv12 I__655 (
            .O(N__5202),
            .I(A_c_27));
    Odrv12 I__654 (
            .O(N__5199),
            .I(A_c_27));
    InMux I__653 (
            .O(N__5194),
            .I(N__5191));
    LocalMux I__652 (
            .O(N__5191),
            .I(\U409_ADDRESS_DECODE.g0_i_a4_1Z0Z_3 ));
    InMux I__651 (
            .O(N__5188),
            .I(N__5185));
    LocalMux I__650 (
            .O(N__5185),
            .I(\U409_ADDRESS_DECODE.g0_i_a4Z0Z_1 ));
    InMux I__649 (
            .O(N__5182),
            .I(N__5178));
    InMux I__648 (
            .O(N__5181),
            .I(N__5175));
    LocalMux I__647 (
            .O(N__5178),
            .I(\U409_AUTOCONFIG.AC_STARTZ0 ));
    LocalMux I__646 (
            .O(N__5175),
            .I(\U409_AUTOCONFIG.AC_STARTZ0 ));
    InMux I__645 (
            .O(N__5170),
            .I(N__5167));
    LocalMux I__644 (
            .O(N__5167),
            .I(N__5164));
    Span4Mux_h I__643 (
            .O(N__5164),
            .I(N__5161));
    Odrv4 I__642 (
            .O(N__5161),
            .I(\U409_AUTOCONFIG.LIDE_OUTc_0_0 ));
    CascadeMux I__641 (
            .O(N__5158),
            .I(N__5155));
    InMux I__640 (
            .O(N__5155),
            .I(N__5152));
    LocalMux I__639 (
            .O(N__5152),
            .I(N__5148));
    InMux I__638 (
            .O(N__5151),
            .I(N__5145));
    Odrv12 I__637 (
            .O(N__5148),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ1Z_0 ));
    LocalMux I__636 (
            .O(N__5145),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ1Z_0 ));
    InMux I__635 (
            .O(N__5140),
            .I(N__5137));
    LocalMux I__634 (
            .O(N__5137),
            .I(\U409_AUTOCONFIG.N_50 ));
    CascadeMux I__633 (
            .O(N__5134),
            .I(N__5131));
    InMux I__632 (
            .O(N__5131),
            .I(N__5128));
    LocalMux I__631 (
            .O(N__5128),
            .I(N__5125));
    Odrv4 I__630 (
            .O(N__5125),
            .I(\U409_AUTOCONFIG.LIDE_OUTc_0_0_0 ));
    InMux I__629 (
            .O(N__5122),
            .I(N__5119));
    LocalMux I__628 (
            .O(N__5119),
            .I(N__5116));
    Span4Mux_v I__627 (
            .O(N__5116),
            .I(N__5112));
    InMux I__626 (
            .O(N__5115),
            .I(N__5109));
    Odrv4 I__625 (
            .O(N__5112),
            .I(\U409_AUTOCONFIG.N_48 ));
    LocalMux I__624 (
            .O(N__5109),
            .I(\U409_AUTOCONFIG.N_48 ));
    InMux I__623 (
            .O(N__5104),
            .I(N__5092));
    InMux I__622 (
            .O(N__5103),
            .I(N__5092));
    InMux I__621 (
            .O(N__5102),
            .I(N__5092));
    InMux I__620 (
            .O(N__5101),
            .I(N__5092));
    LocalMux I__619 (
            .O(N__5092),
            .I(\U409_AUTOCONFIG.AC_START_RNI777KZ0Z2 ));
    InMux I__618 (
            .O(N__5089),
            .I(N__5085));
    CascadeMux I__617 (
            .O(N__5088),
            .I(N__5082));
    LocalMux I__616 (
            .O(N__5085),
            .I(N__5079));
    InMux I__615 (
            .O(N__5082),
            .I(N__5076));
    Odrv4 I__614 (
            .O(N__5079),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ));
    LocalMux I__613 (
            .O(N__5076),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ));
    InMux I__612 (
            .O(N__5071),
            .I(N__5065));
    InMux I__611 (
            .O(N__5070),
            .I(N__5065));
    LocalMux I__610 (
            .O(N__5065),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ));
    InMux I__609 (
            .O(N__5062),
            .I(N__5058));
    InMux I__608 (
            .O(N__5061),
            .I(N__5055));
    LocalMux I__607 (
            .O(N__5058),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ1Z_1 ));
    LocalMux I__606 (
            .O(N__5055),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ1Z_1 ));
    IoInMux I__605 (
            .O(N__5050),
            .I(N__5047));
    LocalMux I__604 (
            .O(N__5047),
            .I(N__5044));
    Span12Mux_s4_v I__603 (
            .O(N__5044),
            .I(N__5041));
    Span12Mux_v I__602 (
            .O(N__5041),
            .I(N__5038));
    Odrv12 I__601 (
            .O(N__5038),
            .I(U409_AUTOCONFIG_D_OUT_0_i_1));
    InMux I__600 (
            .O(N__5035),
            .I(N__5032));
    LocalMux I__599 (
            .O(N__5032),
            .I(N__5028));
    InMux I__598 (
            .O(N__5031),
            .I(N__5025));
    Odrv4 I__597 (
            .O(N__5028),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ));
    LocalMux I__596 (
            .O(N__5025),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ));
    IoInMux I__595 (
            .O(N__5020),
            .I(N__5017));
    LocalMux I__594 (
            .O(N__5017),
            .I(N__5014));
    Span4Mux_s3_v I__593 (
            .O(N__5014),
            .I(N__5011));
    Span4Mux_v I__592 (
            .O(N__5011),
            .I(N__5008));
    Span4Mux_v I__591 (
            .O(N__5008),
            .I(N__5005));
    Odrv4 I__590 (
            .O(N__5005),
            .I(U409_AUTOCONFIG_D_OUT_0_i_0));
    CascadeMux I__589 (
            .O(N__5002),
            .I(\U409_TRANSFER_ACK.G_14_0_a7_1_3_cascade_ ));
    InMux I__588 (
            .O(N__4999),
            .I(N__4994));
    InMux I__587 (
            .O(N__4998),
            .I(N__4991));
    InMux I__586 (
            .O(N__4997),
            .I(N__4988));
    LocalMux I__585 (
            .O(N__4994),
            .I(N__4981));
    LocalMux I__584 (
            .O(N__4991),
            .I(N__4981));
    LocalMux I__583 (
            .O(N__4988),
            .I(N__4981));
    Span4Mux_v I__582 (
            .O(N__4981),
            .I(N__4978));
    Odrv4 I__581 (
            .O(N__4978),
            .I(\U409_AUTOCONFIG.un1_AZ0Z_18 ));
    InMux I__580 (
            .O(N__4975),
            .I(N__4968));
    InMux I__579 (
            .O(N__4974),
            .I(N__4968));
    InMux I__578 (
            .O(N__4973),
            .I(N__4962));
    LocalMux I__577 (
            .O(N__4968),
            .I(N__4959));
    InMux I__576 (
            .O(N__4967),
            .I(N__4956));
    InMux I__575 (
            .O(N__4966),
            .I(N__4953));
    InMux I__574 (
            .O(N__4965),
            .I(N__4950));
    LocalMux I__573 (
            .O(N__4962),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    Odrv4 I__572 (
            .O(N__4959),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__571 (
            .O(N__4956),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__570 (
            .O(N__4953),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__569 (
            .O(N__4950),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    CascadeMux I__568 (
            .O(N__4939),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7_cascade_ ));
    InMux I__567 (
            .O(N__4936),
            .I(N__4933));
    LocalMux I__566 (
            .O(N__4933),
            .I(N__4930));
    Odrv4 I__565 (
            .O(N__4930),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_4 ));
    InMux I__564 (
            .O(N__4927),
            .I(N__4924));
    LocalMux I__563 (
            .O(N__4924),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_10 ));
    CascadeMux I__562 (
            .O(N__4921),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9_cascade_ ));
    InMux I__561 (
            .O(N__4918),
            .I(N__4915));
    LocalMux I__560 (
            .O(N__4915),
            .I(N__4912));
    Span4Mux_v I__559 (
            .O(N__4912),
            .I(N__4909));
    Span4Mux_v I__558 (
            .O(N__4909),
            .I(N__4906));
    IoSpan4Mux I__557 (
            .O(N__4906),
            .I(N__4903));
    Odrv4 I__556 (
            .O(N__4903),
            .I(TT_c_1));
    CascadeMux I__555 (
            .O(N__4900),
            .I(N__4897));
    InMux I__554 (
            .O(N__4897),
            .I(N__4894));
    LocalMux I__553 (
            .O(N__4894),
            .I(N__4891));
    Span4Mux_h I__552 (
            .O(N__4891),
            .I(N__4888));
    Span4Mux_v I__551 (
            .O(N__4888),
            .I(N__4885));
    Span4Mux_v I__550 (
            .O(N__4885),
            .I(N__4882));
    Odrv4 I__549 (
            .O(N__4882),
            .I(TT_c_0));
    InMux I__548 (
            .O(N__4879),
            .I(N__4876));
    LocalMux I__547 (
            .O(N__4876),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8 ));
    InMux I__546 (
            .O(N__4873),
            .I(N__4870));
    LocalMux I__545 (
            .O(N__4870),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3 ));
    CascadeMux I__544 (
            .O(N__4867),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4_cascade_ ));
    CascadeMux I__543 (
            .O(N__4864),
            .I(AUTOCONFIG_SPACE_cascade_));
    IoInMux I__542 (
            .O(N__4861),
            .I(N__4858));
    LocalMux I__541 (
            .O(N__4858),
            .I(N__4853));
    IoInMux I__540 (
            .O(N__4857),
            .I(N__4850));
    IoInMux I__539 (
            .O(N__4856),
            .I(N__4847));
    IoSpan4Mux I__538 (
            .O(N__4853),
            .I(N__4839));
    LocalMux I__537 (
            .O(N__4850),
            .I(N__4839));
    LocalMux I__536 (
            .O(N__4847),
            .I(N__4839));
    IoInMux I__535 (
            .O(N__4846),
            .I(N__4836));
    IoSpan4Mux I__534 (
            .O(N__4839),
            .I(N__4831));
    LocalMux I__533 (
            .O(N__4836),
            .I(N__4831));
    Span4Mux_s3_v I__532 (
            .O(N__4831),
            .I(N__4828));
    Span4Mux_v I__531 (
            .O(N__4828),
            .I(N__4825));
    Span4Mux_v I__530 (
            .O(N__4825),
            .I(N__4822));
    Odrv4 I__529 (
            .O(N__4822),
            .I(D_1_i));
    InMux I__528 (
            .O(N__4819),
            .I(N__4816));
    LocalMux I__527 (
            .O(N__4816),
            .I(N__4813));
    Odrv12 I__526 (
            .O(N__4813),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0 ));
    CascadeMux I__525 (
            .O(N__4810),
            .I(N__4807));
    InMux I__524 (
            .O(N__4807),
            .I(N__4804));
    LocalMux I__523 (
            .O(N__4804),
            .I(N__4801));
    Odrv4 I__522 (
            .O(N__4801),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_1_0 ));
    InMux I__521 (
            .O(N__4798),
            .I(N__4791));
    InMux I__520 (
            .O(N__4797),
            .I(N__4791));
    InMux I__519 (
            .O(N__4796),
            .I(N__4788));
    LocalMux I__518 (
            .O(N__4791),
            .I(\U409_AUTOCONFIG.N_59_1 ));
    LocalMux I__517 (
            .O(N__4788),
            .I(\U409_AUTOCONFIG.N_59_1 ));
    InMux I__516 (
            .O(N__4783),
            .I(N__4780));
    LocalMux I__515 (
            .O(N__4780),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_8_sqmuxa ));
    InMux I__514 (
            .O(N__4777),
            .I(N__4774));
    LocalMux I__513 (
            .O(N__4774),
            .I(N__4771));
    Span4Mux_v I__512 (
            .O(N__4771),
            .I(N__4767));
    InMux I__511 (
            .O(N__4770),
            .I(N__4764));
    Sp12to4 I__510 (
            .O(N__4767),
            .I(N__4759));
    LocalMux I__509 (
            .O(N__4764),
            .I(N__4759));
    Odrv12 I__508 (
            .O(N__4759),
            .I(\U409_AUTOCONFIG.N_57 ));
    InMux I__507 (
            .O(N__4756),
            .I(N__4753));
    LocalMux I__506 (
            .O(N__4753),
            .I(N__4750));
    Span4Mux_h I__505 (
            .O(N__4750),
            .I(N__4747));
    Odrv4 I__504 (
            .O(N__4747),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_1 ));
    CascadeMux I__503 (
            .O(N__4744),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_8_sqmuxa_cascade_ ));
    CascadeMux I__502 (
            .O(N__4741),
            .I(\U409_AUTOCONFIG.LIDE_OUT_7_94_i_i_1_tz_cascade_ ));
    CascadeMux I__501 (
            .O(N__4738),
            .I(\U409_ADDRESS_DECODE.g0_i_a4_0Z0Z_2_cascade_ ));
    CascadeMux I__500 (
            .O(N__4735),
            .I(\U409_AUTOCONFIG.N_55_cascade_ ));
    InMux I__499 (
            .O(N__4732),
            .I(N__4729));
    LocalMux I__498 (
            .O(N__4729),
            .I(N__4725));
    InMux I__497 (
            .O(N__4728),
            .I(N__4722));
    Odrv4 I__496 (
            .O(N__4725),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ));
    LocalMux I__495 (
            .O(N__4722),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ));
    CascadeMux I__494 (
            .O(N__4717),
            .I(N__4714));
    InMux I__493 (
            .O(N__4714),
            .I(N__4710));
    CascadeMux I__492 (
            .O(N__4713),
            .I(N__4707));
    LocalMux I__491 (
            .O(N__4710),
            .I(N__4704));
    InMux I__490 (
            .O(N__4707),
            .I(N__4701));
    Span4Mux_v I__489 (
            .O(N__4704),
            .I(N__4698));
    LocalMux I__488 (
            .O(N__4701),
            .I(N__4695));
    Sp12to4 I__487 (
            .O(N__4698),
            .I(N__4692));
    Span4Mux_h I__486 (
            .O(N__4695),
            .I(N__4689));
    Span12Mux_s10_h I__485 (
            .O(N__4692),
            .I(N__4684));
    Sp12to4 I__484 (
            .O(N__4689),
            .I(N__4684));
    Span12Mux_v I__483 (
            .O(N__4684),
            .I(N__4681));
    Odrv12 I__482 (
            .O(N__4681),
            .I(CPUCONFn_c));
    InMux I__481 (
            .O(N__4678),
            .I(N__4675));
    LocalMux I__480 (
            .O(N__4675),
            .I(N__4672));
    Span4Mux_v I__479 (
            .O(N__4672),
            .I(N__4669));
    Odrv4 I__478 (
            .O(N__4669),
            .I(\U409_AUTOCONFIG.N_40 ));
    CascadeMux I__477 (
            .O(N__4666),
            .I(\U409_AUTOCONFIG.N_59_1_cascade_ ));
    InMux I__476 (
            .O(N__4663),
            .I(N__4660));
    LocalMux I__475 (
            .O(N__4660),
            .I(N__4656));
    InMux I__474 (
            .O(N__4659),
            .I(N__4653));
    Odrv12 I__473 (
            .O(N__4656),
            .I(\U409_AUTOCONFIG.N_61 ));
    LocalMux I__472 (
            .O(N__4653),
            .I(\U409_AUTOCONFIG.N_61 ));
    CascadeMux I__471 (
            .O(N__4648),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_2_cascade_ ));
    InMux I__470 (
            .O(N__4645),
            .I(N__4639));
    InMux I__469 (
            .O(N__4644),
            .I(N__4639));
    LocalMux I__468 (
            .O(N__4639),
            .I(N__4636));
    Odrv4 I__467 (
            .O(N__4636),
            .I(\U409_AUTOCONFIG.N_67 ));
    InMux I__466 (
            .O(N__4633),
            .I(N__4630));
    LocalMux I__465 (
            .O(N__4630),
            .I(\U409_AUTOCONFIG.N_56 ));
    InMux I__464 (
            .O(N__4627),
            .I(N__4624));
    LocalMux I__463 (
            .O(N__4624),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ));
    CascadeMux I__462 (
            .O(N__4621),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5_cascade_ ));
    InMux I__461 (
            .O(N__4618),
            .I(N__4615));
    LocalMux I__460 (
            .O(N__4615),
            .I(N__4612));
    Span4Mux_h I__459 (
            .O(N__4612),
            .I(N__4609));
    Odrv4 I__458 (
            .O(N__4609),
            .I(\U409_AUTOCONFIG.ATA_BASE10Z0Z_2 ));
    CascadeMux I__457 (
            .O(N__4606),
            .I(\U409_AUTOCONFIG.ATA_BASE10_cascade_ ));
    IoInMux I__456 (
            .O(N__4603),
            .I(N__4600));
    LocalMux I__455 (
            .O(N__4600),
            .I(N__4597));
    Span12Mux_s2_v I__454 (
            .O(N__4597),
            .I(N__4594));
    Span12Mux_v I__453 (
            .O(N__4594),
            .I(N__4591));
    Odrv12 I__452 (
            .O(N__4591),
            .I(U409_AUTOCONFIG_D_OUT_0_i_3));
    InMux I__451 (
            .O(N__4588),
            .I(N__4585));
    LocalMux I__450 (
            .O(N__4585),
            .I(N__4580));
    CascadeMux I__449 (
            .O(N__4584),
            .I(N__4577));
    CascadeMux I__448 (
            .O(N__4583),
            .I(N__4573));
    Span4Mux_v I__447 (
            .O(N__4580),
            .I(N__4568));
    InMux I__446 (
            .O(N__4577),
            .I(N__4559));
    InMux I__445 (
            .O(N__4576),
            .I(N__4559));
    InMux I__444 (
            .O(N__4573),
            .I(N__4559));
    InMux I__443 (
            .O(N__4572),
            .I(N__4559));
    InMux I__442 (
            .O(N__4571),
            .I(N__4556));
    Sp12to4 I__441 (
            .O(N__4568),
            .I(N__4549));
    LocalMux I__440 (
            .O(N__4559),
            .I(N__4549));
    LocalMux I__439 (
            .O(N__4556),
            .I(N__4549));
    Odrv12 I__438 (
            .O(N__4549),
            .I(A_c_6));
    InMux I__437 (
            .O(N__4546),
            .I(N__4534));
    InMux I__436 (
            .O(N__4545),
            .I(N__4534));
    InMux I__435 (
            .O(N__4544),
            .I(N__4534));
    InMux I__434 (
            .O(N__4543),
            .I(N__4534));
    LocalMux I__433 (
            .O(N__4534),
            .I(N__4529));
    InMux I__432 (
            .O(N__4533),
            .I(N__4526));
    InMux I__431 (
            .O(N__4532),
            .I(N__4523));
    Span4Mux_v I__430 (
            .O(N__4529),
            .I(N__4520));
    LocalMux I__429 (
            .O(N__4526),
            .I(N__4515));
    LocalMux I__428 (
            .O(N__4523),
            .I(N__4515));
    Sp12to4 I__427 (
            .O(N__4520),
            .I(N__4510));
    Span12Mux_v I__426 (
            .O(N__4515),
            .I(N__4510));
    Odrv12 I__425 (
            .O(N__4510),
            .I(A_c_7));
    CascadeMux I__424 (
            .O(N__4507),
            .I(\U409_AUTOCONFIG.un1_A_18Z0Z_0_cascade_ ));
    CascadeMux I__423 (
            .O(N__4504),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_cascade_ ));
    InMux I__422 (
            .O(N__4501),
            .I(N__4498));
    LocalMux I__421 (
            .O(N__4498),
            .I(\U409_AUTOCONFIG.N_63 ));
    CascadeMux I__420 (
            .O(N__4495),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_1_2_0_cascade_ ));
    CascadeMux I__419 (
            .O(N__4492),
            .I(\U409_AUTOCONFIG.N_196_1_cascade_ ));
    InMux I__418 (
            .O(N__4489),
            .I(N__4486));
    LocalMux I__417 (
            .O(N__4486),
            .I(\U409_AUTOCONFIG.LIDE_OUT_7_0_62_i_i_a3_0 ));
    CascadeMux I__416 (
            .O(N__4483),
            .I(\U409_AUTOCONFIG.N_67_cascade_ ));
    CascadeMux I__415 (
            .O(N__4480),
            .I(N__4476));
    InMux I__414 (
            .O(N__4479),
            .I(N__4473));
    InMux I__413 (
            .O(N__4476),
            .I(N__4470));
    LocalMux I__412 (
            .O(N__4473),
            .I(\U409_AUTOCONFIG.N_214_1 ));
    LocalMux I__411 (
            .O(N__4470),
            .I(\U409_AUTOCONFIG.N_214_1 ));
    IoInMux I__410 (
            .O(N__4465),
            .I(N__4462));
    LocalMux I__409 (
            .O(N__4462),
            .I(N__4459));
    Span4Mux_s2_h I__408 (
            .O(N__4459),
            .I(N__4456));
    Sp12to4 I__407 (
            .O(N__4456),
            .I(N__4453));
    Span12Mux_v I__406 (
            .O(N__4453),
            .I(N__4450));
    Span12Mux_v I__405 (
            .O(N__4450),
            .I(N__4447));
    Odrv12 I__404 (
            .O(N__4447),
            .I(PIO_P0_c));
    IoInMux I__403 (
            .O(N__4444),
            .I(N__4441));
    LocalMux I__402 (
            .O(N__4441),
            .I(N__4438));
    IoSpan4Mux I__401 (
            .O(N__4438),
            .I(N__4435));
    Span4Mux_s2_h I__400 (
            .O(N__4435),
            .I(N__4432));
    Sp12to4 I__399 (
            .O(N__4432),
            .I(N__4429));
    Span12Mux_v I__398 (
            .O(N__4429),
            .I(N__4426));
    Span12Mux_v I__397 (
            .O(N__4426),
            .I(N__4423));
    Odrv12 I__396 (
            .O(N__4423),
            .I(PIO_S0_c));
    ClkMux I__395 (
            .O(N__4420),
            .I(N__4384));
    ClkMux I__394 (
            .O(N__4419),
            .I(N__4384));
    ClkMux I__393 (
            .O(N__4418),
            .I(N__4384));
    ClkMux I__392 (
            .O(N__4417),
            .I(N__4384));
    ClkMux I__391 (
            .O(N__4416),
            .I(N__4384));
    ClkMux I__390 (
            .O(N__4415),
            .I(N__4384));
    ClkMux I__389 (
            .O(N__4414),
            .I(N__4384));
    ClkMux I__388 (
            .O(N__4413),
            .I(N__4384));
    ClkMux I__387 (
            .O(N__4412),
            .I(N__4384));
    ClkMux I__386 (
            .O(N__4411),
            .I(N__4384));
    ClkMux I__385 (
            .O(N__4410),
            .I(N__4384));
    ClkMux I__384 (
            .O(N__4409),
            .I(N__4384));
    GlobalMux I__383 (
            .O(N__4384),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .I(N__4409));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .I(N__4415));
    INV \INVU409_TRANSFER_ACK.TACK_OUTnC  (
            .O(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .I(N__4413));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__4411));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .I(N__4410));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .I(N__4418));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .I(N__4417));
    INV \INVU409_TRANSFER_ACK.CIA_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .I(N__4416));
    INV \INVU409_TRANSFER_ACK.TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .I(N__4414));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net ),
            .I(N__4412));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .I(N__4420));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net ),
            .I(N__4419));
    INV \INVU409_AUTOCONFIG.ATA_BASE_7C  (
            .O(\INVU409_AUTOCONFIG.ATA_BASE_7C_net ),
            .I(N__10351));
    INV \INVU409_AUTOCONFIG.ATA_BASE_2C  (
            .O(\INVU409_AUTOCONFIG.ATA_BASE_2C_net ),
            .I(N__10357));
    INV \INVU409_AUTOCONFIG.LIDE_OUT_0C  (
            .O(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .I(N__10348));
    INV \INVU409_AUTOCONFIG.BRIDGE_BASE_1C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net ),
            .I(N__10359));
    INV \INVU409_AUTOCONFIG.BRIDGE_OUT_0C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .I(N__10349));
    INV \INVU409_AUTOCONFIG.BRIDGE_OUT_3C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .I(N__10352));
    INV \INVU409_AUTOCONFIG.STATE_0C  (
            .O(\INVU409_AUTOCONFIG.STATE_0C_net ),
            .I(N__10358));
    INV \INVU409_AUTOCONFIG.LIDE_CONFC  (
            .O(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .I(N__10363));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__10636),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_4_1_0_a2_LC_2_11_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_4_1_0_a2_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_4_1_0_a2_LC_2_11_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_AUTOCONFIG.un1_A_4_1_0_a2_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__5564),
            .in2(_gnd_net_),
            .in3(N__6270),
            .lcout(\U409_AUTOCONFIG.N_214_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.ATA_BASE10_2_LC_2_11_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE10_2_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.ATA_BASE10_2_LC_2_11_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE10_2_LC_2_11_7  (
            .in0(N__4532),
            .in1(N__4571),
            .in2(N__5802),
            .in3(N__5450),
            .lcout(\U409_AUTOCONFIG.ATA_BASE10Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_2_0__m2_0_123_i_i_a3_LC_2_12_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_2_0__m2_0_123_i_i_a3_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_2_0__m2_0_123_i_i_a3_LC_2_12_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_cnst_2_0__m2_0_123_i_i_a3_LC_2_12_3  (
            .in0(N__5541),
            .in1(N__6244),
            .in2(N__5451),
            .in3(N__5693),
            .lcout(\U409_AUTOCONFIG.N_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_2_12_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_2_12_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_2_12_4  (
            .in0(N__6243),
            .in1(N__5694),
            .in2(_gnd_net_),
            .in3(N__5540),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_7_0_62_i_i_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_o2_LC_2_12_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_o2_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_o2_LC_2_12_6 .LUT_INIT=16'b0011111000111111;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_o2_LC_2_12_6  (
            .in0(N__4479),
            .in1(N__5814),
            .in2(N__5712),
            .in3(N__5433),
            .lcout(\U409_AUTOCONFIG.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_2_12_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_2_12_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_2_12_7  (
            .in0(N__4588),
            .in1(N__5432),
            .in2(_gnd_net_),
            .in3(N__4533),
            .lcout(\U409_AUTOCONFIG.N_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_2_0_LC_3_11_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_2_0_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_2_0_LC_3_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_2_0_LC_3_11_0  (
            .in0(N__4544),
            .in1(N__5788),
            .in2(N__4583),
            .in3(N__5466),
            .lcout(\U409_AUTOCONFIG.N_67 ),
            .ltout(\U409_AUTOCONFIG.N_67_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_3_11_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_3_11_1 .LUT_INIT=16'b0011001110110011;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_3_11_1  (
            .in0(N__6294),
            .in1(N__10809),
            .in2(N__4483),
            .in3(N__5578),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_0_LC_3_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_0_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_0_LC_3_11_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_0_LC_3_11_3  (
            .in0(_gnd_net_),
            .in1(N__4543),
            .in2(_gnd_net_),
            .in3(N__4572),
            .lcout(\U409_AUTOCONFIG.N_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_2_LC_3_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_2_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_2_LC_3_11_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_2_LC_3_11_5  (
            .in0(N__5597),
            .in1(N__4545),
            .in2(N__4480),
            .in3(N__4576),
            .lcout(\U409_AUTOCONFIG.N_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_18_0_LC_3_11_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_18_0_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_18_0_LC_3_11_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_AUTOCONFIG.un1_A_18_0_LC_3_11_6  (
            .in0(N__5579),
            .in1(N__6295),
            .in2(N__4584),
            .in3(N__5467),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.un1_A_18Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_18_LC_3_11_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_18_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_18_LC_3_11_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_AUTOCONFIG.un1_A_18_LC_3_11_7  (
            .in0(N__5727),
            .in1(N__4546),
            .in2(N__4507),
            .in3(N__5789),
            .lcout(\U409_AUTOCONFIG.un1_AZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_4_0_LC_3_12_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_4_0_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_4_0_LC_3_12_1 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_4_0_LC_3_12_1  (
            .in0(N__5816),
            .in1(N__6246),
            .in2(N__5464),
            .in3(N__5696),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_3_12_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_3_12_2 .LUT_INIT=16'b0101010111010101;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_3_12_2  (
            .in0(N__10832),
            .in1(N__4659),
            .in2(N__4504),
            .in3(N__5542),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_3_12_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_3_12_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_3_12_3  (
            .in0(N__5543),
            .in1(N__6245),
            .in2(_gnd_net_),
            .in3(N__5695),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_3_12_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_3_12_4 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_3_12_4  (
            .in0(N__5115),
            .in1(N__4501),
            .in2(N__4495),
            .in3(N__5815),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_18_3_0_a2_LC_3_12_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_18_3_0_a2_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_18_3_0_a2_LC_3_12_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_AUTOCONFIG.un1_A_18_3_0_a2_LC_3_12_5  (
            .in0(N__5817),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5697),
            .lcout(\U409_AUTOCONFIG.N_196_1 ),
            .ltout(\U409_AUTOCONFIG.N_196_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_3_12_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_3_12_6 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_3_12_6  (
            .in0(N__6247),
            .in1(N__5455),
            .in2(N__4492),
            .in3(N__4489),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTc_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_3_15_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_3_15_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_3_15_0  (
            .in0(N__6074),
            .in1(N__10833),
            .in2(_gnd_net_),
            .in3(N__6026),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_3_15_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_3_15_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_3_15_4  (
            .in0(N__6507),
            .in1(N__5279),
            .in2(N__5242),
            .in3(N__5341),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_3_15_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_3_15_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_LC_3_15_5  (
            .in0(N__6607),
            .in1(N__4627),
            .in2(N__4621),
            .in3(N__5978),
            .lcout(U409_ADDRESS_DECODE_Z2_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_5_7_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_5_7_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_5_7_3  (
            .in0(N__8017),
            .in1(N__7489),
            .in2(_gnd_net_),
            .in3(N__7822),
            .lcout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_5_8_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_5_8_1 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_LC_5_8_1  (
            .in0(N__4998),
            .in1(N__4974),
            .in2(N__6406),
            .in3(N__6160),
            .lcout(\U409_AUTOCONFIG.LIDE_CONFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__9736));
    defparam \U409_AUTOCONFIG.AC_TACK_LC_5_8_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_TACK_LC_5_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_TACK_LC_5_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_AUTOCONFIG.AC_TACK_LC_5_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4975),
            .lcout(AC_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__9736));
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_5_8_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_5_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_5_8_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_CONF_LC_5_8_7  (
            .in0(_gnd_net_),
            .in1(N__5922),
            .in2(_gnd_net_),
            .in3(N__6782),
            .lcout(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__9736));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0EA21_LC_5_9_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0EA21_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0EA21_LC_5_9_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNI0EA21_LC_5_9_0  (
            .in0(N__5577),
            .in1(N__6154),
            .in2(N__5734),
            .in3(N__4618),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.ATA_BASE10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIH7AQ2_0_LC_5_9_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIH7AQ2_0_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIH7AQ2_0_LC_5_9_1 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIH7AQ2_0_LC_5_9_1  (
            .in0(N__4997),
            .in1(N__6372),
            .in2(N__4606),
            .in3(N__4966),
            .lcout(\U409_AUTOCONFIG.un1_STATE_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNISS061_3_LC_5_9_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNISS061_3_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNISS061_3_LC_5_9_2 .LUT_INIT=16'b1110111111100000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNISS061_3_LC_5_9_2  (
            .in0(N__5923),
            .in1(N__4732),
            .in2(N__6170),
            .in3(N__5089),
            .lcout(U409_AUTOCONFIG_D_OUT_0_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g0_i_a4_0_2_LC_5_10_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g0_i_a4_0_2_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g0_i_a4_0_2_LC_5_10_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.g0_i_a4_0_2_LC_5_10_3  (
            .in0(N__7862),
            .in1(N__8215),
            .in2(_gnd_net_),
            .in3(N__8004),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.g0_i_a4_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g0_i_0_0_LC_5_10_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g0_i_0_0_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g0_i_0_0_LC_5_10_4 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \U409_ADDRESS_DECODE.g0_i_0_0_LC_5_10_4  (
            .in0(N__8522),
            .in1(N__7450),
            .in2(N__4738),
            .in3(N__5188),
            .lcout(\U409_ADDRESS_DECODE.g0_i_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_0_LC_5_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_0_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.STATE_0_LC_5_10_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_0_LC_5_10_6  (
            .in0(N__10822),
            .in1(N__4973),
            .in2(N__4717),
            .in3(N__5182),
            .lcout(\U409_AUTOCONFIG.STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_5_11_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_5_11_1 .LUT_INIT=16'b1000000000100000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_5_11_1  (
            .in0(N__4644),
            .in1(N__5580),
            .in2(N__6297),
            .in3(N__5728),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.N_55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_5_11_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_5_11_2 .LUT_INIT=16'b0000101010001000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_5_11_2  (
            .in0(N__10825),
            .in1(N__4728),
            .in2(N__4735),
            .in3(N__4798),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_RNIJJLA1_LC_5_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_RNIJJLA1_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.AC_START_RNIJJLA1_LC_5_11_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_AUTOCONFIG.AC_START_RNIJJLA1_LC_5_11_3  (
            .in0(N__6396),
            .in1(N__4965),
            .in2(N__4713),
            .in3(N__5181),
            .lcout(\U409_AUTOCONFIG.N_59_1 ),
            .ltout(\U409_AUTOCONFIG.N_59_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_RNI777K2_LC_5_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_RNI777K2_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.AC_START_RNI777K2_LC_5_11_4 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \U409_AUTOCONFIG.AC_START_RNI777K2_LC_5_11_4  (
            .in0(N__10823),
            .in1(N__4678),
            .in2(N__4666),
            .in3(N__4663),
            .lcout(\U409_AUTOCONFIG.AC_START_RNI777KZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_5_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_5_11_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_5_11_5  (
            .in0(N__4770),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4633),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_5_11_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_5_11_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_5_11_6 .LUT_INIT=16'b0000101010001000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_5_11_6  (
            .in0(N__10824),
            .in1(N__5898),
            .in2(N__4648),
            .in3(N__4797),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_2_LC_5_11_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_2_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_2_LC_5_11_7 .LUT_INIT=16'b0000100010000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_2_LC_5_11_7  (
            .in0(N__4645),
            .in1(N__5581),
            .in2(N__6298),
            .in3(N__5729),
            .lcout(\U409_AUTOCONFIG.N_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_5_12_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_5_12_0 .LUT_INIT=16'b1100110000000101;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_5_12_0  (
            .in0(N__4819),
            .in1(N__5031),
            .in2(N__4810),
            .in3(N__4783),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_5_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_5_12_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_5_12_1  (
            .in0(N__7876),
            .in1(N__7661),
            .in2(N__7780),
            .in3(N__7556),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_RNI9THQ1_LC_5_12_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_RNI9THQ1_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.AC_START_RNI9THQ1_LC_5_12_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U409_AUTOCONFIG.AC_START_RNI9THQ1_LC_5_12_4  (
            .in0(N__10836),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4796),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUT_8_sqmuxa ),
            .ltout(\U409_AUTOCONFIG.BRIDGE_OUT_8_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_5_12_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_5_12_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_5_12_5 .LUT_INIT=16'b1111000100000001;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_5_12_5  (
            .in0(N__4777),
            .in1(N__4756),
            .in2(N__4744),
            .in3(N__5061),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_5_12_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_5_12_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_5_12_7  (
            .in0(N__5560),
            .in1(N__5701),
            .in2(N__6296),
            .in3(N__5448),
            .lcout(\U409_AUTOCONFIG.N_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_0_LC_5_13_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_0_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_0_LC_5_13_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_4_0_LC_5_13_1  (
            .in0(N__7973),
            .in1(N__7414),
            .in2(N__8237),
            .in3(N__8488),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_13_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_13_5 .LUT_INIT=16'b1100110000010001;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_13_5  (
            .in0(N__5733),
            .in1(N__5818),
            .in2(_gnd_net_),
            .in3(N__5465),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.LIDE_OUT_7_94_i_i_1_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_13_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_13_6 .LUT_INIT=16'b1000100000110000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_13_6  (
            .in0(N__5610),
            .in1(N__5559),
            .in2(N__4741),
            .in3(N__6233),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTc_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_5_15_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_5_15_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_5_15_0  (
            .in0(N__6619),
            .in1(N__6528),
            .in2(N__5293),
            .in3(N__5338),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_15_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_15_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__5239),
            .in2(N__4939),
            .in3(N__6081),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_5_15_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_5_15_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_5_15_6  (
            .in0(N__4936),
            .in1(N__6032),
            .in2(_gnd_net_),
            .in3(N__5991),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_LC_5_15_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_LC_5_15_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_LC_5_15_7  (
            .in0(N__4927),
            .in1(_gnd_net_),
            .in2(N__4921),
            .in3(N__4879),
            .lcout(AUTOVECTOR),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_5_16_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_5_16_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_5_16_5  (
            .in0(N__6564),
            .in1(N__4918),
            .in2(N__4900),
            .in3(N__10840),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_6_7_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_6_7_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_6_7_1  (
            .in0(N__8418),
            .in1(N__8536),
            .in2(N__8236),
            .in3(N__7540),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_6_7_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_6_7_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_6_7_2  (
            .in0(N__4873),
            .in1(N__7770),
            .in2(N__4867),
            .in3(N__7621),
            .lcout(AUTOCONFIG_SPACE),
            .ltout(AUTOCONFIG_SPACE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_6_7_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_6_7_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.D_1_i_LC_6_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4864),
            .in3(N__6401),
            .lcout(D_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_6_7_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_6_7_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_6_7_4  (
            .in0(N__6402),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9919),
            .lcout(un1_AUTOCONFIG_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_6_8_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_6_8_0 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_6_8_0 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_6_8_0  (
            .in0(N__7267),
            .in1(N__6778),
            .in2(N__6892),
            .in3(N__5844),
            .lcout(BRIDGE_BASE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net ),
            .ce(),
            .sr(N__9735));
    defparam \U409_AUTOCONFIG.ATA_BASE_5_LC_6_8_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_5_LC_6_8_2 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_5_LC_6_8_2 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_5_LC_6_8_2  (
            .in0(N__7265),
            .in1(N__6803),
            .in2(N__6891),
            .in3(N__6659),
            .lcout(ATA_BASE_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net ),
            .ce(),
            .sr(N__9735));
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_6_8_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_6_8_3 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_6_8_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_AUTOCONFIG.CONFIGENn_LC_6_8_3  (
            .in0(_gnd_net_),
            .in1(N__6777),
            .in2(_gnd_net_),
            .in3(N__6710),
            .lcout(CONFIGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net ),
            .ce(),
            .sr(N__9735));
    defparam \U409_AUTOCONFIG.ATA_BASE_4_LC_6_8_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_4_LC_6_8_4 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_4_LC_6_8_4 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_4_LC_6_8_4  (
            .in0(N__7264),
            .in1(N__6802),
            .in2(N__6930),
            .in3(N__8096),
            .lcout(ATA_BASE_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net ),
            .ce(),
            .sr(N__9735));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_6_8_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_6_8_5 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_6_8_5 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_6_8_5  (
            .in0(N__6108),
            .in1(N__7266),
            .in2(N__6786),
            .in3(N__6926),
            .lcout(BRIDGE_BASE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net ),
            .ce(),
            .sr(N__9735));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_6_8_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_6_8_6 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_6_8_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_6_8_6  (
            .in0(N__6776),
            .in1(N__6850),
            .in2(N__7277),
            .in3(N__5829),
            .lcout(BRIDGE_BASE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net ),
            .ce(),
            .sr(N__9735));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_6_9_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_6_9_1 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_6_9_1  (
            .in0(N__5035),
            .in1(N__5924),
            .in2(N__5158),
            .in3(N__6159),
            .lcout(U409_AUTOCONFIG_D_OUT_0_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g0_i_a4_1_3_LC_6_9_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g0_i_a4_1_3_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g0_i_a4_1_3_LC_6_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.g0_i_a4_1_3_LC_6_9_2  (
            .in0(N__7451),
            .in1(N__8542),
            .in2(N__7877),
            .in3(N__8222),
            .lcout(\U409_ADDRESS_DECODE.g0_i_a4_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_12_LC_6_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_12_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_12_LC_6_9_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_12_LC_6_9_3  (
            .in0(N__8388),
            .in1(N__7869),
            .in2(N__7486),
            .in3(N__8033),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.G_14_0_a7_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_10_LC_6_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_10_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_10_LC_6_9_4 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_10_LC_6_9_4  (
            .in0(_gnd_net_),
            .in1(N__8543),
            .in2(N__5002),
            .in3(N__8223),
            .lcout(\U409_TRANSFER_ACK.N_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNI25A42_0_LC_6_9_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNI25A42_0_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNI25A42_0_LC_6_9_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNI25A42_0_LC_6_9_5  (
            .in0(N__4999),
            .in1(N__4967),
            .in2(N__6387),
            .in3(N__6158),
            .lcout(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g0_i_a4_1_LC_6_10_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g0_i_a4_1_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g0_i_a4_1_LC_6_10_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U409_ADDRESS_DECODE.g0_i_a4_1_LC_6_10_2  (
            .in0(N__5194),
            .in1(N__8389),
            .in2(_gnd_net_),
            .in3(N__8010),
            .lcout(\U409_ADDRESS_DECODE.g0_i_a4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_1_LC_6_10_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_1_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_1_LC_6_10_5 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_1_LC_6_10_5  (
            .in0(N__7040),
            .in1(N__9291),
            .in2(_gnd_net_),
            .in3(N__7109),
            .lcout(U409_ADDRESS_DECODE_ROMEN_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_LC_6_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_START_LC_6_10_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_AUTOCONFIG.AC_START_LC_6_10_7  (
            .in0(N__9929),
            .in1(N__9475),
            .in2(N__10808),
            .in3(N__6717),
            .lcout(\U409_AUTOCONFIG.AC_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10350),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_11_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_11_1 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_11_1  (
            .in0(N__5170),
            .in1(N__5151),
            .in2(N__5362),
            .in3(N__5101),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .ce(),
            .sr(N__9728));
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_11_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_11_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_11_2 .LUT_INIT=16'b0101011100000010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_11_2  (
            .in0(N__5102),
            .in1(N__5140),
            .in2(N__5134),
            .in3(N__5070),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .ce(),
            .sr(N__9728));
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_11_3 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_11_3  (
            .in0(N__5122),
            .in1(N__5883),
            .in2(N__5746),
            .in3(N__5103),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .ce(),
            .sr(N__9728));
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_11_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_11_4 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_11_4  (
            .in0(N__5104),
            .in1(N__5641),
            .in2(N__5088),
            .in3(N__5745),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_0C_net ),
            .ce(),
            .sr(N__9728));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_6_11_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_6_11_6 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_6_11_6  (
            .in0(N__6177),
            .in1(N__5071),
            .in2(N__5935),
            .in3(N__5062),
            .lcout(U409_AUTOCONFIG_D_OUT_0_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIQQ061_2_LC_6_11_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIQQ061_2_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIQQ061_2_LC_6_11_7 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIQQ061_2_LC_6_11_7  (
            .in0(N__5934),
            .in1(N__5899),
            .in2(N__5887),
            .in3(N__6178),
            .lcout(U409_AUTOCONFIG_D_OUT_0_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_0_LC_6_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_0_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_0_LC_6_12_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_0_LC_6_12_1  (
            .in0(N__5278),
            .in1(N__5334),
            .in2(N__5851),
            .in3(N__5833),
            .lcout(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_0_3_144_i_i_a2_LC_6_12_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_0_3_144_i_i_a2_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_0_3_144_i_i_a2_LC_6_12_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_0_3_144_i_i_a2_LC_6_12_3  (
            .in0(N__5555),
            .in1(N__5810),
            .in2(N__6299),
            .in3(N__5702),
            .lcout(\U409_AUTOCONFIG.N_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_12_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_12_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_12_7  (
            .in0(N__6288),
            .in1(N__5449),
            .in2(N__5576),
            .in3(N__5703),
            .lcout(\U409_AUTOCONFIG.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_6_13_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_6_13_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_6_13_7  (
            .in0(N__5635),
            .in1(N__5611),
            .in2(N__5575),
            .in3(N__5431),
            .lcout(\U409_AUTOCONFIG.N_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g2_LC_6_15_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g2_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g2_LC_6_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.g2_LC_6_15_0  (
            .in0(N__6088),
            .in1(N__6621),
            .in2(N__5992),
            .in3(N__6036),
            .lcout(\U409_ADDRESS_DECODE.g2_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g2_0_LC_6_15_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g2_0_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g2_0_LC_6_15_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_ADDRESS_DECODE.g2_0_LC_6_15_2  (
            .in0(N__5339),
            .in1(N__5291),
            .in2(N__10834),
            .in3(N__5240),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.g2_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g2_9_LC_6_15_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g2_9_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g2_9_LC_6_15_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.g2_9_LC_6_15_3  (
            .in0(N__5350),
            .in1(N__5944),
            .in2(N__5344),
            .in3(N__6716),
            .lcout(\U409_ADDRESS_DECODE.g2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g2_6_LC_6_15_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g2_6_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g2_6_LC_6_15_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_ADDRESS_DECODE.g2_6_LC_6_15_6  (
            .in0(N__5340),
            .in1(N__5292),
            .in2(N__10835),
            .in3(N__5241),
            .lcout(U409_ADDRESS_DECODE_g2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g2_5_LC_6_15_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g2_5_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g2_5_LC_6_15_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.g2_5_LC_6_15_7  (
            .in0(N__6620),
            .in1(N__6087),
            .in2(N__6037),
            .in3(N__5987),
            .lcout(\U409_ADDRESS_DECODE.g2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g2_4_LC_6_16_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g2_4_LC_6_16_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g2_4_LC_6_16_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_ADDRESS_DECODE.g2_4_LC_6_16_5  (
            .in0(N__7013),
            .in1(N__7086),
            .in2(_gnd_net_),
            .in3(N__6529),
            .lcout(\U409_ADDRESS_DECODE.g2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_6_1_LC_7_7_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_6_1_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_6_1_LC_7_7_1 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.un1_Z2_SPACE_6_1_LC_7_7_1  (
            .in0(N__8537),
            .in1(N__6658),
            .in2(N__8252),
            .in3(N__8092),
            .lcout(\U409_ADDRESS_DECODE.un1_Z2_SPACE_6Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_9_LC_7_7_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_9_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_9_LC_7_7_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_9_LC_7_7_2  (
            .in0(N__7824),
            .in1(N__7491),
            .in2(N__8253),
            .in3(N__8538),
            .lcout(\U409_TRANSFER_ACK.G_14_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g2_10_LC_7_7_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g2_10_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g2_10_LC_7_7_6 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.g2_10_LC_7_7_6  (
            .in0(N__7823),
            .in1(N__7185),
            .in2(N__7779),
            .in3(N__6946),
            .lcout(\U409_ADDRESS_DECODE.g2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g0_i_o4_1_LC_7_8_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g0_i_o4_1_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g0_i_o4_1_LC_7_8_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \U409_ADDRESS_DECODE.g0_i_o4_1_LC_7_8_1  (
            .in0(N__7343),
            .in1(N__7658),
            .in2(N__7596),
            .in3(N__7552),
            .lcout(\U409_ADDRESS_DECODE.g0_i_o4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_6_0_LC_7_8_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_6_0_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_6_0_LC_7_8_2 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.un1_Z2_SPACE_6_0_LC_7_8_2  (
            .in0(N__7659),
            .in1(N__7588),
            .in2(N__7558),
            .in3(N__7342),
            .lcout(\U409_ADDRESS_DECODE.un1_Z2_SPACE_6Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_1_LC_7_8_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_1_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_1_LC_7_8_3 .LUT_INIT=16'b0000000010000100;
    LogicCell40 \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_1_LC_7_8_3  (
            .in0(N__8119),
            .in1(N__8419),
            .in2(N__8028),
            .in3(N__6698),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.un1_Z2_SPACE_7Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_3_LC_7_8_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_3_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_3_LC_7_8_4 .LUT_INIT=16'b1100000000110000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_3_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(N__7481),
            .in2(N__5938),
            .in3(N__7318),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.un1_Z2_SPACE_7Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_LC_7_8_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_LC_7_8_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_Z2_SPACE_LC_7_8_5  (
            .in0(N__6421),
            .in1(N__6415),
            .in2(N__6409),
            .in3(N__7570),
            .lcout(\U409_ADDRESS_DECODE.un1_Z2_SPACEZ0 ),
            .ltout(\U409_ADDRESS_DECODE.un1_Z2_SPACEZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_ROM_EN_LC_7_8_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_ROM_EN_LC_7_8_6 .SEQ_MODE=4'b1001;
    defparam \U409_ADDRESS_DECODE.ATA_ROM_EN_LC_7_8_6 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_ROM_EN_LC_7_8_6  (
            .in0(N__6400),
            .in1(N__9492),
            .in2(N__6328),
            .in3(N__10014),
            .lcout(U409_ADDRESS_DECODE_ATA_ROM_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10356),
            .ce(),
            .sr(N__9733));
    defparam \U409_ADDRESS_DECODE.g2_11_LC_7_9_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g2_11_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g2_11_LC_7_9_0 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.g2_11_LC_7_9_0  (
            .in0(N__7490),
            .in1(N__7323),
            .in2(N__8040),
            .in3(N__8126),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.g2Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_ROM_EN_RNITNPB5_LC_7_9_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_ROM_EN_RNITNPB5_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_ROM_EN_RNITNPB5_LC_7_9_1 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_ROM_EN_RNITNPB5_LC_7_9_1  (
            .in0(N__10015),
            .in1(N__6325),
            .in2(N__6316),
            .in3(N__6313),
            .lcout(U409_ADDRESS_DECODE_ATA_ROM_d),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNI0FVT2_0_LC_7_9_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNI0FVT2_0_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNI0FVT2_0_LC_7_9_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNI0FVT2_0_LC_7_9_4  (
            .in0(N__6120),
            .in1(N__6301),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_AUTOCONFIG.STATE_RNI0FVT2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIHQ9A3_LC_7_9_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIHQ9A3_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIHQ9A3_LC_7_9_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIHQ9A3_LC_7_9_5  (
            .in0(N__6300),
            .in1(N__6176),
            .in2(_gnd_net_),
            .in3(N__6121),
            .lcout(\U409_AUTOCONFIG.LIDE_CONF_RNIHQ9AZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_0_LC_7_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_0_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_0_LC_7_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_0_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(N__8626),
            .in2(_gnd_net_),
            .in3(N__8753),
            .lcout(\U409_TRANSFER_ACK.CO1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_2_LC_7_10_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_2_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_2_LC_7_10_0 .LUT_INIT=16'b0100010000010001;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_2_LC_7_10_0  (
            .in0(N__6715),
            .in1(N__6527),
            .in2(_gnd_net_),
            .in3(N__6109),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_4_LC_7_10_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_4_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_4_LC_7_10_1 .LUT_INIT=16'b0110000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_4_LC_7_10_1  (
            .in0(N__7041),
            .in1(N__7110),
            .in2(N__6091),
            .in3(N__10776),
            .lcout(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_8_LC_7_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_8_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_8_LC_7_10_5 .LUT_INIT=16'b1111111111011110;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_8_LC_7_10_5  (
            .in0(N__8532),
            .in1(N__6451),
            .in2(N__6670),
            .in3(N__6714),
            .lcout(\U409_TRANSFER_ACK.G_14_0_o7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g0_i_o4_0_LC_7_10_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g0_i_o4_0_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g0_i_o4_0_LC_7_10_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \U409_ADDRESS_DECODE.g0_i_o4_0_LC_7_10_6  (
            .in0(N__6669),
            .in1(N__8098),
            .in2(N__8241),
            .in3(N__8531),
            .lcout(\U409_ADDRESS_DECODE.g0_i_o4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_7_11_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_7_11_3 .LUT_INIT=16'b0111111110111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_7_11_3  (
            .in0(N__6748),
            .in1(N__6640),
            .in2(N__6634),
            .in3(N__6625),
            .lcout(U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_0_LC_7_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_0_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_0_LC_7_13_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_0_LC_7_13_3  (
            .in0(N__6565),
            .in1(N__8505),
            .in2(_gnd_net_),
            .in3(N__8221),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_13_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_13_4  (
            .in0(N__6541),
            .in1(N__7487),
            .in2(N__6544),
            .in3(N__9276),
            .lcout(CIA_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_7_13_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_7_13_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_7_13_7  (
            .in0(N__7030),
            .in1(N__7099),
            .in2(_gnd_net_),
            .in3(N__8018),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.g2_7_LC_7_15_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.g2_7_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.g2_7_LC_7_15_3 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \U409_ADDRESS_DECODE.g2_7_LC_7_15_3  (
            .in0(N__7029),
            .in1(N__6535),
            .in2(N__7085),
            .in3(N__6517),
            .lcout(),
            .ltout(U409_ADDRESS_DECODE_g2_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_11_LC_7_15_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_11_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_11_LC_7_15_4 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_11_LC_7_15_4  (
            .in0(N__6460),
            .in1(_gnd_net_),
            .in2(N__6454),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.G_14_0_o7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_8_6_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_8_6_0 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_8_6_0  (
            .in0(N__9304),
            .in1(N__6967),
            .in2(N__7665),
            .in3(N__6955),
            .lcout(U409_ADDRESS_DECODE_un1_RTC_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_8_6_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_8_6_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_8_6_4  (
            .in0(N__8251),
            .in1(N__8548),
            .in2(N__7870),
            .in3(N__7734),
            .lcout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3 ),
            .ltout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_8_6_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_8_6_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_8_6_5  (
            .in0(N__6966),
            .in1(N__9303),
            .in2(N__6949),
            .in3(N__7654),
            .lcout(U409_ADDRESS_DECODE_un1_RTC_ENn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_2_LC_8_7_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_2_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_2_LC_8_7_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_2_LC_8_7_1  (
            .in0(N__7735),
            .in1(N__7838),
            .in2(N__7186),
            .in3(N__6944),
            .lcout(U409_ADDRESS_DECODE_un1_Z2_SPACE_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.ATA_BASE_2_LC_8_7_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_2_LC_8_7_2 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_2_LC_8_7_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_2_LC_8_7_2  (
            .in0(N__6945),
            .in1(N__7278),
            .in2(N__6846),
            .in3(N__7240),
            .lcout(ATA_BASE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_2C_net ),
            .ce(),
            .sr(N__9734));
    defparam \U409_AUTOCONFIG.ATA_BASE_7_LC_8_8_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_7_LC_8_8_0 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_7_LC_8_8_0 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_7_LC_8_8_0  (
            .in0(N__7217),
            .in1(N__6805),
            .in2(N__8127),
            .in3(N__7296),
            .lcout(ATA_BASE_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_7C_net ),
            .ce(),
            .sr(N__9730));
    defparam \U409_AUTOCONFIG.ATA_BASE_0_LC_8_8_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_0_LC_8_8_1 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_0_LC_8_8_1 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_0_LC_8_8_1  (
            .in0(N__7292),
            .in1(N__7234),
            .in2(N__6931),
            .in3(N__7344),
            .lcout(ATA_BASE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_7C_net ),
            .ce(),
            .sr(N__9730));
    defparam \U409_AUTOCONFIG.ATA_BASE_1_LC_8_8_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_1_LC_8_8_3 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_1_LC_8_8_3 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_1_LC_8_8_3  (
            .in0(N__7293),
            .in1(N__7235),
            .in2(N__7597),
            .in3(N__6873),
            .lcout(ATA_BASE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_7C_net ),
            .ce(),
            .sr(N__9730));
    defparam \U409_AUTOCONFIG.ATA_BASE_6_LC_8_8_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_6_LC_8_8_4 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_6_LC_8_8_4 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_6_LC_8_8_4  (
            .in0(N__6836),
            .in1(N__6804),
            .in2(N__7324),
            .in3(N__7295),
            .lcout(ATA_BASE_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_7C_net ),
            .ce(),
            .sr(N__9730));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_8_8_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_8_8_6 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_8_8_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_8_8_6  (
            .in0(N__7218),
            .in1(N__7297),
            .in2(N__6747),
            .in3(N__6787),
            .lcout(BRIDGE_BASE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_7C_net ),
            .ce(),
            .sr(N__9730));
    defparam \U409_AUTOCONFIG.ATA_BASE_3_LC_8_8_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_3_LC_8_8_7 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.ATA_BASE_3_LC_8_8_7 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_3_LC_8_8_7  (
            .in0(N__7294),
            .in1(N__7236),
            .in2(N__7219),
            .in3(N__7184),
            .lcout(ATA_BASE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_7C_net ),
            .ce(),
            .sr(N__9730));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_8_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_8_9_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__8627),
            .in2(_gnd_net_),
            .in3(N__8754),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__9729));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_8_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_8_9_2 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_8_9_2  (
            .in0(N__7132),
            .in1(N__8062),
            .in2(N__7165),
            .in3(N__8056),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__9729));
    defparam \U409_ADDRESS_DECODE.ATA_ROM_EN_RNITAAO4_LC_8_10_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_ROM_EN_RNITAAO4_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_ROM_EN_RNITAAO4_LC_8_10_2 .LUT_INIT=16'b0000010100010101;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_ROM_EN_RNITAAO4_LC_8_10_2  (
            .in0(N__7156),
            .in1(N__7147),
            .in2(N__10034),
            .in3(N__7138),
            .lcout(U409_ADDRESS_DECODE_ATA_ROM_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_8_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_8_10_6 .LUT_INIT=16'b0011110000010100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_8_10_6  (
            .in0(N__8590),
            .in1(N__7125),
            .in2(N__8668),
            .in3(N__8572),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__9726));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_8_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_8_10_7 .LUT_INIT=16'b0100110010000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_8_10_7  (
            .in0(N__8663),
            .in1(N__8554),
            .in2(N__7126),
            .in3(N__8795),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__9726));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_8_11_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_8_11_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_8_11_2  (
            .in0(N__7111),
            .in1(N__7488),
            .in2(N__7042),
            .in3(N__7969),
            .lcout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_8_12_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_8_12_0 .LUT_INIT=16'b1110101011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_8_12_0  (
            .in0(N__8217),
            .in1(N__7879),
            .in2(N__7778),
            .in3(N__7687),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.un2_REGSPACEn_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_LC_8_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_LC_8_12_1 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \U409_ADDRESS_DECODE.un2_REGSPACEn_LC_8_12_1  (
            .in0(N__8545),
            .in1(N__7693),
            .in2(N__7882),
            .in3(N__7699),
            .lcout(U409_ADDRESS_DECODE_un2_REGSPACEn_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.REG_SPACE_2_LC_8_12_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.REG_SPACE_2_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.REG_SPACE_2_LC_8_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.REG_SPACE_2_LC_8_12_4  (
            .in0(N__8216),
            .in1(N__7878),
            .in2(N__7777),
            .in3(N__7666),
            .lcout(\U409_ADDRESS_DECODE.REG_SPACEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_8_12_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_8_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_8_12_5  (
            .in0(N__8029),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7461),
            .lcout(\U409_ADDRESS_DECODE.REG_SPACE_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_8_12_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_8_12_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_8_12_6  (
            .in0(N__7462),
            .in1(N__8030),
            .in2(_gnd_net_),
            .in3(N__8544),
            .lcout(\U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.LOWROM_3_LC_9_6_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.LOWROM_3_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.LOWROM_3_LC_9_6_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_ADDRESS_DECODE.LOWROM_3_LC_9_6_4  (
            .in0(N__8041),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7492),
            .lcout(\U409_ADDRESS_DECODE.LOWROMZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_0_LC_9_7_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_0_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_0_LC_9_7_4 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_0_LC_9_7_4  (
            .in0(N__8925),
            .in1(N__8940),
            .in2(_gnd_net_),
            .in3(N__9498),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_7_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_7_5 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_7_5  (
            .in0(N__8547),
            .in1(N__8434),
            .in2(N__8387),
            .in3(N__8304),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_4_LC_9_8_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_4_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_4_LC_9_8_1 .LUT_INIT=16'b0110011011111111;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_4_LC_9_8_1  (
            .in0(N__7660),
            .in1(N__7595),
            .in2(_gnd_net_),
            .in3(N__7569),
            .lcout(\U409_TRANSFER_ACK.g0_0_0_o6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_6_LC_9_8_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_6_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_6_LC_9_8_5 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_6_LC_9_8_5  (
            .in0(N__7557),
            .in1(N__7482),
            .in2(N__7348),
            .in3(N__7322),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.G_14_0_o7_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_3_LC_9_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_3_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_3_LC_9_8_6 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_3_LC_9_8_6  (
            .in0(N__8068),
            .in1(_gnd_net_),
            .in2(N__8269),
            .in3(N__8266),
            .lcout(\U409_TRANSFER_ACK.G_14_0_o7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_7_LC_9_8_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_7_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_7_LC_9_8_7 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_7_LC_9_8_7  (
            .in0(N__8032),
            .in1(N__8254),
            .in2(N__8128),
            .in3(N__8097),
            .lcout(\U409_TRANSFER_ACK.G_14_0_o7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_9_0 .LUT_INIT=16'b0011000100010001;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_9_0  (
            .in0(N__8055),
            .in1(N__8589),
            .in2(N__8680),
            .in3(N__8571),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_LC_9_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_LC_9_9_1 .LUT_INIT=16'b1010101010101011;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_LC_9_9_1  (
            .in0(N__8750),
            .in1(N__8623),
            .in2(N__8667),
            .in3(N__8787),
            .lcout(\U409_TRANSFER_ACK.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_1_0_LC_9_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_1_0_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_1_0_LC_9_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_1_0_LC_9_9_2  (
            .in0(N__8786),
            .in1(N__8657),
            .in2(N__8629),
            .in3(N__8749),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20 ),
            .ltout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_9_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_9_9_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_9_9_3  (
            .in0(N__8588),
            .in1(_gnd_net_),
            .in2(N__8044),
            .in3(N__8676),
            .lcout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_9_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_9_4  (
            .in0(N__8625),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8662),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER20_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_5_LC_9_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_5_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_5_LC_9_9_5 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_5_LC_9_9_5  (
            .in0(N__8031),
            .in1(N__7909),
            .in2(N__7900),
            .in3(N__8788),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.G_14_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_9_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_9_9_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_9_9_6  (
            .in0(N__8624),
            .in1(N__8661),
            .in2(N__7885),
            .in3(N__8751),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.G_14_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_9_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_9_9_7 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_9_9_7  (
            .in0(N__8698),
            .in1(N__10035),
            .in2(N__8689),
            .in3(N__8686),
            .lcout(\U409_TRANSFER_ACK.ROMENn_1_sqmuxa_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_s_LC_9_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_s_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_s_LC_9_10_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_s_LC_9_10_3  (
            .in0(N__8420),
            .in1(N__9488),
            .in2(_gnd_net_),
            .in3(N__10388),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER15_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_0_LC_9_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_0_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_0_LC_9_10_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_0_LC_9_10_6  (
            .in0(N__8656),
            .in1(N__8752),
            .in2(N__8628),
            .in3(N__8789),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_3_LC_9_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_3_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_3_LC_9_10_7 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_3_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8575),
            .in3(N__8570),
            .lcout(\U409_TRANSFER_ACK.ROMENn_1_sqmuxa_0_c ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_9_11_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_9_11_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_9_11_7  (
            .in0(N__8546),
            .in1(N__8433),
            .in2(N__8377),
            .in3(N__8311),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_9_13_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_9_13_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__9295),
            .in2(_gnd_net_),
            .in3(N__9315),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn),
            .ltout(U409_ADDRESS_DECODE_un1_REGSPACEn_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_9_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_9_13_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_9_13_3  (
            .in0(N__9947),
            .in1(N__8956),
            .in2(N__8293),
            .in3(N__9896),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_6_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_6_1 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_6_1  (
            .in0(N__8902),
            .in1(N__8965),
            .in2(N__8881),
            .in3(N__10391),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net ),
            .ce(),
            .sr(N__9731));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_6_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_6_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_6_3  (
            .in0(N__8971),
            .in1(N__10390),
            .in2(_gnd_net_),
            .in3(N__8964),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net ),
            .ce(),
            .sr(N__9731));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_10_7_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_10_7_2 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_10_7_2  (
            .in0(N__10741),
            .in1(N__8952),
            .in2(N__8929),
            .in3(N__9499),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_7_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_7_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_7_3  (
            .in0(N__10752),
            .in1(N__9652),
            .in2(_gnd_net_),
            .in3(N__9674),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNI7KT7_LC_10_7_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNI7KT7_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNI7KT7_LC_10_7_5 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNI7KT7_LC_10_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8860),
            .in3(N__8709),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIBQIN_LC_10_7_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIBQIN_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIBQIN_LC_10_7_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIBQIN_LC_10_7_6  (
            .in0(N__8896),
            .in1(N__8877),
            .in2(N__8866),
            .in3(N__9510),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER6 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_7_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_7_7 .LUT_INIT=16'b0000000010001010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_7_7  (
            .in0(N__10751),
            .in1(N__9653),
            .in2(N__8863),
            .in3(N__9675),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_8_0 .LUT_INIT=16'b0101111100001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_8_0  (
            .in0(N__10207),
            .in1(N__9688),
            .in2(N__10237),
            .in3(N__8859),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__9727));
    defparam \U409_TRANSFER_ACK.ROMENn_LC_10_8_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_10_8_1 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_10_8_1 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_LC_10_8_1  (
            .in0(N__8817),
            .in1(N__8845),
            .in2(N__8806),
            .in3(N__8839),
            .lcout(ROMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__9727));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_8_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_8_2 .LUT_INIT=16'b0111111100100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_8_2  (
            .in0(N__8802),
            .in1(N__8761),
            .in2(N__8719),
            .in3(N__8710),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__9727));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_10_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_10_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_10_8_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_10_8_3  (
            .in0(N__10431),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__9727));
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_10_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_10_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_10_8_4 .LUT_INIT=16'b0111000001110001;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_LC_10_8_4  (
            .in0(N__9655),
            .in1(N__9676),
            .in2(N__9848),
            .in3(N__9628),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__9727));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_10_8_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_10_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_10_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9550),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__9727));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CKM1_7_LC_10_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CKM1_7_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CKM1_7_LC_10_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CKM1_7_LC_10_9_0  (
            .in0(N__9022),
            .in1(N__9046),
            .in2(N__9127),
            .in3(N__8987),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_4_LC_10_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_4_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_4_LC_10_9_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_4_LC_10_9_1  (
            .in0(N__9412),
            .in1(N__10105),
            .in2(N__8992),
            .in3(N__9106),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_9_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_9_2 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_9_2  (
            .in0(N__10106),
            .in1(N__9025),
            .in2(N__10156),
            .in3(N__10134),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__10080));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_3 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_3 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_3  (
            .in0(N__9126),
            .in1(N__9004),
            .in2(N__10138),
            .in3(N__8989),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__10080));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_3_LC_10_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_3_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_3_LC_10_9_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_3_LC_10_9_4  (
            .in0(N__9023),
            .in1(N__9413),
            .in2(N__9052),
            .in3(N__10104),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_7_LC_10_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_7_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_7_LC_10_9_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_7_LC_10_9_5  (
            .in0(N__9125),
            .in1(N__8988),
            .in2(N__8974),
            .in3(N__9105),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_7_LC_10_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_7_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_7_LC_10_9_6 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_7_LC_10_9_6  (
            .in0(N__9493),
            .in1(N__10387),
            .in2(N__9133),
            .in3(N__9527),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__9124),
            .in2(N__9130),
            .in3(N__9003),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__10080));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_10_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_10_0 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_10_0  (
            .in0(N__9416),
            .in1(N__9094),
            .in2(_gnd_net_),
            .in3(N__10132),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__10076));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_1 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_1  (
            .in0(N__9093),
            .in1(_gnd_net_),
            .in2(N__9076),
            .in3(N__9418),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__10076));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_10_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_10_2  (
            .in0(_gnd_net_),
            .in1(N__9090),
            .in2(_gnd_net_),
            .in3(N__9064),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_10_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_10_10_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_10_10_3  (
            .in0(N__9092),
            .in1(_gnd_net_),
            .in2(N__9075),
            .in3(N__9415),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_10_4 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_10_4  (
            .in0(N__9051),
            .in1(_gnd_net_),
            .in2(N__9097),
            .in3(N__10131),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__10076));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_10_5  (
            .in0(N__9091),
            .in1(N__9414),
            .in2(N__9074),
            .in3(N__9050),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_10_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__10111),
            .in2(N__9028),
            .in3(N__9024),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_7 .LUT_INIT=16'b0001000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_7  (
            .in0(N__9497),
            .in1(N__9417),
            .in2(N__10393),
            .in3(N__9529),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__10076));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_13_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_13_5 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_13_5  (
            .in0(N__9391),
            .in1(N__9354),
            .in2(N__9385),
            .in3(N__10767),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_DATA_BUFFERS.un1_BUFENn_LC_10_14_3 .C_ON=1'b0;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_LC_10_14_3 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \U409_DATA_BUFFERS.un1_BUFENn_LC_10_14_3  (
            .in0(N__9325),
            .in1(N__9297),
            .in2(N__9361),
            .in3(N__9948),
            .lcout(BUFENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_10_14_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_10_14_5 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_10_14_5  (
            .in0(N__9324),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9296),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNI692L_0_LC_11_3_3 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNI692L_0_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNI692L_0_LC_11_3_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_CIA.VMA_RNI692L_0_LC_11_3_3  (
            .in0(N__10695),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9970),
            .lcout(CIA_ENABLE),
            .ltout(CIA_ENABLE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_11_3_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_11_3_4 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_11_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9220),
            .in3(N__9217),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS0n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_3_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_3_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_3_6  (
            .in0(N__9178),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9172),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS1n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_5_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10270),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .ce(),
            .sr(N__9732));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_5_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_5_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_5_6  (
            .in0(N__10724),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9969),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .ce(),
            .sr(N__9732));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_6_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_6_0 .LUT_INIT=16'b0000011111110111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_6_0  (
            .in0(N__10283),
            .in1(N__10268),
            .in2(N__10202),
            .in3(N__9687),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_6_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_6_1 .LUT_INIT=16'b0000001010001010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_6_1  (
            .in0(N__10739),
            .in1(N__10230),
            .in2(N__9697),
            .in3(N__9694),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_6_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_6_6 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_6_6  (
            .in0(N__10284),
            .in1(N__10267),
            .in2(N__10203),
            .in3(N__10248),
            .lcout(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_11_7_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_11_7_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_11_7_2  (
            .in0(N__9549),
            .in1(N__10389),
            .in2(_gnd_net_),
            .in3(N__9562),
            .lcout(\U409_TRANSFER_ACK.N_17_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_7_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_7_3 .LUT_INIT=16'b0010001100100111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_7_3  (
            .in0(N__9673),
            .in1(N__9575),
            .in2(N__9654),
            .in3(N__9627),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_7_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_7_4 .LUT_INIT=16'b0010111000101110;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_11_7_4  (
            .in0(N__9576),
            .in1(N__10740),
            .in2(N__9616),
            .in3(_gnd_net_),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_11_7_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_11_7_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__9561),
            .in2(_gnd_net_),
            .in3(N__9548),
            .lcout(\U409_TRANSFER_ACK.N_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_8_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_8_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_8_1 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_8_1  (
            .in0(N__9511),
            .in1(N__9535),
            .in2(_gnd_net_),
            .in3(N__9528),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .ce(),
            .sr(N__10081));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_8_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_8_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_8_6  (
            .in0(N__10155),
            .in1(N__10110),
            .in2(_gnd_net_),
            .in3(N__10133),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .ce(),
            .sr(N__10081));
    defparam \U409_ADDRESS_DECODE.ATA_ROM_EN_RNIBHHS6_LC_11_9_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_ROM_EN_RNIBHHS6_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_ROM_EN_RNIBHHS6_LC_11_9_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_ROM_EN_RNIBHHS6_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__10048),
            .in2(_gnd_net_),
            .in3(N__10036),
            .lcout(U409_ADDRESS_DECODE_un1_ATA_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__10884),
            .in2(_gnd_net_),
            .in3(N__10537),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10480),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_11_10_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_11_10_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__10556),
            .in2(_gnd_net_),
            .in3(N__10577),
            .lcout(\U409_CIA.CLK_CIA6_4 ),
            .ltout(\U409_CIA.CLK_CIA6_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_11_10_1 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_11_10_1 .LUT_INIT=16'b0010000010000000;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_11_10_1  (
            .in0(N__10591),
            .in1(N__10462),
            .in2(N__9976),
            .in3(N__10535),
            .lcout(),
            .ltout(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_11_10_2 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_11_10_2 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \U409_CIA.VMA_LC_11_10_2  (
            .in0(N__10536),
            .in1(N__9901),
            .in2(N__9973),
            .in3(N__9962),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10478),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_11_10_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_11_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10883),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10478),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_11_13_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_11_13_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_11_13_2  (
            .in0(N__9949),
            .in1(N__9897),
            .in2(_gnd_net_),
            .in3(N__9855),
            .lcout(TCIn_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_7.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_7.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10392),
            .lcout(GB_BUFFER_CLK40_IN_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_6_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_6_0 .LUT_INIT=16'b0001000000011111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_6_0  (
            .in0(N__10285),
            .in1(N__10269),
            .in2(N__10201),
            .in3(N__10249),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.N_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_6_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_6_1 .LUT_INIT=16'b0010101000001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_6_1  (
            .in0(N__10714),
            .in1(N__10229),
            .in2(N__10210),
            .in3(N__10191),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__10532),
            .in2(N__10885),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__10924),
            .in2(_gnd_net_),
            .in3(N__10168),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__10479),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_12_9_2 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_12_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__10942),
            .in2(_gnd_net_),
            .in3(N__10165),
            .lcout(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__10459),
            .in2(_gnd_net_),
            .in3(N__10162),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__10479),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__10903),
            .in2(_gnd_net_),
            .in3(N__10159),
            .lcout(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_12_9_5 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_12_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_6_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(N__10579),
            .in2(_gnd_net_),
            .in3(N__10597),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ),
            .clk(N__10479),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_12_9_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_12_9_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_7_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__10560),
            .in2(_gnd_net_),
            .in3(N__10594),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10479),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_1_LC_12_9_7 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_1_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_1_LC_12_9_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_CIA.VMA_RNO_1_LC_12_9_7  (
            .in0(N__10943),
            .in1(N__10925),
            .in2(N__10908),
            .in3(N__10880),
            .lcout(\U409_CIA.un1_CIA_CLK_COUNT_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_12_10_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_12_10_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_12_10_0  (
            .in0(N__10852),
            .in1(N__10507),
            .in2(N__10501),
            .in3(N__10585),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10477),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_12_10_1 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_12_10_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_0_LC_12_10_1  (
            .in0(N__10578),
            .in1(N__10882),
            .in2(N__10561),
            .in3(N__10534),
            .lcout(),
            .ltout(\U409_CIA.CLK_CIA6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_LC_12_10_2 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLK_CIA_LC_12_10_2 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \U409_CIA.CLK_CIA_LC_12_10_2  (
            .in0(N__10399),
            .in1(N__10417),
            .in2(N__10540),
            .in3(N__10907),
            .lcout(CLK_CIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10477),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_12_10_3 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_12_10_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__10460),
            .in2(_gnd_net_),
            .in3(N__10533),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_2 ),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_10_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_12_10_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_12_10_4  (
            .in0(N__10497),
            .in1(N__10851),
            .in2(N__10489),
            .in3(N__10486),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10477),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_12_10_5 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_12_10_5 .LUT_INIT=16'b0000000000011000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_1_LC_12_10_5  (
            .in0(N__10945),
            .in1(N__10461),
            .in2(N__10424),
            .in3(N__10927),
            .lcout(\U409_CIA.CLK_CIA_r_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_12_10_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_12_10_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_12_10_7  (
            .in0(N__10944),
            .in1(N__10926),
            .in2(N__10909),
            .in3(N__10881),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_6.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_6.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_18_6 (
            .in0(N__10745),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_13_5_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_13_5_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_13_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_13_5_0  (
            .in0(_gnd_net_),
            .in1(N__11193),
            .in2(_gnd_net_),
            .in3(N__11214),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11846),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_13_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_13_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_13_5_1 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_13_5_1  (
            .in0(N__11043),
            .in1(N__10997),
            .in2(N__11461),
            .in3(N__11069),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11846),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_13_5_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_13_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_13_5_3 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_13_5_3  (
            .in0(N__11042),
            .in1(N__11125),
            .in2(N__11002),
            .in3(N__11068),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11846),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNINQJI1_4_LC_13_5_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNINQJI1_4_LC_13_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNINQJI1_4_LC_13_5_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNINQJI1_4_LC_13_5_4  (
            .in0(N__11098),
            .in1(N__11137),
            .in2(N__11116),
            .in3(N__11473),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(\U409_TICK.TICK603_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_13_5_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_13_5_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_13_5_5 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_13_5_5  (
            .in0(N__11497),
            .in1(N__11045),
            .in2(N__10624),
            .in3(N__10998),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11846),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_13_5_6 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_13_5_6 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK60_LC_13_5_6  (
            .in0(N__10996),
            .in1(N__10608),
            .in2(N__11077),
            .in3(N__11044),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11846),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_13_6_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_13_6_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_13_6_0  (
            .in0(N__11075),
            .in1(N__10995),
            .in2(N__11047),
            .in3(N__11662),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11847),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIA84S_11_LC_13_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIA84S_11_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIA84S_11_LC_13_6_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIA84S_11_LC_13_6_1  (
            .in0(N__11410),
            .in1(N__11152),
            .in2(N__11170),
            .in3(N__11395),
            .lcout(\U409_TICK.TICK603_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_13_6_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_13_6_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_13_6_2  (
            .in0(N__11074),
            .in1(N__10994),
            .in2(N__11046),
            .in3(N__11350),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11847),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIRP4S_14_LC_13_6_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIRP4S_14_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIRP4S_14_LC_13_6_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_TICK.COUNTER60_RNIRP4S_14_LC_13_6_3  (
            .in0(N__11674),
            .in1(N__11449),
            .in2(N__11365),
            .in3(N__11488),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_13_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_13_6_4 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_13_6_4  (
            .in0(N__11073),
            .in1(N__10993),
            .in2(N__11080),
            .in3(N__11192),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11847),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_13_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_13_6_5 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_13_6_5  (
            .in0(N__10992),
            .in1(N__11076),
            .in2(N__11437),
            .in3(N__11041),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11847),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDAFF_10_LC_13_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDAFF_10_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDAFF_10_LC_13_6_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDAFF_10_LC_13_6_6  (
            .in0(N__11380),
            .in1(N__11425),
            .in2(_gnd_net_),
            .in3(N__11191),
            .lcout(),
            .ltout(\U409_TICK.TICK603_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIVPLP1_16_LC_13_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIVPLP1_16_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIVPLP1_16_LC_13_6_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNIVPLP1_16_LC_13_6_7  (
            .in0(N__11215),
            .in1(N__11649),
            .in2(N__11011),
            .in3(N__11008),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_13_7_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_13_7_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_13_7_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_13_7_0  (
            .in0(N__11290),
            .in1(N__11323),
            .in2(N__11536),
            .in3(N__11248),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11849),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_13_7_1 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_13_7_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK50_LC_13_7_1  (
            .in0(N__11247),
            .in1(N__10956),
            .in2(N__11329),
            .in3(N__11292),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11849),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_13_7_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_13_7_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_13_7_2  (
            .in0(N__11291),
            .in1(N__11324),
            .in2(N__11509),
            .in3(N__11249),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11849),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNI3J3V_10_LC_13_7_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNI3J3V_10_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNI3J3V_10_LC_13_7_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNI3J3V_10_LC_13_7_4  (
            .in0(N__11770),
            .in1(N__11596),
            .in2(N__11638),
            .in3(N__11731),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_13_7_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_13_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_13_7_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_13_7_5  (
            .in0(N__11322),
            .in1(N__11289),
            .in2(N__11258),
            .in3(N__11740),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11849),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_13_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_13_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_13_7_7  (
            .in0(_gnd_net_),
            .in1(N__11637),
            .in2(_gnd_net_),
            .in3(N__11619),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11849),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_13_8_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_13_8_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_13_8_0  (
            .in0(N__11286),
            .in1(N__11320),
            .in2(N__11260),
            .in3(N__11704),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11851),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIJAR11_3_LC_13_8_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIJAR11_3_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIJAR11_3_LC_13_8_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIJAR11_3_LC_13_8_1  (
            .in0(N__11524),
            .in1(N__11581),
            .in2(N__11551),
            .in3(N__11791),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_13_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_13_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_13_8_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_13_8_2  (
            .in0(N__11287),
            .in1(N__11257),
            .in2(N__11086),
            .in3(N__11878),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11851),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIDMCS_11_LC_13_8_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIDMCS_11_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIDMCS_11_LC_13_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIDMCS_11_LC_13_8_3  (
            .in0(N__11695),
            .in1(N__11716),
            .in2(N__11755),
            .in3(N__11890),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_13_8_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_13_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_13_8_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_13_8_4  (
            .in0(N__11288),
            .in1(N__11321),
            .in2(N__11083),
            .in3(N__11779),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11851),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIG9CP_4_LC_13_8_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIG9CP_4_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIG9CP_4_LC_13_8_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TICK.COUNTER50_RNIG9CP_4_LC_13_8_5  (
            .in0(N__11821),
            .in1(N__11566),
            .in2(_gnd_net_),
            .in3(N__11617),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNI02282_16_LC_13_8_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNI02282_16_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNI02282_16_LC_13_8_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TICK.COUNTER50_RNI02282_16_LC_13_8_6  (
            .in0(N__11865),
            .in1(N__11341),
            .in2(N__11335),
            .in3(N__11806),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_13_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_13_8_7 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_13_8_7  (
            .in0(N__11319),
            .in1(N__11253),
            .in2(N__11332),
            .in3(N__11618),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11851),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_13_9_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_13_9_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_13_9_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_13_9_2  (
            .in0(N__11328),
            .in1(N__11293),
            .in2(N__11259),
            .in3(N__11683),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11853),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_5_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_5_0  (
            .in0(_gnd_net_),
            .in1(N__11210),
            .in2(N__11194),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_14_5_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_14_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_14_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_14_5_1  (
            .in0(_gnd_net_),
            .in1(N__11166),
            .in2(_gnd_net_),
            .in3(N__11155),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__11848),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_14_5_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_14_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_14_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(N__11151),
            .in2(_gnd_net_),
            .in3(N__11140),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__11848),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_14_5_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_14_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_14_5_3  (
            .in0(_gnd_net_),
            .in1(N__11136),
            .in2(_gnd_net_),
            .in3(N__11119),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_14_5_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_14_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_14_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_14_5_4  (
            .in0(_gnd_net_),
            .in1(N__11112),
            .in2(_gnd_net_),
            .in3(N__11101),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__11848),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_14_5_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_14_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(N__11097),
            .in2(_gnd_net_),
            .in3(N__11491),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_14_5_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_14_5_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_14_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_14_5_6  (
            .in0(_gnd_net_),
            .in1(N__11487),
            .in2(_gnd_net_),
            .in3(N__11476),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__11848),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_14_5_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_14_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_14_5_7  (
            .in0(_gnd_net_),
            .in1(N__11472),
            .in2(_gnd_net_),
            .in3(N__11452),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_14_6_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_14_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_14_6_0  (
            .in0(_gnd_net_),
            .in1(N__11448),
            .in2(_gnd_net_),
            .in3(N__11428),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_14_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_14_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(N__11424),
            .in2(_gnd_net_),
            .in3(N__11413),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__11850),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_14_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_14_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_14_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(N__11409),
            .in2(_gnd_net_),
            .in3(N__11398),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__11850),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_14_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_14_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_14_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(N__11394),
            .in2(_gnd_net_),
            .in3(N__11383),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__11850),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_14_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_14_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_14_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(N__11379),
            .in2(_gnd_net_),
            .in3(N__11368),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__11850),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_14_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_14_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_14_6_5  (
            .in0(_gnd_net_),
            .in1(N__11361),
            .in2(_gnd_net_),
            .in3(N__11344),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_14_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_14_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_14_6_6  (
            .in0(_gnd_net_),
            .in1(N__11673),
            .in2(_gnd_net_),
            .in3(N__11656),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_14_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_14_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_14_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(N__11650),
            .in2(_gnd_net_),
            .in3(N__11653),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11850),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_7_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(N__11633),
            .in2(N__11620),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_14_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_14_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(N__11595),
            .in2(_gnd_net_),
            .in3(N__11584),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__11852),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_14_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_14_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__11580),
            .in2(_gnd_net_),
            .in3(N__11569),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__11852),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_14_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_14_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(N__11565),
            .in2(_gnd_net_),
            .in3(N__11554),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__11852),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(N__11547),
            .in2(_gnd_net_),
            .in3(N__11527),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(N__11520),
            .in2(_gnd_net_),
            .in3(N__11500),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_14_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_14_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(N__11820),
            .in2(_gnd_net_),
            .in3(N__11809),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__11852),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_14_7_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_14_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(N__11805),
            .in2(_gnd_net_),
            .in3(N__11794),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__11852),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_8_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__11790),
            .in2(_gnd_net_),
            .in3(N__11773),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_14_8_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_14_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_14_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_14_8_1  (
            .in0(_gnd_net_),
            .in1(N__11769),
            .in2(_gnd_net_),
            .in3(N__11758),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__11854),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_8_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_14_8_2  (
            .in0(_gnd_net_),
            .in1(N__11751),
            .in2(_gnd_net_),
            .in3(N__11734),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_14_8_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_14_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(N__11730),
            .in2(_gnd_net_),
            .in3(N__11719),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__11854),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_8_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(N__11715),
            .in2(_gnd_net_),
            .in3(N__11698),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_8_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(N__11694),
            .in2(_gnd_net_),
            .in3(N__11677),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_8_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(N__11889),
            .in2(_gnd_net_),
            .in3(N__11872),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_14_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_14_8_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(N__11866),
            .in2(_gnd_net_),
            .in3(N__11869),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11854),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

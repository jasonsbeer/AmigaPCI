-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 22 2025 01:34:21

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U400_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U400_TOP
entity U400_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    MA : out std_logic_vector(12 downto 0);
    A : in std_logic_vector(31 downto 0);
    LBENn : out std_logic;
    CS0n : out std_logic;
    UUBEn : out std_logic;
    TAn : out std_logic;
    CLK40 : in std_logic;
    RnW : in std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    WEn : out std_logic;
    LLBEn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    RASn : out std_logic;
    CS1n : out std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic);
end U400_TOP;

-- Architecture of U400_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U400_TOP is

signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2569\ : std_logic;
signal \CLK40_ibuf_gb_io_gb_input\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_29\ : std_logic;
signal \A_c_28\ : std_logic;
signal \A_c_27\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_\ : std_logic;
signal \U400_SDRAM.un1_TA_COUNTER26_0_cascade_\ : std_logic;
signal \U400_SDRAM.TA_COUNTER23_cascade_\ : std_logic;
signal \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0\ : std_logic;
signal \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_\ : std_logic;
signal \U400_SDRAM.CO1\ : std_logic;
signal \U400_SDRAM.CO1_cascade_\ : std_logic;
signal \A_c_21\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \A_c_22\ : std_logic;
signal \BANK1_c\ : std_logic;
signal \INVU400_SDRAM.BANK0C_net\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_a3_0_cascade_\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_1\ : std_logic;
signal \U400_SDRAM.N_208_cascade_\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \CASn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \INVU400_SDRAM.RASnC_net\ : std_logic;
signal \A_c_24\ : std_logic;
signal \A_c_18\ : std_logic;
signal \MA_c_8\ : std_logic;
signal \A_c_17\ : std_logic;
signal \A_c_9\ : std_logic;
signal \MA_c_7\ : std_logic;
signal \INVU400_SDRAM.MA_8C_net\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_16\ : std_logic;
signal \MA_c_6\ : std_logic;
signal \INVU400_SDRAM.MA_6C_net\ : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_1\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_2\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_3\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_4\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_5\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_6\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_7\ : std_logic;
signal \INVU400_SDRAM.REFRESH_COUNTER_2C_net\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_2\ : std_logic;
signal \U400_SDRAM.un1_TA_COUNTER26_2_0\ : std_logic;
signal \TA_OUT\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_1\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_3\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_0_sqmuxa\ : std_logic;
signal \U400_SDRAM.TA_COUNTER27\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_\ : std_logic;
signal \INVU400_SDRAM.BURSTC_net\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER52_2_0_i_1_cascade_\ : std_logic;
signal \U400_SDRAM.N_23\ : std_logic;
signal \U400_SDRAM.N_255\ : std_logic;
signal \U400_SDRAM.TACK_7_iv_i_i_0_cascade_\ : std_logic;
signal \U400_SDRAM.TACK_7_iv_i_i_1\ : std_logic;
signal \U400_SDRAM.N_15\ : std_logic;
signal \U400_SDRAM.RAM_CYCLE_e_1\ : std_logic;
signal \U400_SDRAM.N_6\ : std_logic;
signal \RnW_c\ : std_logic;
signal \INVU400_SDRAM.RAM_CYCLEC_net\ : std_logic;
signal \CS0n_c\ : std_logic;
signal \A_c_19\ : std_logic;
signal \MA_c_9\ : std_logic;
signal \INVU400_SDRAM.CS0_ENC_net\ : std_logic;
signal \INVU400_SDRAM.REFRESH_COUNTER_0C_net\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_0\ : std_logic;
signal \U400_SDRAM.BURSTZ0\ : std_logic;
signal \U400_SDRAM.TA_EN11_m\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U400_SDRAM.N_205_cascade_\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CMD_1C_net\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en\ : std_logic;
signal \U400_SDRAM.un1_REFRESH_COUNTERlto7_4\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_8\ : std_logic;
signal \U400_SDRAM.un1_REFRESH_COUNTERlto7_5\ : std_logic;
signal \U400_SDRAM.N_189\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_1_32_i_0_i_1_1_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_1_32_i_0_i_1_cascade_\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CMD_0C_net\ : std_logic;
signal \U400_SDRAM.N_128\ : std_logic;
signal \U400_SDRAM.N_185\ : std_logic;
signal \U400_SDRAM.RAM_CYCLEZ0\ : std_logic;
signal \U400_SDRAM.N_75_cascade_\ : std_logic;
signal \U400_SDRAM.CS1_EN_0\ : std_logic;
signal \U400_SDRAM.CS1_EN_7_i_0_o3_0_cascade_\ : std_logic;
signal \U400_SDRAM.N_159\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U400_SDRAM.CS0_ENZ0\ : std_logic;
signal \U400_SDRAM.N_159_cascade_\ : std_logic;
signal \U400_SDRAM.N_75\ : std_logic;
signal \U400_SDRAM.CS0_EN_0\ : std_logic;
signal \U400_SDRAM.N_250\ : std_logic;
signal \U400_SDRAM.N_176_cascade_\ : std_logic;
signal \U400_SDRAM.CS1_ENZ0\ : std_logic;
signal \CS1n_c\ : std_logic;
signal \A_c_26\ : std_logic;
signal \MA_c_12\ : std_logic;
signal \INVU400_SDRAM.CS1nC_net\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \UUBEn_c\ : std_logic;
signal \U400_SDRAM.TA_COUNTER23\ : std_logic;
signal \U400_SDRAM.TACKZ0\ : std_logic;
signal \CLK40_c_g\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0\ : std_logic;
signal \U400_SDRAM.N_252_cascade_\ : std_logic;
signal \U400_SDRAM.N_200_cascade_\ : std_logic;
signal \U400_SDRAM.N_199\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_61_i_i_1_cascade_\ : std_logic;
signal \U400_SDRAM.N_17\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CMD_2C_net\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_i_a2_0_1_1\ : std_logic;
signal \U400_SDRAM.N_228\ : std_logic;
signal \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5Z0Z_0_cascade_\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_3C_net\ : std_logic;
signal \U400_SDRAM.N_203\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_i_0\ : std_logic;
signal \U400_SDRAM.N_126_cascade_\ : std_logic;
signal \U400_SDRAM.N_129_cascade_\ : std_logic;
signal \U400_SDRAM.N_257_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_1_0\ : std_logic;
signal \U400_SDRAM.N_133\ : std_logic;
signal \U400_SDRAM.N_133_cascade_\ : std_logic;
signal \U400_SDRAM.N_139\ : std_logic;
signal \U400_SDRAM.N_141_cascade_\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTER_RNIVV903Z0Z_8\ : std_logic;
signal \U400_SDRAM.RAM_CYCLE_STARTZ0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_2_0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U400_SDRAM.N_181_cascade_\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_0C_net\ : std_logic;
signal \A_c_25\ : std_logic;
signal \MA_c_11\ : std_logic;
signal \U400_SDRAM.N_257\ : std_logic;
signal \INVU400_SDRAM.MA_11C_net\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_14\ : std_logic;
signal \MA_c_4\ : std_logic;
signal \MA_c_5\ : std_logic;
signal \INVU400_SDRAM.MA_4C_net\ : std_logic;
signal \U400_SDRAM.N_150\ : std_logic;
signal \U400_SDRAM.N_150_cascade_\ : std_logic;
signal \U400_SDRAM.N_252\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_61_i_i_a3_1_0_cascade_\ : std_logic;
signal \U400_SDRAM.N_201\ : std_logic;
signal \TA_EN_i_ess\ : std_logic;
signal \N_529_i\ : std_logic;
signal \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5Z0Z_0\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_1C_net\ : std_logic;
signal \U400_SDRAM.N_129\ : std_logic;
signal \U400_SDRAM.N_260\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_1\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_3\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U400_SDRAM.N_37\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_2C_net\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U400_SDRAM.WRITE_CYCLEZ0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U400_SDRAM.N_161_cascade_\ : std_logic;
signal \U400_SDRAM.N_183\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U400_SDRAM.N_126\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U400_SDRAM.N_138\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a3_1_0_0\ : std_logic;
signal \U400_SDRAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7JZ0\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U400_SDRAM.MAc_0_0\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_10\ : std_logic;
signal \MA_c_0\ : std_logic;
signal \A_c_20\ : std_logic;
signal \MA_c_10\ : std_logic;
signal \INVU400_SDRAM.MA_0C_net\ : std_logic;
signal \UMBEn_c\ : std_logic;
signal \LLBEn_c\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \LMBEn_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U400_SDRAM.N_220\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U400_SDRAM.BURST8\ : std_logic;
signal \A_c_31\ : std_logic;
signal \U400_ADDRESS_DECODE_RAM_SPACE_0_a3_3\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \N_220_3_i\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_13\ : std_logic;
signal \MA_c_3\ : std_logic;
signal \INVU400_SDRAM.MA_3C_net\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U400_SDRAM.MAc_1_0\ : std_logic;
signal \MA_c_2\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ1Z_0\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U400_SDRAM.MAc_9_0\ : std_logic;
signal \MA_c_1\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \INVU400_SDRAM.MA_2C_net\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \MA_wire\ : std_logic_vector(12 downto 0);
signal \A_wire\ : std_logic_vector(31 downto 0);
signal \CASn_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \UUBEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \LLBEn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \TAn_wire\ : std_logic;
signal \LBENn_wire\ : std_logic;
signal \CS1n_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CS0n_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CLK40_wire\ : std_logic;

begin
    MA <= \MA_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    BANK1 <= \BANK1_wire\;
    UUBEn <= \UUBEn_wire\;
    \SIZ_wire\ <= SIZ;
    LLBEn <= \LLBEn_wire\;
    \TSn_wire\ <= TSn;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    \RESETn_wire\ <= RESETn;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    TAn <= \TAn_wire\;
    LBENn <= \LBENn_wire\;
    CS1n <= \CS1n_wire\;
    WEn <= \WEn_wire\;
    \RnW_wire\ <= RnW;
    CS0n <= \CS0n_wire\;
    LMBEn <= \LMBEn_wire\;
    \CLK40_wire\ <= CLK40;

    \MA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7004\,
            DIN => \N__7003\,
            DOUT => \N__7002\,
            PACKAGEPIN => \MA_wire\(7)
        );

    \MA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7004\,
            PADOUT => \N__7003\,
            PADIN => \N__7002\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2797\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6995\,
            DIN => \N__6994\,
            DOUT => \N__6993\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6995\,
            PADOUT => \N__6994\,
            PADIN => \N__6993\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6986\,
            DIN => \N__6985\,
            DOUT => \N__6984\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6986\,
            PADOUT => \N__6985\,
            PADIN => \N__6984\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2881\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6977\,
            DIN => \N__6976\,
            DOUT => \N__6975\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6977\,
            PADOUT => \N__6976\,
            PADIN => \N__6975\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2677\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6968\,
            DIN => \N__6967\,
            DOUT => \N__6966\,
            PACKAGEPIN => \MA_wire\(8)
        );

    \MA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6968\,
            PADOUT => \N__6967\,
            PADIN => \N__6966\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2830\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6959\,
            DIN => \N__6958\,
            DOUT => \N__6957\,
            PACKAGEPIN => \MA_wire\(10)
        );

    \MA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6959\,
            PADOUT => \N__6958\,
            PADIN => \N__6957\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5881\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6950\,
            DIN => \N__6949\,
            DOUT => \N__6948\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6950\,
            PADOUT => \N__6949\,
            PADIN => \N__6948\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6941\,
            DIN => \N__6940\,
            DOUT => \N__6939\,
            PACKAGEPIN => \MA_wire\(2)
        );

    \MA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6941\,
            PADOUT => \N__6940\,
            PADIN => \N__6939\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6325\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6932\,
            DIN => \N__6931\,
            DOUT => \N__6930\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6932\,
            PADOUT => \N__6931\,
            PADIN => \N__6930\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6923\,
            DIN => \N__6922\,
            DOUT => \N__6921\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6923\,
            PADOUT => \N__6922\,
            PADIN => \N__6921\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6914\,
            DIN => \N__6913\,
            DOUT => \N__6912\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6914\,
            PADOUT => \N__6913\,
            PADIN => \N__6912\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3727\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6905\,
            DIN => \N__6904\,
            DOUT => \N__6903\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6905\,
            PADOUT => \N__6904\,
            PADIN => \N__6903\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6896\,
            DIN => \N__6895\,
            DOUT => \N__6894\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6896\,
            PADOUT => \N__6895\,
            PADIN => \N__6894\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6887\,
            DIN => \N__6886\,
            DOUT => \N__6885\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6887\,
            PADOUT => \N__6886\,
            PADIN => \N__6885\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6878\,
            DIN => \N__6877\,
            DOUT => \N__6876\,
            PACKAGEPIN => \MA_wire\(12)
        );

    \MA_obuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6878\,
            PADOUT => \N__6877\,
            PADIN => \N__6876\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3763\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6869\,
            DIN => \N__6868\,
            DOUT => \N__6867\,
            PACKAGEPIN => \MA_wire\(1)
        );

    \MA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6869\,
            PADOUT => \N__6868\,
            PADIN => \N__6867\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5947\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6860\,
            DIN => \N__6859\,
            DOUT => \N__6858\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6860\,
            PADOUT => \N__6859\,
            PADIN => \N__6858\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6851\,
            DIN => \N__6850\,
            DOUT => \N__6849\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6851\,
            PADOUT => \N__6850\,
            PADIN => \N__6849\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6842\,
            DIN => \N__6841\,
            DOUT => \N__6840\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6842\,
            PADOUT => \N__6841\,
            PADIN => \N__6840\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6833\,
            DIN => \N__6832\,
            DOUT => \N__6831\,
            PACKAGEPIN => \MA_wire\(4)
        );

    \MA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6833\,
            PADOUT => \N__6832\,
            PADIN => \N__6831\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4186\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6824\,
            DIN => \N__6823\,
            DOUT => \N__6822\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6824\,
            PADOUT => \N__6823\,
            PADIN => \N__6822\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6815\,
            DIN => \N__6814\,
            DOUT => \N__6813\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6815\,
            PADOUT => \N__6814\,
            PADIN => \N__6813\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6806\,
            DIN => \N__6805\,
            DOUT => \N__6804\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6806\,
            PADOUT => \N__6805\,
            PADIN => \N__6804\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5866\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6797\,
            DIN => \N__6796\,
            DOUT => \N__6795\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6797\,
            PADOUT => \N__6796\,
            PADIN => \N__6795\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6788\,
            DIN => \N__6787\,
            DOUT => \N__6786\,
            PACKAGEPIN => \MA_wire\(9)
        );

    \MA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6788\,
            PADOUT => \N__6787\,
            PADIN => \N__6786\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3091\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6779\,
            DIN => \N__6778\,
            DOUT => \N__6777\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6779\,
            PADOUT => \N__6778\,
            PADIN => \N__6777\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5875\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6770\,
            DIN => \N__6769\,
            DOUT => \N__6768\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6770\,
            PADOUT => \N__6769\,
            PADIN => \N__6768\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6761\,
            DIN => \N__6760\,
            DOUT => \N__6759\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6761\,
            PADOUT => \N__6760\,
            PADIN => \N__6759\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6752\,
            DIN => \N__6751\,
            DOUT => \N__6750\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6752\,
            PADOUT => \N__6751\,
            PADIN => \N__6750\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3751\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6743\,
            DIN => \N__6742\,
            DOUT => \N__6741\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6743\,
            PADOUT => \N__6742\,
            PADIN => \N__6741\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6734\,
            DIN => \N__6733\,
            DOUT => \N__6732\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6734\,
            PADOUT => \N__6733\,
            PADIN => \N__6732\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6725\,
            DIN => \N__6724\,
            DOUT => \N__6723\,
            PACKAGEPIN => \MA_wire\(3)
        );

    \MA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6725\,
            PADOUT => \N__6724\,
            PADIN => \N__6723\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5371\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6716\,
            DIN => \N__6715\,
            DOUT => \N__6714\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6716\,
            PADOUT => \N__6715\,
            PADIN => \N__6714\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6707\,
            DIN => \N__6706\,
            DOUT => \N__6705\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6707\,
            PADOUT => \N__6706\,
            PADIN => \N__6705\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6698\,
            DIN => \N__6697\,
            DOUT => \N__6696\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6698\,
            PADOUT => \N__6697\,
            PADIN => \N__6696\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6689\,
            DIN => \N__6688\,
            DOUT => \N__6687\,
            PACKAGEPIN => \MA_wire\(6)
        );

    \MA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6689\,
            PADOUT => \N__6688\,
            PADIN => \N__6687\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2761\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6680\,
            DIN => \N__6679\,
            DOUT => \N__6678\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6680\,
            PADOUT => \N__6679\,
            PADIN => \N__6678\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6671\,
            DIN => \N__6670\,
            DOUT => \N__6669\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6671\,
            PADOUT => \N__6670\,
            PADIN => \N__6669\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6662\,
            DIN => \N__6661\,
            DOUT => \N__6660\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6662\,
            PADOUT => \N__6661\,
            PADIN => \N__6660\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6653\,
            DIN => \N__6652\,
            DOUT => \N__6651\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6653\,
            PADOUT => \N__6652\,
            PADIN => \N__6651\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2893\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6644\,
            DIN => \N__6643\,
            DOUT => \N__6642\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6644\,
            PADOUT => \N__6643\,
            PADIN => \N__6642\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6635\,
            DIN => \N__6634\,
            DOUT => \N__6633\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6635\,
            PADOUT => \N__6634\,
            PADIN => \N__6633\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2716\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6626\,
            DIN => \N__6625\,
            DOUT => \N__6624\,
            PACKAGEPIN => \MA_wire\(11)
        );

    \MA_obuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6626\,
            PADOUT => \N__6625\,
            PADIN => \N__6624\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4258\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6617\,
            DIN => \N__6616\,
            DOUT => \N__6615\,
            PACKAGEPIN => \TAn_wire\
        );

    \TAn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6617\,
            PADOUT => \N__6616\,
            PADIN => \N__6615\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4117\,
            DIN0 => OPEN,
            DOUT0 => \N__2926\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6608\,
            DIN => \N__6607\,
            DOUT => \N__6606\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6608\,
            PADOUT => \N__6607\,
            PADIN => \N__6606\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6599\,
            DIN => \N__6598\,
            DOUT => \N__6597\,
            PACKAGEPIN => \MA_wire\(5)
        );

    \MA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6599\,
            PADOUT => \N__6598\,
            PADIN => \N__6597\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4171\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6590\,
            DIN => \N__6589\,
            DOUT => \N__6588\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6590\,
            PADOUT => \N__6589\,
            PADIN => \N__6588\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6581\,
            DIN => \N__6580\,
            DOUT => \N__6579\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6581\,
            PADOUT => \N__6580\,
            PADIN => \N__6579\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LBENn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6572\,
            DIN => \N__6571\,
            DOUT => \N__6570\,
            PACKAGEPIN => \LBENn_wire\
        );

    \LBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6572\,
            PADOUT => \N__6571\,
            PADIN => \N__6570\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5404\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6563\,
            DIN => \N__6562\,
            DOUT => \N__6561\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6563\,
            PADOUT => \N__6562\,
            PADIN => \N__6561\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6554\,
            DIN => \N__6553\,
            DOUT => \N__6552\,
            PACKAGEPIN => \CS1n_wire\
        );

    \CS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6554\,
            PADOUT => \N__6553\,
            PADIN => \N__6552\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3793\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6545\,
            DIN => \N__6544\,
            DOUT => \N__6543\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6545\,
            PADOUT => \N__6544\,
            PADIN => \N__6543\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6536\,
            DIN => \N__6535\,
            DOUT => \N__6534\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6536\,
            PADOUT => \N__6535\,
            PADIN => \N__6534\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6527\,
            DIN => \N__6526\,
            DOUT => \N__6525\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6527\,
            PADOUT => \N__6526\,
            PADIN => \N__6525\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6518\,
            DIN => \N__6517\,
            DOUT => \N__6516\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6518\,
            PADOUT => \N__6517\,
            PADIN => \N__6516\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6509\,
            DIN => \N__6508\,
            DOUT => \N__6507\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6509\,
            PADOUT => \N__6508\,
            PADIN => \N__6507\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2872\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6500\,
            DIN => \N__6499\,
            DOUT => \N__6498\,
            PACKAGEPIN => \MA_wire\(0)
        );

    \MA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6500\,
            PADOUT => \N__6499\,
            PADIN => \N__6498\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4468\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6491\,
            DIN => \N__6490\,
            DOUT => \N__6489\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6491\,
            PADOUT => \N__6490\,
            PADIN => \N__6489\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6482\,
            DIN => \N__6481\,
            DOUT => \N__6480\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6482\,
            PADOUT => \N__6481\,
            PADIN => \N__6480\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6473\,
            DIN => \N__6472\,
            DOUT => \N__6471\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6473\,
            PADOUT => \N__6472\,
            PADIN => \N__6471\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6464\,
            DIN => \N__6463\,
            DOUT => \N__6462\,
            PACKAGEPIN => \CS0n_wire\
        );

    \CS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6464\,
            PADOUT => \N__6463\,
            PADIN => \N__6462\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3124\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6455\,
            DIN => \N__6454\,
            DOUT => \N__6453\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6455\,
            PADOUT => \N__6454\,
            PADIN => \N__6453\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6446\,
            DIN => \N__6445\,
            DOUT => \N__6444\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6446\,
            PADOUT => \N__6445\,
            PADIN => \N__6444\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5785\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6437\,
            DIN => \N__6436\,
            DOUT => \N__6435\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6437\,
            PADOUT => \N__6436\,
            PADIN => \N__6435\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6428\,
            DIN => \N__6427\,
            DOUT => \N__6426\,
            PACKAGEPIN => \CLK40_wire\
        );

    \CLK40_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6428\,
            PADOUT => \N__6427\,
            PADIN => \N__6426\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_ibuf_gb_io_gb_input\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1516\ : InMux
    port map (
            O => \N__6409\,
            I => \N__6406\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__6406\,
            I => \N__6403\
        );

    \I__1514\ : Span4Mux_s2_v
    port map (
            O => \N__6403\,
            I => \N__6400\
        );

    \I__1513\ : IoSpan4Mux
    port map (
            O => \N__6400\,
            I => \N__6397\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__6397\,
            I => \A_c_4\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__6394\,
            I => \N__6391\
        );

    \I__1510\ : InMux
    port map (
            O => \N__6391\,
            I => \N__6388\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__6388\,
            I => \A_c_12\
        );

    \I__1508\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6380\
        );

    \I__1507\ : InMux
    port map (
            O => \N__6384\,
            I => \N__6377\
        );

    \I__1506\ : InMux
    port map (
            O => \N__6383\,
            I => \N__6372\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__6380\,
            I => \N__6367\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__6377\,
            I => \N__6367\
        );

    \I__1503\ : InMux
    port map (
            O => \N__6376\,
            I => \N__6364\
        );

    \I__1502\ : InMux
    port map (
            O => \N__6375\,
            I => \N__6361\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__6372\,
            I => \N__6356\
        );

    \I__1500\ : Span4Mux_h
    port map (
            O => \N__6367\,
            I => \N__6351\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__6364\,
            I => \N__6351\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__6361\,
            I => \N__6348\
        );

    \I__1497\ : InMux
    port map (
            O => \N__6360\,
            I => \N__6343\
        );

    \I__1496\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6343\
        );

    \I__1495\ : Span4Mux_v
    port map (
            O => \N__6356\,
            I => \N__6338\
        );

    \I__1494\ : Span4Mux_v
    port map (
            O => \N__6351\,
            I => \N__6338\
        );

    \I__1493\ : Span4Mux_h
    port map (
            O => \N__6348\,
            I => \N__6335\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__6343\,
            I => \N__6332\
        );

    \I__1491\ : Odrv4
    port map (
            O => \N__6338\,
            I => \U400_SDRAM.MAc_1_0\
        );

    \I__1490\ : Odrv4
    port map (
            O => \N__6335\,
            I => \U400_SDRAM.MAc_1_0\
        );

    \I__1489\ : Odrv4
    port map (
            O => \N__6332\,
            I => \U400_SDRAM.MAc_1_0\
        );

    \I__1488\ : IoInMux
    port map (
            O => \N__6325\,
            I => \N__6322\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__6322\,
            I => \MA_c_2\
        );

    \I__1486\ : CascadeMux
    port map (
            O => \N__6319\,
            I => \N__6315\
        );

    \I__1485\ : InMux
    port map (
            O => \N__6318\,
            I => \N__6311\
        );

    \I__1484\ : InMux
    port map (
            O => \N__6315\,
            I => \N__6308\
        );

    \I__1483\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6305\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__6311\,
            I => \N__6292\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__6308\,
            I => \N__6292\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__6305\,
            I => \N__6289\
        );

    \I__1479\ : InMux
    port map (
            O => \N__6304\,
            I => \N__6286\
        );

    \I__1478\ : InMux
    port map (
            O => \N__6303\,
            I => \N__6283\
        );

    \I__1477\ : InMux
    port map (
            O => \N__6302\,
            I => \N__6278\
        );

    \I__1476\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6278\
        );

    \I__1475\ : InMux
    port map (
            O => \N__6300\,
            I => \N__6275\
        );

    \I__1474\ : InMux
    port map (
            O => \N__6299\,
            I => \N__6272\
        );

    \I__1473\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6267\
        );

    \I__1472\ : InMux
    port map (
            O => \N__6297\,
            I => \N__6267\
        );

    \I__1471\ : Span4Mux_s2_v
    port map (
            O => \N__6292\,
            I => \N__6264\
        );

    \I__1470\ : Span4Mux_s1_v
    port map (
            O => \N__6289\,
            I => \N__6257\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__6286\,
            I => \N__6257\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__6283\,
            I => \N__6257\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__6278\,
            I => \N__6250\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__6275\,
            I => \N__6250\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__6272\,
            I => \N__6247\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__6267\,
            I => \N__6244\
        );

    \I__1463\ : Sp12to4
    port map (
            O => \N__6264\,
            I => \N__6241\
        );

    \I__1462\ : Span4Mux_h
    port map (
            O => \N__6257\,
            I => \N__6238\
        );

    \I__1461\ : InMux
    port map (
            O => \N__6256\,
            I => \N__6235\
        );

    \I__1460\ : InMux
    port map (
            O => \N__6255\,
            I => \N__6232\
        );

    \I__1459\ : Span4Mux_v
    port map (
            O => \N__6250\,
            I => \N__6229\
        );

    \I__1458\ : Span4Mux_v
    port map (
            O => \N__6247\,
            I => \N__6226\
        );

    \I__1457\ : Sp12to4
    port map (
            O => \N__6244\,
            I => \N__6217\
        );

    \I__1456\ : Span12Mux_s6_h
    port map (
            O => \N__6241\,
            I => \N__6217\
        );

    \I__1455\ : Sp12to4
    port map (
            O => \N__6238\,
            I => \N__6217\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__6235\,
            I => \N__6217\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__6232\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__6229\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__6226\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1450\ : Odrv12
    port map (
            O => \N__6217\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1449\ : InMux
    port map (
            O => \N__6208\,
            I => \N__6205\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__6205\,
            I => \N__6200\
        );

    \I__1447\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6195\
        );

    \I__1446\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6192\
        );

    \I__1445\ : Span4Mux_h
    port map (
            O => \N__6200\,
            I => \N__6185\
        );

    \I__1444\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6182\
        );

    \I__1443\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6179\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__6195\,
            I => \N__6176\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__6192\,
            I => \N__6173\
        );

    \I__1440\ : InMux
    port map (
            O => \N__6191\,
            I => \N__6168\
        );

    \I__1439\ : InMux
    port map (
            O => \N__6190\,
            I => \N__6168\
        );

    \I__1438\ : InMux
    port map (
            O => \N__6189\,
            I => \N__6163\
        );

    \I__1437\ : InMux
    port map (
            O => \N__6188\,
            I => \N__6163\
        );

    \I__1436\ : Sp12to4
    port map (
            O => \N__6185\,
            I => \N__6156\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__6182\,
            I => \N__6156\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__6179\,
            I => \N__6153\
        );

    \I__1433\ : Span4Mux_s3_v
    port map (
            O => \N__6176\,
            I => \N__6150\
        );

    \I__1432\ : Span4Mux_h
    port map (
            O => \N__6173\,
            I => \N__6143\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__6168\,
            I => \N__6143\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6163\,
            I => \N__6143\
        );

    \I__1429\ : InMux
    port map (
            O => \N__6162\,
            I => \N__6140\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6137\
        );

    \I__1427\ : Span12Mux_s10_v
    port map (
            O => \N__6156\,
            I => \N__6134\
        );

    \I__1426\ : Span4Mux_h
    port map (
            O => \N__6153\,
            I => \N__6129\
        );

    \I__1425\ : Span4Mux_v
    port map (
            O => \N__6150\,
            I => \N__6129\
        );

    \I__1424\ : Sp12to4
    port map (
            O => \N__6143\,
            I => \N__6124\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__6140\,
            I => \N__6124\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__6137\,
            I => \U400_SDRAM.SDRAM_CMDZ1Z_0\
        );

    \I__1421\ : Odrv12
    port map (
            O => \N__6134\,
            I => \U400_SDRAM.SDRAM_CMDZ1Z_0\
        );

    \I__1420\ : Odrv4
    port map (
            O => \N__6129\,
            I => \U400_SDRAM.SDRAM_CMDZ1Z_0\
        );

    \I__1419\ : Odrv12
    port map (
            O => \N__6124\,
            I => \U400_SDRAM.SDRAM_CMDZ1Z_0\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__6115\,
            I => \N__6110\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__6114\,
            I => \N__6105\
        );

    \I__1416\ : InMux
    port map (
            O => \N__6113\,
            I => \N__6100\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6097\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6109\,
            I => \N__6094\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__6108\,
            I => \N__6091\
        );

    \I__1412\ : InMux
    port map (
            O => \N__6105\,
            I => \N__6082\
        );

    \I__1411\ : InMux
    port map (
            O => \N__6104\,
            I => \N__6082\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6103\,
            I => \N__6079\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__6100\,
            I => \N__6073\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__6097\,
            I => \N__6073\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__6094\,
            I => \N__6070\
        );

    \I__1406\ : InMux
    port map (
            O => \N__6091\,
            I => \N__6065\
        );

    \I__1405\ : InMux
    port map (
            O => \N__6090\,
            I => \N__6065\
        );

    \I__1404\ : InMux
    port map (
            O => \N__6089\,
            I => \N__6060\
        );

    \I__1403\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6060\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6087\,
            I => \N__6057\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__6082\,
            I => \N__6050\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__6079\,
            I => \N__6050\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6043\
        );

    \I__1398\ : Span4Mux_v
    port map (
            O => \N__6073\,
            I => \N__6037\
        );

    \I__1397\ : Span4Mux_s3_v
    port map (
            O => \N__6070\,
            I => \N__6037\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__6065\,
            I => \N__6030\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__6060\,
            I => \N__6030\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6057\,
            I => \N__6030\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6056\,
            I => \N__6026\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6055\,
            I => \N__6023\
        );

    \I__1391\ : Span4Mux_s2_v
    port map (
            O => \N__6050\,
            I => \N__6020\
        );

    \I__1390\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6017\
        );

    \I__1389\ : InMux
    port map (
            O => \N__6048\,
            I => \N__6012\
        );

    \I__1388\ : InMux
    port map (
            O => \N__6047\,
            I => \N__6012\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6046\,
            I => \N__6009\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__6043\,
            I => \N__6006\
        );

    \I__1385\ : InMux
    port map (
            O => \N__6042\,
            I => \N__6003\
        );

    \I__1384\ : Span4Mux_h
    port map (
            O => \N__6037\,
            I => \N__5998\
        );

    \I__1383\ : Span4Mux_s3_v
    port map (
            O => \N__6030\,
            I => \N__5998\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6029\,
            I => \N__5995\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__6026\,
            I => \N__5990\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__6023\,
            I => \N__5990\
        );

    \I__1379\ : Span4Mux_v
    port map (
            O => \N__6020\,
            I => \N__5987\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6017\,
            I => \N__5984\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__6012\,
            I => \N__5975\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__6009\,
            I => \N__5975\
        );

    \I__1375\ : Span4Mux_h
    port map (
            O => \N__6006\,
            I => \N__5975\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__6003\,
            I => \N__5975\
        );

    \I__1373\ : Span4Mux_v
    port map (
            O => \N__5998\,
            I => \N__5972\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__5995\,
            I => \N__5965\
        );

    \I__1371\ : Span4Mux_v
    port map (
            O => \N__5990\,
            I => \N__5965\
        );

    \I__1370\ : Span4Mux_v
    port map (
            O => \N__5987\,
            I => \N__5965\
        );

    \I__1369\ : Span4Mux_h
    port map (
            O => \N__5984\,
            I => \N__5960\
        );

    \I__1368\ : Span4Mux_v
    port map (
            O => \N__5975\,
            I => \N__5960\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__5972\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1366\ : Odrv4
    port map (
            O => \N__5965\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1365\ : Odrv4
    port map (
            O => \N__5960\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1364\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5950\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__5950\,
            I => \U400_SDRAM.MAc_9_0\
        );

    \I__1362\ : IoInMux
    port map (
            O => \N__5947\,
            I => \N__5944\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__5944\,
            I => \MA_c_1\
        );

    \I__1360\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5938\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__5938\,
            I => \N__5929\
        );

    \I__1358\ : SRMux
    port map (
            O => \N__5937\,
            I => \N__5887\
        );

    \I__1357\ : SRMux
    port map (
            O => \N__5936\,
            I => \N__5887\
        );

    \I__1356\ : SRMux
    port map (
            O => \N__5935\,
            I => \N__5887\
        );

    \I__1355\ : SRMux
    port map (
            O => \N__5934\,
            I => \N__5887\
        );

    \I__1354\ : SRMux
    port map (
            O => \N__5933\,
            I => \N__5887\
        );

    \I__1353\ : SRMux
    port map (
            O => \N__5932\,
            I => \N__5887\
        );

    \I__1352\ : Glb2LocalMux
    port map (
            O => \N__5929\,
            I => \N__5887\
        );

    \I__1351\ : SRMux
    port map (
            O => \N__5928\,
            I => \N__5887\
        );

    \I__1350\ : SRMux
    port map (
            O => \N__5927\,
            I => \N__5887\
        );

    \I__1349\ : SRMux
    port map (
            O => \N__5926\,
            I => \N__5887\
        );

    \I__1348\ : SRMux
    port map (
            O => \N__5925\,
            I => \N__5887\
        );

    \I__1347\ : SRMux
    port map (
            O => \N__5924\,
            I => \N__5887\
        );

    \I__1346\ : SRMux
    port map (
            O => \N__5923\,
            I => \N__5887\
        );

    \I__1345\ : SRMux
    port map (
            O => \N__5922\,
            I => \N__5887\
        );

    \I__1344\ : SRMux
    port map (
            O => \N__5921\,
            I => \N__5887\
        );

    \I__1343\ : SRMux
    port map (
            O => \N__5920\,
            I => \N__5887\
        );

    \I__1342\ : GlobalMux
    port map (
            O => \N__5887\,
            I => \N__5884\
        );

    \I__1341\ : gio2CtrlBuf
    port map (
            O => \N__5884\,
            I => \RESETn_c_i_g\
        );

    \I__1340\ : IoInMux
    port map (
            O => \N__5881\,
            I => \N__5878\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__5878\,
            I => \MA_c_10\
        );

    \I__1338\ : IoInMux
    port map (
            O => \N__5875\,
            I => \N__5872\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__5872\,
            I => \N__5869\
        );

    \I__1336\ : Odrv12
    port map (
            O => \N__5869\,
            I => \UMBEn_c\
        );

    \I__1335\ : IoInMux
    port map (
            O => \N__5866\,
            I => \N__5863\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__5863\,
            I => \N__5860\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__5860\,
            I => \LLBEn_c\
        );

    \I__1332\ : CascadeMux
    port map (
            O => \N__5857\,
            I => \N__5853\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__5856\,
            I => \N__5850\
        );

    \I__1330\ : InMux
    port map (
            O => \N__5853\,
            I => \N__5842\
        );

    \I__1329\ : InMux
    port map (
            O => \N__5850\,
            I => \N__5842\
        );

    \I__1328\ : InMux
    port map (
            O => \N__5849\,
            I => \N__5842\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__5842\,
            I => \N__5838\
        );

    \I__1326\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5835\
        );

    \I__1325\ : Span4Mux_h
    port map (
            O => \N__5838\,
            I => \N__5832\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__5835\,
            I => \N__5829\
        );

    \I__1323\ : Sp12to4
    port map (
            O => \N__5832\,
            I => \N__5824\
        );

    \I__1322\ : Sp12to4
    port map (
            O => \N__5829\,
            I => \N__5824\
        );

    \I__1321\ : Span12Mux_v
    port map (
            O => \N__5824\,
            I => \N__5821\
        );

    \I__1320\ : Odrv12
    port map (
            O => \N__5821\,
            I => \A_c_1\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__5818\,
            I => \N__5813\
        );

    \I__1318\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5805\
        );

    \I__1317\ : InMux
    port map (
            O => \N__5816\,
            I => \N__5805\
        );

    \I__1316\ : InMux
    port map (
            O => \N__5813\,
            I => \N__5805\
        );

    \I__1315\ : InMux
    port map (
            O => \N__5812\,
            I => \N__5802\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__5805\,
            I => \N__5797\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5802\,
            I => \N__5797\
        );

    \I__1312\ : Span4Mux_h
    port map (
            O => \N__5797\,
            I => \N__5794\
        );

    \I__1311\ : Sp12to4
    port map (
            O => \N__5794\,
            I => \N__5791\
        );

    \I__1310\ : Span12Mux_v
    port map (
            O => \N__5791\,
            I => \N__5788\
        );

    \I__1309\ : Odrv12
    port map (
            O => \N__5788\,
            I => \A_c_0\
        );

    \I__1308\ : IoInMux
    port map (
            O => \N__5785\,
            I => \N__5782\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__5782\,
            I => \N__5779\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__5779\,
            I => \LMBEn_c\
        );

    \I__1305\ : InMux
    port map (
            O => \N__5776\,
            I => \N__5773\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__5773\,
            I => \N__5770\
        );

    \I__1303\ : Span4Mux_v
    port map (
            O => \N__5770\,
            I => \N__5767\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__5767\,
            I => \TSn_c\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5764\,
            I => \N__5761\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__5761\,
            I => \N__5758\
        );

    \I__1299\ : Span4Mux_h
    port map (
            O => \N__5758\,
            I => \N__5755\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__5755\,
            I => \U400_SDRAM.N_220\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__5752\,
            I => \N__5748\
        );

    \I__1296\ : InMux
    port map (
            O => \N__5751\,
            I => \N__5745\
        );

    \I__1295\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5738\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__5745\,
            I => \N__5735\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5744\,
            I => \N__5728\
        );

    \I__1292\ : InMux
    port map (
            O => \N__5743\,
            I => \N__5728\
        );

    \I__1291\ : InMux
    port map (
            O => \N__5742\,
            I => \N__5728\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5741\,
            I => \N__5725\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5738\,
            I => \N__5721\
        );

    \I__1288\ : Span4Mux_v
    port map (
            O => \N__5735\,
            I => \N__5718\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__5728\,
            I => \N__5715\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__5725\,
            I => \N__5712\
        );

    \I__1285\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5709\
        );

    \I__1284\ : Span4Mux_h
    port map (
            O => \N__5721\,
            I => \N__5706\
        );

    \I__1283\ : Span4Mux_h
    port map (
            O => \N__5718\,
            I => \N__5697\
        );

    \I__1282\ : Span4Mux_v
    port map (
            O => \N__5715\,
            I => \N__5697\
        );

    \I__1281\ : Span4Mux_v
    port map (
            O => \N__5712\,
            I => \N__5697\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__5709\,
            I => \N__5697\
        );

    \I__1279\ : Span4Mux_v
    port map (
            O => \N__5706\,
            I => \N__5694\
        );

    \I__1278\ : IoSpan4Mux
    port map (
            O => \N__5697\,
            I => \N__5691\
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__5694\,
            I => \SIZ_c_1\
        );

    \I__1276\ : Odrv4
    port map (
            O => \N__5691\,
            I => \SIZ_c_1\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__5686\,
            I => \N__5682\
        );

    \I__1274\ : InMux
    port map (
            O => \N__5685\,
            I => \N__5676\
        );

    \I__1273\ : InMux
    port map (
            O => \N__5682\,
            I => \N__5672\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5681\,
            I => \N__5665\
        );

    \I__1271\ : InMux
    port map (
            O => \N__5680\,
            I => \N__5665\
        );

    \I__1270\ : InMux
    port map (
            O => \N__5679\,
            I => \N__5665\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__5676\,
            I => \N__5661\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5675\,
            I => \N__5658\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__5672\,
            I => \N__5655\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__5665\,
            I => \N__5652\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5649\
        );

    \I__1264\ : Sp12to4
    port map (
            O => \N__5661\,
            I => \N__5646\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5658\,
            I => \N__5643\
        );

    \I__1262\ : Span4Mux_v
    port map (
            O => \N__5655\,
            I => \N__5640\
        );

    \I__1261\ : Span4Mux_s3_v
    port map (
            O => \N__5652\,
            I => \N__5635\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__5649\,
            I => \N__5635\
        );

    \I__1259\ : Span12Mux_s7_v
    port map (
            O => \N__5646\,
            I => \N__5632\
        );

    \I__1258\ : Span4Mux_v
    port map (
            O => \N__5643\,
            I => \N__5629\
        );

    \I__1257\ : Span4Mux_h
    port map (
            O => \N__5640\,
            I => \N__5624\
        );

    \I__1256\ : Span4Mux_v
    port map (
            O => \N__5635\,
            I => \N__5624\
        );

    \I__1255\ : Odrv12
    port map (
            O => \N__5632\,
            I => \SIZ_c_0\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__5629\,
            I => \SIZ_c_0\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__5624\,
            I => \SIZ_c_0\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5614\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__5614\,
            I => \N__5610\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__5613\,
            I => \N__5607\
        );

    \I__1249\ : Span4Mux_v
    port map (
            O => \N__5610\,
            I => \N__5604\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5607\,
            I => \N__5601\
        );

    \I__1247\ : Odrv4
    port map (
            O => \N__5604\,
            I => \U400_SDRAM.BURST8\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__5601\,
            I => \U400_SDRAM.BURST8\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5590\
        );

    \I__1244\ : InMux
    port map (
            O => \N__5595\,
            I => \N__5590\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__5590\,
            I => \N__5587\
        );

    \I__1242\ : Span4Mux_h
    port map (
            O => \N__5587\,
            I => \N__5584\
        );

    \I__1241\ : Span4Mux_h
    port map (
            O => \N__5584\,
            I => \N__5581\
        );

    \I__1240\ : Span4Mux_v
    port map (
            O => \N__5581\,
            I => \N__5578\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__5578\,
            I => \A_c_31\
        );

    \I__1238\ : CascadeMux
    port map (
            O => \N__5575\,
            I => \N__5572\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5572\,
            I => \N__5566\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5571\,
            I => \N__5566\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__5566\,
            I => \N__5563\
        );

    \I__1234\ : Span12Mux_v
    port map (
            O => \N__5563\,
            I => \N__5560\
        );

    \I__1233\ : Odrv12
    port map (
            O => \N__5560\,
            I => \U400_ADDRESS_DECODE_RAM_SPACE_0_a3_3\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__5557\,
            I => \N__5548\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5545\
        );

    \I__1230\ : InMux
    port map (
            O => \N__5555\,
            I => \N__5542\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__5554\,
            I => \N__5538\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__5553\,
            I => \N__5535\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5552\,
            I => \N__5528\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5551\,
            I => \N__5528\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5548\,
            I => \N__5528\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5545\,
            I => \N__5519\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5542\,
            I => \N__5516\
        );

    \I__1222\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5513\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5538\,
            I => \N__5510\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5507\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5528\,
            I => \N__5504\
        );

    \I__1218\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5499\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5526\,
            I => \N__5499\
        );

    \I__1216\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5494\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5494\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5491\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5485\
        );

    \I__1212\ : Span4Mux_v
    port map (
            O => \N__5519\,
            I => \N__5482\
        );

    \I__1211\ : Span4Mux_v
    port map (
            O => \N__5516\,
            I => \N__5479\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__5513\,
            I => \N__5474\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__5510\,
            I => \N__5474\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__5507\,
            I => \N__5471\
        );

    \I__1207\ : Span4Mux_h
    port map (
            O => \N__5504\,
            I => \N__5464\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__5499\,
            I => \N__5464\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__5494\,
            I => \N__5464\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__5491\,
            I => \N__5461\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5456\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5456\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5453\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5485\,
            I => \N__5450\
        );

    \I__1199\ : Span4Mux_v
    port map (
            O => \N__5482\,
            I => \N__5443\
        );

    \I__1198\ : Span4Mux_h
    port map (
            O => \N__5479\,
            I => \N__5443\
        );

    \I__1197\ : Span4Mux_v
    port map (
            O => \N__5474\,
            I => \N__5443\
        );

    \I__1196\ : Span4Mux_v
    port map (
            O => \N__5471\,
            I => \N__5440\
        );

    \I__1195\ : Span4Mux_v
    port map (
            O => \N__5464\,
            I => \N__5437\
        );

    \I__1194\ : Span4Mux_h
    port map (
            O => \N__5461\,
            I => \N__5432\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5456\,
            I => \N__5432\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5453\,
            I => \N__5429\
        );

    \I__1191\ : Span12Mux_s8_v
    port map (
            O => \N__5450\,
            I => \N__5426\
        );

    \I__1190\ : Span4Mux_h
    port map (
            O => \N__5443\,
            I => \N__5423\
        );

    \I__1189\ : Span4Mux_h
    port map (
            O => \N__5440\,
            I => \N__5418\
        );

    \I__1188\ : Span4Mux_h
    port map (
            O => \N__5437\,
            I => \N__5418\
        );

    \I__1187\ : Span4Mux_v
    port map (
            O => \N__5432\,
            I => \N__5413\
        );

    \I__1186\ : Span4Mux_v
    port map (
            O => \N__5429\,
            I => \N__5413\
        );

    \I__1185\ : Odrv12
    port map (
            O => \N__5426\,
            I => \RESETn_c\
        );

    \I__1184\ : Odrv4
    port map (
            O => \N__5423\,
            I => \RESETn_c\
        );

    \I__1183\ : Odrv4
    port map (
            O => \N__5418\,
            I => \RESETn_c\
        );

    \I__1182\ : Odrv4
    port map (
            O => \N__5413\,
            I => \RESETn_c\
        );

    \I__1181\ : IoInMux
    port map (
            O => \N__5404\,
            I => \N__5401\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__5401\,
            I => \N__5398\
        );

    \I__1179\ : Odrv12
    port map (
            O => \N__5398\,
            I => \N_220_3_i\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5392\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__5392\,
            I => \N__5389\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__5389\,
            I => \A_c_5\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__5386\,
            I => \N__5383\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5383\,
            I => \N__5380\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5380\,
            I => \N__5377\
        );

    \I__1172\ : Span4Mux_v
    port map (
            O => \N__5377\,
            I => \N__5374\
        );

    \I__1171\ : Odrv4
    port map (
            O => \N__5374\,
            I => \A_c_13\
        );

    \I__1170\ : IoInMux
    port map (
            O => \N__5371\,
            I => \N__5368\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__5368\,
            I => \N__5365\
        );

    \I__1168\ : Span12Mux_s3_v
    port map (
            O => \N__5365\,
            I => \N__5362\
        );

    \I__1167\ : Odrv12
    port map (
            O => \N__5362\,
            I => \MA_c_3\
        );

    \I__1166\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5356\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5356\,
            I => \N__5353\
        );

    \I__1164\ : Span4Mux_h
    port map (
            O => \N__5353\,
            I => \N__5350\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__5350\,
            I => \A_c_3\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__5347\,
            I => \N__5344\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5344\,
            I => \N__5341\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5341\,
            I => \N__5338\
        );

    \I__1159\ : Odrv4
    port map (
            O => \N__5338\,
            I => \A_c_11\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__5335\,
            I => \N__5331\
        );

    \I__1157\ : InMux
    port map (
            O => \N__5334\,
            I => \N__5328\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5331\,
            I => \N__5325\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__5328\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5325\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1153\ : CEMux
    port map (
            O => \N__5320\,
            I => \N__5316\
        );

    \I__1152\ : CEMux
    port map (
            O => \N__5319\,
            I => \N__5311\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5316\,
            I => \N__5308\
        );

    \I__1150\ : CEMux
    port map (
            O => \N__5315\,
            I => \N__5305\
        );

    \I__1149\ : CEMux
    port map (
            O => \N__5314\,
            I => \N__5302\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__5311\,
            I => \N__5299\
        );

    \I__1147\ : Span4Mux_v
    port map (
            O => \N__5308\,
            I => \N__5294\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5305\,
            I => \N__5294\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5302\,
            I => \N__5291\
        );

    \I__1144\ : Span4Mux_v
    port map (
            O => \N__5299\,
            I => \N__5286\
        );

    \I__1143\ : Span4Mux_h
    port map (
            O => \N__5294\,
            I => \N__5286\
        );

    \I__1142\ : Odrv12
    port map (
            O => \N__5291\,
            I => \U400_SDRAM.SDRAM_COUNTERe_0_i\
        );

    \I__1141\ : Odrv4
    port map (
            O => \N__5286\,
            I => \U400_SDRAM.SDRAM_COUNTERe_0_i\
        );

    \I__1140\ : CascadeMux
    port map (
            O => \N__5281\,
            I => \N__5277\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5280\,
            I => \N__5263\
        );

    \I__1138\ : InMux
    port map (
            O => \N__5277\,
            I => \N__5260\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5257\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5252\
        );

    \I__1135\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5252\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5243\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5243\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5271\,
            I => \N__5243\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5270\,
            I => \N__5243\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5237\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5233\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5229\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5226\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5263\,
            I => \N__5220\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__5260\,
            I => \N__5220\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5257\,
            I => \N__5213\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__5252\,
            I => \N__5213\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__5243\,
            I => \N__5213\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5242\,
            I => \N__5210\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5205\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5240\,
            I => \N__5205\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5237\,
            I => \N__5202\
        );

    \I__1117\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5199\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5233\,
            I => \N__5196\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5193\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__5229\,
            I => \N__5188\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__5226\,
            I => \N__5188\
        );

    \I__1112\ : InMux
    port map (
            O => \N__5225\,
            I => \N__5185\
        );

    \I__1111\ : Span4Mux_v
    port map (
            O => \N__5220\,
            I => \N__5178\
        );

    \I__1110\ : Span4Mux_v
    port map (
            O => \N__5213\,
            I => \N__5178\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__5210\,
            I => \N__5178\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__5205\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1107\ : Odrv12
    port map (
            O => \N__5202\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__5199\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1105\ : Odrv4
    port map (
            O => \N__5196\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5193\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1103\ : Odrv12
    port map (
            O => \N__5188\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5185\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1101\ : Odrv4
    port map (
            O => \N__5178\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__5161\,
            I => \N__5156\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__5160\,
            I => \N__5153\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__5159\,
            I => \N__5146\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5143\
        );

    \I__1096\ : InMux
    port map (
            O => \N__5153\,
            I => \N__5139\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__5152\,
            I => \N__5136\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__5151\,
            I => \N__5132\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__5150\,
            I => \N__5128\
        );

    \I__1092\ : InMux
    port map (
            O => \N__5149\,
            I => \N__5122\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5146\,
            I => \N__5122\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__5143\,
            I => \N__5119\
        );

    \I__1089\ : InMux
    port map (
            O => \N__5142\,
            I => \N__5116\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5139\,
            I => \N__5113\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5136\,
            I => \N__5110\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5135\,
            I => \N__5103\
        );

    \I__1085\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5103\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5131\,
            I => \N__5103\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5128\,
            I => \N__5098\
        );

    \I__1082\ : InMux
    port map (
            O => \N__5127\,
            I => \N__5098\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__5122\,
            I => \N__5093\
        );

    \I__1080\ : Span4Mux_v
    port map (
            O => \N__5119\,
            I => \N__5093\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__5116\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__1078\ : Odrv4
    port map (
            O => \N__5113\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5110\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5103\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__5098\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__1074\ : Odrv4
    port map (
            O => \N__5093\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5080\,
            I => \N__5065\
        );

    \I__1072\ : InMux
    port map (
            O => \N__5079\,
            I => \N__5065\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5065\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5062\
        );

    \I__1069\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5059\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__5075\,
            I => \N__5056\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__5074\,
            I => \N__5053\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5050\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5072\,
            I => \N__5047\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__5065\,
            I => \N__5044\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__5062\,
            I => \N__5033\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__5059\,
            I => \N__5033\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5056\,
            I => \N__5028\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5053\,
            I => \N__5028\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5050\,
            I => \N__5023\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__5047\,
            I => \N__5023\
        );

    \I__1057\ : Span4Mux_h
    port map (
            O => \N__5044\,
            I => \N__5018\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5013\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5042\,
            I => \N__5013\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5010\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5007\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5004\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5001\
        );

    \I__1050\ : Span4Mux_h
    port map (
            O => \N__5033\,
            I => \N__4994\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__5028\,
            I => \N__4994\
        );

    \I__1048\ : Span4Mux_h
    port map (
            O => \N__5023\,
            I => \N__4994\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5022\,
            I => \N__4989\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5021\,
            I => \N__4989\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__5018\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__5013\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5010\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5007\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5004\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5001\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1039\ : Odrv4
    port map (
            O => \N__4994\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__4989\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__4972\,
            I => \U400_SDRAM.N_161_cascade_\
        );

    \I__1036\ : InMux
    port map (
            O => \N__4969\,
            I => \N__4966\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__4966\,
            I => \U400_SDRAM.N_183\
        );

    \I__1034\ : InMux
    port map (
            O => \N__4963\,
            I => \N__4952\
        );

    \I__1033\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4952\
        );

    \I__1032\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4952\
        );

    \I__1031\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4941\
        );

    \I__1030\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4941\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__4952\,
            I => \N__4935\
        );

    \I__1028\ : InMux
    port map (
            O => \N__4951\,
            I => \N__4930\
        );

    \I__1027\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4930\
        );

    \I__1026\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4923\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4948\,
            I => \N__4920\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4947\,
            I => \N__4917\
        );

    \I__1023\ : InMux
    port map (
            O => \N__4946\,
            I => \N__4914\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__4941\,
            I => \N__4911\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4940\,
            I => \N__4908\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4939\,
            I => \N__4903\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4903\
        );

    \I__1018\ : Span4Mux_h
    port map (
            O => \N__4935\,
            I => \N__4898\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__4930\,
            I => \N__4898\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4929\,
            I => \N__4895\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4888\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4888\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4888\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__4923\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4920\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4917\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__4914\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1008\ : Odrv12
    port map (
            O => \N__4911\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4908\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4903\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__4898\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__4895\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__4888\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4863\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4859\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4863\,
            I => \N__4856\
        );

    \I__999\ : InMux
    port map (
            O => \N__4862\,
            I => \N__4851\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__4859\,
            I => \N__4848\
        );

    \I__997\ : Span4Mux_h
    port map (
            O => \N__4856\,
            I => \N__4845\
        );

    \I__996\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4842\
        );

    \I__995\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4839\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4851\,
            I => \U400_SDRAM.N_126\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__4848\,
            I => \U400_SDRAM.N_126\
        );

    \I__992\ : Odrv4
    port map (
            O => \N__4845\,
            I => \U400_SDRAM.N_126\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__4842\,
            I => \U400_SDRAM.N_126\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__4839\,
            I => \U400_SDRAM.N_126\
        );

    \I__989\ : CascadeMux
    port map (
            O => \N__4828\,
            I => \N__4821\
        );

    \I__988\ : InMux
    port map (
            O => \N__4827\,
            I => \N__4818\
        );

    \I__987\ : InMux
    port map (
            O => \N__4826\,
            I => \N__4815\
        );

    \I__986\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4812\
        );

    \I__985\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4809\
        );

    \I__984\ : InMux
    port map (
            O => \N__4821\,
            I => \N__4806\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4818\,
            I => \N__4799\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4815\,
            I => \N__4796\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4812\,
            I => \N__4789\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4809\,
            I => \N__4789\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4806\,
            I => \N__4789\
        );

    \I__978\ : InMux
    port map (
            O => \N__4805\,
            I => \N__4786\
        );

    \I__977\ : InMux
    port map (
            O => \N__4804\,
            I => \N__4781\
        );

    \I__976\ : InMux
    port map (
            O => \N__4803\,
            I => \N__4781\
        );

    \I__975\ : InMux
    port map (
            O => \N__4802\,
            I => \N__4775\
        );

    \I__974\ : Span4Mux_h
    port map (
            O => \N__4799\,
            I => \N__4772\
        );

    \I__973\ : Span4Mux_v
    port map (
            O => \N__4796\,
            I => \N__4767\
        );

    \I__972\ : Span4Mux_v
    port map (
            O => \N__4789\,
            I => \N__4767\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4786\,
            I => \N__4762\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4781\,
            I => \N__4762\
        );

    \I__969\ : InMux
    port map (
            O => \N__4780\,
            I => \N__4757\
        );

    \I__968\ : InMux
    port map (
            O => \N__4779\,
            I => \N__4757\
        );

    \I__967\ : InMux
    port map (
            O => \N__4778\,
            I => \N__4754\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4775\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__965\ : Odrv4
    port map (
            O => \N__4772\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__964\ : Odrv4
    port map (
            O => \N__4767\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__963\ : Odrv4
    port map (
            O => \N__4762\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__4757\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4754\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__960\ : InMux
    port map (
            O => \N__4741\,
            I => \N__4738\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4738\,
            I => \N__4735\
        );

    \I__958\ : Span4Mux_v
    port map (
            O => \N__4735\,
            I => \N__4731\
        );

    \I__957\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4728\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__4731\,
            I => \U400_SDRAM.N_138\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4728\,
            I => \U400_SDRAM.N_138\
        );

    \I__954\ : CascadeMux
    port map (
            O => \N__4723\,
            I => \N__4720\
        );

    \I__953\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4717\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4717\,
            I => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a3_1_0_0\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__4714\,
            I => \N__4703\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__4713\,
            I => \N__4700\
        );

    \I__949\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4697\
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__4711\,
            I => \N__4694\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__4710\,
            I => \N__4691\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__4709\,
            I => \N__4688\
        );

    \I__945\ : CascadeMux
    port map (
            O => \N__4708\,
            I => \N__4685\
        );

    \I__944\ : CascadeMux
    port map (
            O => \N__4707\,
            I => \N__4681\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__4706\,
            I => \N__4677\
        );

    \I__942\ : InMux
    port map (
            O => \N__4703\,
            I => \N__4674\
        );

    \I__941\ : InMux
    port map (
            O => \N__4700\,
            I => \N__4671\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4697\,
            I => \N__4668\
        );

    \I__939\ : InMux
    port map (
            O => \N__4694\,
            I => \N__4661\
        );

    \I__938\ : InMux
    port map (
            O => \N__4691\,
            I => \N__4661\
        );

    \I__937\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4661\
        );

    \I__936\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4654\
        );

    \I__935\ : InMux
    port map (
            O => \N__4684\,
            I => \N__4654\
        );

    \I__934\ : InMux
    port map (
            O => \N__4681\,
            I => \N__4647\
        );

    \I__933\ : InMux
    port map (
            O => \N__4680\,
            I => \N__4647\
        );

    \I__932\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4647\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4674\,
            I => \N__4642\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4671\,
            I => \N__4642\
        );

    \I__929\ : Span4Mux_v
    port map (
            O => \N__4668\,
            I => \N__4635\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4661\,
            I => \N__4635\
        );

    \I__927\ : InMux
    port map (
            O => \N__4660\,
            I => \N__4630\
        );

    \I__926\ : InMux
    port map (
            O => \N__4659\,
            I => \N__4630\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4654\,
            I => \N__4622\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4647\,
            I => \N__4622\
        );

    \I__923\ : Span4Mux_h
    port map (
            O => \N__4642\,
            I => \N__4619\
        );

    \I__922\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4616\
        );

    \I__921\ : InMux
    port map (
            O => \N__4640\,
            I => \N__4613\
        );

    \I__920\ : Span4Mux_h
    port map (
            O => \N__4635\,
            I => \N__4608\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__4630\,
            I => \N__4608\
        );

    \I__918\ : InMux
    port map (
            O => \N__4629\,
            I => \N__4603\
        );

    \I__917\ : InMux
    port map (
            O => \N__4628\,
            I => \N__4603\
        );

    \I__916\ : InMux
    port map (
            O => \N__4627\,
            I => \N__4600\
        );

    \I__915\ : Span4Mux_v
    port map (
            O => \N__4622\,
            I => \N__4597\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__4619\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4616\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__4613\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__911\ : Odrv4
    port map (
            O => \N__4608\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4603\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__4600\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__4597\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__4582\,
            I => \N__4578\
        );

    \I__906\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4573\
        );

    \I__905\ : InMux
    port map (
            O => \N__4578\,
            I => \N__4570\
        );

    \I__904\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4567\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__4576\,
            I => \N__4562\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4573\,
            I => \N__4559\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4570\,
            I => \N__4556\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4567\,
            I => \N__4553\
        );

    \I__899\ : InMux
    port map (
            O => \N__4566\,
            I => \N__4548\
        );

    \I__898\ : InMux
    port map (
            O => \N__4565\,
            I => \N__4548\
        );

    \I__897\ : InMux
    port map (
            O => \N__4562\,
            I => \N__4545\
        );

    \I__896\ : Span4Mux_h
    port map (
            O => \N__4559\,
            I => \N__4542\
        );

    \I__895\ : Span4Mux_h
    port map (
            O => \N__4556\,
            I => \N__4533\
        );

    \I__894\ : Span4Mux_h
    port map (
            O => \N__4553\,
            I => \N__4533\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4548\,
            I => \N__4533\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4545\,
            I => \N__4533\
        );

    \I__891\ : Odrv4
    port map (
            O => \N__4542\,
            I => \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7JZ0\
        );

    \I__890\ : Odrv4
    port map (
            O => \N__4533\,
            I => \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7JZ0\
        );

    \I__889\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4525\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4525\,
            I => \N__4522\
        );

    \I__887\ : Span4Mux_s2_v
    port map (
            O => \N__4522\,
            I => \N__4519\
        );

    \I__886\ : Odrv4
    port map (
            O => \N__4519\,
            I => \A_c_7\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__4516\,
            I => \N__4513\
        );

    \I__884\ : InMux
    port map (
            O => \N__4513\,
            I => \N__4510\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__4510\,
            I => \N__4507\
        );

    \I__882\ : IoSpan4Mux
    port map (
            O => \N__4507\,
            I => \N__4504\
        );

    \I__881\ : Odrv4
    port map (
            O => \N__4504\,
            I => \A_c_15\
        );

    \I__880\ : InMux
    port map (
            O => \N__4501\,
            I => \N__4498\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4498\,
            I => \U400_SDRAM.MAc_0_0\
        );

    \I__878\ : InMux
    port map (
            O => \N__4495\,
            I => \N__4492\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__4492\,
            I => \N__4489\
        );

    \I__876\ : Span4Mux_h
    port map (
            O => \N__4489\,
            I => \N__4486\
        );

    \I__875\ : Odrv4
    port map (
            O => \N__4486\,
            I => \A_c_2\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__4483\,
            I => \N__4480\
        );

    \I__873\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4477\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4477\,
            I => \N__4474\
        );

    \I__871\ : Span4Mux_s1_v
    port map (
            O => \N__4474\,
            I => \N__4471\
        );

    \I__870\ : Odrv4
    port map (
            O => \N__4471\,
            I => \A_c_10\
        );

    \I__869\ : IoInMux
    port map (
            O => \N__4468\,
            I => \N__4465\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4465\,
            I => \MA_c_0\
        );

    \I__867\ : InMux
    port map (
            O => \N__4462\,
            I => \N__4459\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4459\,
            I => \N__4456\
        );

    \I__865\ : Span12Mux_s10_h
    port map (
            O => \N__4456\,
            I => \N__4453\
        );

    \I__864\ : Span12Mux_v
    port map (
            O => \N__4453\,
            I => \N__4450\
        );

    \I__863\ : Odrv12
    port map (
            O => \N__4450\,
            I => \A_c_20\
        );

    \I__862\ : InMux
    port map (
            O => \N__4447\,
            I => \N__4444\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4444\,
            I => \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5Z0Z_0\
        );

    \I__860\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4438\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4438\,
            I => \N__4435\
        );

    \I__858\ : Span4Mux_h
    port map (
            O => \N__4435\,
            I => \N__4428\
        );

    \I__857\ : InMux
    port map (
            O => \N__4434\,
            I => \N__4425\
        );

    \I__856\ : InMux
    port map (
            O => \N__4433\,
            I => \N__4422\
        );

    \I__855\ : InMux
    port map (
            O => \N__4432\,
            I => \N__4419\
        );

    \I__854\ : InMux
    port map (
            O => \N__4431\,
            I => \N__4416\
        );

    \I__853\ : Odrv4
    port map (
            O => \N__4428\,
            I => \U400_SDRAM.N_129\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__4425\,
            I => \U400_SDRAM.N_129\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4422\,
            I => \U400_SDRAM.N_129\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4419\,
            I => \U400_SDRAM.N_129\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4416\,
            I => \U400_SDRAM.N_129\
        );

    \I__848\ : InMux
    port map (
            O => \N__4405\,
            I => \N__4401\
        );

    \I__847\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4397\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4401\,
            I => \N__4394\
        );

    \I__845\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4391\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4397\,
            I => \U400_SDRAM.N_260\
        );

    \I__843\ : Odrv4
    port map (
            O => \N__4394\,
            I => \U400_SDRAM.N_260\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4391\,
            I => \U400_SDRAM.N_260\
        );

    \I__841\ : InMux
    port map (
            O => \N__4384\,
            I => \N__4381\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4381\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_1\
        );

    \I__839\ : InMux
    port map (
            O => \N__4378\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_0\
        );

    \I__838\ : InMux
    port map (
            O => \N__4375\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_1\
        );

    \I__837\ : InMux
    port map (
            O => \N__4372\,
            I => \N__4369\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4369\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_3\
        );

    \I__835\ : InMux
    port map (
            O => \N__4366\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_2\
        );

    \I__834\ : InMux
    port map (
            O => \N__4363\,
            I => \N__4359\
        );

    \I__833\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4356\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4359\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4356\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__830\ : InMux
    port map (
            O => \N__4351\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_3\
        );

    \I__829\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4344\
        );

    \I__828\ : InMux
    port map (
            O => \N__4347\,
            I => \N__4341\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4344\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4341\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__825\ : InMux
    port map (
            O => \N__4336\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_4\
        );

    \I__824\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4329\
        );

    \I__823\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4326\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4329\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4326\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__820\ : InMux
    port map (
            O => \N__4321\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_5\
        );

    \I__819\ : InMux
    port map (
            O => \N__4318\,
            I => \N__4307\
        );

    \I__818\ : InMux
    port map (
            O => \N__4317\,
            I => \N__4307\
        );

    \I__817\ : InMux
    port map (
            O => \N__4316\,
            I => \N__4307\
        );

    \I__816\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4301\
        );

    \I__815\ : InMux
    port map (
            O => \N__4314\,
            I => \N__4298\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4307\,
            I => \N__4295\
        );

    \I__813\ : InMux
    port map (
            O => \N__4306\,
            I => \N__4292\
        );

    \I__812\ : InMux
    port map (
            O => \N__4305\,
            I => \N__4287\
        );

    \I__811\ : InMux
    port map (
            O => \N__4304\,
            I => \N__4287\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__4301\,
            I => \U400_SDRAM.N_37\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4298\,
            I => \U400_SDRAM.N_37\
        );

    \I__808\ : Odrv4
    port map (
            O => \N__4295\,
            I => \U400_SDRAM.N_37\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4292\,
            I => \U400_SDRAM.N_37\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4287\,
            I => \U400_SDRAM.N_37\
        );

    \I__805\ : InMux
    port map (
            O => \N__4276\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_6\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__4273\,
            I => \N__4270\
        );

    \I__803\ : InMux
    port map (
            O => \N__4270\,
            I => \N__4267\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__4267\,
            I => \N__4264\
        );

    \I__801\ : Span12Mux_v
    port map (
            O => \N__4264\,
            I => \N__4261\
        );

    \I__800\ : Odrv12
    port map (
            O => \N__4261\,
            I => \A_c_25\
        );

    \I__799\ : IoInMux
    port map (
            O => \N__4258\,
            I => \N__4255\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4255\,
            I => \N__4252\
        );

    \I__797\ : Span4Mux_s3_v
    port map (
            O => \N__4252\,
            I => \N__4249\
        );

    \I__796\ : Odrv4
    port map (
            O => \N__4249\,
            I => \MA_c_11\
        );

    \I__795\ : InMux
    port map (
            O => \N__4246\,
            I => \N__4243\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4243\,
            I => \N__4236\
        );

    \I__793\ : InMux
    port map (
            O => \N__4242\,
            I => \N__4233\
        );

    \I__792\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4230\
        );

    \I__791\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4225\
        );

    \I__790\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4225\
        );

    \I__789\ : Odrv4
    port map (
            O => \N__4236\,
            I => \U400_SDRAM.N_257\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4233\,
            I => \U400_SDRAM.N_257\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4230\,
            I => \U400_SDRAM.N_257\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4225\,
            I => \U400_SDRAM.N_257\
        );

    \I__785\ : InMux
    port map (
            O => \N__4216\,
            I => \N__4213\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4213\,
            I => \N__4210\
        );

    \I__783\ : Span4Mux_s3_v
    port map (
            O => \N__4210\,
            I => \N__4207\
        );

    \I__782\ : Span4Mux_h
    port map (
            O => \N__4207\,
            I => \N__4204\
        );

    \I__781\ : Odrv4
    port map (
            O => \N__4204\,
            I => \A_c_6\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__4201\,
            I => \N__4198\
        );

    \I__779\ : InMux
    port map (
            O => \N__4198\,
            I => \N__4195\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4195\,
            I => \N__4192\
        );

    \I__777\ : Span4Mux_h
    port map (
            O => \N__4192\,
            I => \N__4189\
        );

    \I__776\ : Odrv4
    port map (
            O => \N__4189\,
            I => \A_c_14\
        );

    \I__775\ : IoInMux
    port map (
            O => \N__4186\,
            I => \N__4183\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4183\,
            I => \N__4180\
        );

    \I__773\ : Span4Mux_s0_v
    port map (
            O => \N__4180\,
            I => \N__4177\
        );

    \I__772\ : Span4Mux_h
    port map (
            O => \N__4177\,
            I => \N__4174\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__4174\,
            I => \MA_c_4\
        );

    \I__770\ : IoInMux
    port map (
            O => \N__4171\,
            I => \N__4168\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4168\,
            I => \N__4165\
        );

    \I__768\ : IoSpan4Mux
    port map (
            O => \N__4165\,
            I => \N__4162\
        );

    \I__767\ : Odrv4
    port map (
            O => \N__4162\,
            I => \MA_c_5\
        );

    \I__766\ : InMux
    port map (
            O => \N__4159\,
            I => \N__4156\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__764\ : Odrv4
    port map (
            O => \N__4153\,
            I => \U400_SDRAM.N_150\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__4150\,
            I => \U400_SDRAM.N_150_cascade_\
        );

    \I__762\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4143\
        );

    \I__761\ : InMux
    port map (
            O => \N__4146\,
            I => \N__4140\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4143\,
            I => \U400_SDRAM.N_252\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4140\,
            I => \U400_SDRAM.N_252\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__4135\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_61_i_i_a3_1_0_cascade_\
        );

    \I__757\ : InMux
    port map (
            O => \N__4132\,
            I => \N__4126\
        );

    \I__756\ : InMux
    port map (
            O => \N__4131\,
            I => \N__4126\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4126\,
            I => \U400_SDRAM.N_201\
        );

    \I__754\ : InMux
    port map (
            O => \N__4123\,
            I => \N__4120\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4120\,
            I => \TA_EN_i_ess\
        );

    \I__752\ : IoInMux
    port map (
            O => \N__4117\,
            I => \N__4114\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4114\,
            I => \N__4111\
        );

    \I__750\ : Odrv12
    port map (
            O => \N__4111\,
            I => \N_529_i\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__4108\,
            I => \U400_SDRAM.N_126_cascade_\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__4105\,
            I => \U400_SDRAM.N_129_cascade_\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__4102\,
            I => \U400_SDRAM.N_257_cascade_\
        );

    \I__746\ : InMux
    port map (
            O => \N__4099\,
            I => \N__4096\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4096\,
            I => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_1_0\
        );

    \I__744\ : InMux
    port map (
            O => \N__4093\,
            I => \N__4088\
        );

    \I__743\ : InMux
    port map (
            O => \N__4092\,
            I => \N__4083\
        );

    \I__742\ : InMux
    port map (
            O => \N__4091\,
            I => \N__4083\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4088\,
            I => \U400_SDRAM.N_133\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4083\,
            I => \U400_SDRAM.N_133\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__4078\,
            I => \U400_SDRAM.N_133_cascade_\
        );

    \I__738\ : CascadeMux
    port map (
            O => \N__4075\,
            I => \N__4070\
        );

    \I__737\ : InMux
    port map (
            O => \N__4074\,
            I => \N__4060\
        );

    \I__736\ : InMux
    port map (
            O => \N__4073\,
            I => \N__4060\
        );

    \I__735\ : InMux
    port map (
            O => \N__4070\,
            I => \N__4055\
        );

    \I__734\ : InMux
    port map (
            O => \N__4069\,
            I => \N__4055\
        );

    \I__733\ : InMux
    port map (
            O => \N__4068\,
            I => \N__4052\
        );

    \I__732\ : InMux
    port map (
            O => \N__4067\,
            I => \N__4047\
        );

    \I__731\ : InMux
    port map (
            O => \N__4066\,
            I => \N__4047\
        );

    \I__730\ : InMux
    port map (
            O => \N__4065\,
            I => \N__4044\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__4060\,
            I => \U400_SDRAM.N_139\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4055\,
            I => \U400_SDRAM.N_139\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__4052\,
            I => \U400_SDRAM.N_139\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4047\,
            I => \U400_SDRAM.N_139\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4044\,
            I => \U400_SDRAM.N_139\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__4033\,
            I => \U400_SDRAM.N_141_cascade_\
        );

    \I__723\ : InMux
    port map (
            O => \N__4030\,
            I => \N__4023\
        );

    \I__722\ : InMux
    port map (
            O => \N__4029\,
            I => \N__4023\
        );

    \I__721\ : InMux
    port map (
            O => \N__4028\,
            I => \N__4020\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4023\,
            I => \N__4009\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__4020\,
            I => \N__4006\
        );

    \I__718\ : InMux
    port map (
            O => \N__4019\,
            I => \N__4003\
        );

    \I__717\ : InMux
    port map (
            O => \N__4018\,
            I => \N__3998\
        );

    \I__716\ : InMux
    port map (
            O => \N__4017\,
            I => \N__3998\
        );

    \I__715\ : InMux
    port map (
            O => \N__4016\,
            I => \N__3995\
        );

    \I__714\ : InMux
    port map (
            O => \N__4015\,
            I => \N__3988\
        );

    \I__713\ : InMux
    port map (
            O => \N__4014\,
            I => \N__3988\
        );

    \I__712\ : InMux
    port map (
            O => \N__4013\,
            I => \N__3988\
        );

    \I__711\ : InMux
    port map (
            O => \N__4012\,
            I => \N__3985\
        );

    \I__710\ : Span4Mux_h
    port map (
            O => \N__4009\,
            I => \N__3976\
        );

    \I__709\ : Span4Mux_v
    port map (
            O => \N__4006\,
            I => \N__3976\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4003\,
            I => \N__3976\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__3998\,
            I => \N__3976\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3995\,
            I => \U400_SDRAM.REFRESH_COUNTER_RNIVV903Z0Z_8\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3988\,
            I => \U400_SDRAM.REFRESH_COUNTER_RNIVV903Z0Z_8\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__3985\,
            I => \U400_SDRAM.REFRESH_COUNTER_RNIVV903Z0Z_8\
        );

    \I__703\ : Odrv4
    port map (
            O => \N__3976\,
            I => \U400_SDRAM.REFRESH_COUNTER_RNIVV903Z0Z_8\
        );

    \I__702\ : InMux
    port map (
            O => \N__3967\,
            I => \N__3960\
        );

    \I__701\ : InMux
    port map (
            O => \N__3966\,
            I => \N__3960\
        );

    \I__700\ : InMux
    port map (
            O => \N__3965\,
            I => \N__3955\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3960\,
            I => \N__3952\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__3959\,
            I => \N__3945\
        );

    \I__697\ : InMux
    port map (
            O => \N__3958\,
            I => \N__3941\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3955\,
            I => \N__3938\
        );

    \I__695\ : Span4Mux_h
    port map (
            O => \N__3952\,
            I => \N__3935\
        );

    \I__694\ : InMux
    port map (
            O => \N__3951\,
            I => \N__3930\
        );

    \I__693\ : InMux
    port map (
            O => \N__3950\,
            I => \N__3930\
        );

    \I__692\ : InMux
    port map (
            O => \N__3949\,
            I => \N__3927\
        );

    \I__691\ : InMux
    port map (
            O => \N__3948\,
            I => \N__3924\
        );

    \I__690\ : InMux
    port map (
            O => \N__3945\,
            I => \N__3919\
        );

    \I__689\ : InMux
    port map (
            O => \N__3944\,
            I => \N__3919\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3941\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__687\ : Odrv4
    port map (
            O => \N__3938\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__686\ : Odrv4
    port map (
            O => \N__3935\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__3930\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3927\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__3924\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__3919\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__681\ : InMux
    port map (
            O => \N__3904\,
            I => \N__3901\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3901\,
            I => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_2_0\
        );

    \I__679\ : InMux
    port map (
            O => \N__3898\,
            I => \N__3895\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3895\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_0\
        );

    \I__677\ : CascadeMux
    port map (
            O => \N__3892\,
            I => \U400_SDRAM.N_181_cascade_\
        );

    \I__676\ : CascadeMux
    port map (
            O => \N__3889\,
            I => \U400_SDRAM.N_200_cascade_\
        );

    \I__675\ : InMux
    port map (
            O => \N__3886\,
            I => \N__3883\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3883\,
            I => \N__3880\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__3880\,
            I => \U400_SDRAM.N_199\
        );

    \I__672\ : CascadeMux
    port map (
            O => \N__3877\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_61_i_i_1_cascade_\
        );

    \I__671\ : InMux
    port map (
            O => \N__3874\,
            I => \N__3870\
        );

    \I__670\ : InMux
    port map (
            O => \N__3873\,
            I => \N__3866\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3870\,
            I => \N__3863\
        );

    \I__668\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3860\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3866\,
            I => \U400_SDRAM.N_17\
        );

    \I__666\ : Odrv4
    port map (
            O => \N__3863\,
            I => \U400_SDRAM.N_17\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3860\,
            I => \U400_SDRAM.N_17\
        );

    \I__664\ : InMux
    port map (
            O => \N__3853\,
            I => \N__3850\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__3850\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_0_1_1\
        );

    \I__662\ : InMux
    port map (
            O => \N__3847\,
            I => \N__3842\
        );

    \I__661\ : InMux
    port map (
            O => \N__3846\,
            I => \N__3839\
        );

    \I__660\ : InMux
    port map (
            O => \N__3845\,
            I => \N__3836\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3842\,
            I => \U400_SDRAM.N_228\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3839\,
            I => \U400_SDRAM.N_228\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3836\,
            I => \U400_SDRAM.N_228\
        );

    \I__656\ : CascadeMux
    port map (
            O => \N__3829\,
            I => \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5Z0Z_0_cascade_\
        );

    \I__655\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3823\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3823\,
            I => \U400_SDRAM.N_203\
        );

    \I__653\ : InMux
    port map (
            O => \N__3820\,
            I => \N__3817\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3817\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_i_0\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__3814\,
            I => \U400_SDRAM.N_176_cascade_\
        );

    \I__650\ : CascadeMux
    port map (
            O => \N__3811\,
            I => \N__3808\
        );

    \I__649\ : InMux
    port map (
            O => \N__3808\,
            I => \N__3805\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__3805\,
            I => \N__3801\
        );

    \I__647\ : InMux
    port map (
            O => \N__3804\,
            I => \N__3798\
        );

    \I__646\ : Odrv4
    port map (
            O => \N__3801\,
            I => \U400_SDRAM.CS1_ENZ0\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3798\,
            I => \U400_SDRAM.CS1_ENZ0\
        );

    \I__644\ : IoInMux
    port map (
            O => \N__3793\,
            I => \N__3790\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__3790\,
            I => \N__3787\
        );

    \I__642\ : Odrv12
    port map (
            O => \N__3787\,
            I => \CS1n_c\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__3784\,
            I => \N__3781\
        );

    \I__640\ : InMux
    port map (
            O => \N__3781\,
            I => \N__3778\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__3778\,
            I => \N__3775\
        );

    \I__638\ : Span4Mux_h
    port map (
            O => \N__3775\,
            I => \N__3772\
        );

    \I__637\ : Span4Mux_v
    port map (
            O => \N__3772\,
            I => \N__3769\
        );

    \I__636\ : Span4Mux_v
    port map (
            O => \N__3769\,
            I => \N__3766\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__3766\,
            I => \A_c_26\
        );

    \I__634\ : IoInMux
    port map (
            O => \N__3763\,
            I => \N__3760\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3760\,
            I => \N__3757\
        );

    \I__632\ : Span12Mux_s0_v
    port map (
            O => \N__3757\,
            I => \N__3754\
        );

    \I__631\ : Odrv12
    port map (
            O => \N__3754\,
            I => \MA_c_12\
        );

    \I__630\ : IoInMux
    port map (
            O => \N__3751\,
            I => \N__3748\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3748\,
            I => \N__3745\
        );

    \I__628\ : IoSpan4Mux
    port map (
            O => \N__3745\,
            I => \N__3741\
        );

    \I__627\ : InMux
    port map (
            O => \N__3744\,
            I => \N__3738\
        );

    \I__626\ : Span4Mux_s2_h
    port map (
            O => \N__3741\,
            I => \N__3735\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3738\,
            I => \N__3732\
        );

    \I__624\ : Odrv4
    port map (
            O => \N__3735\,
            I => \CONSTANT_ONE_NET\
        );

    \I__623\ : Odrv4
    port map (
            O => \N__3732\,
            I => \CONSTANT_ONE_NET\
        );

    \I__622\ : IoInMux
    port map (
            O => \N__3727\,
            I => \N__3724\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3724\,
            I => \N__3721\
        );

    \I__620\ : Odrv12
    port map (
            O => \N__3721\,
            I => \UUBEn_c\
        );

    \I__619\ : InMux
    port map (
            O => \N__3718\,
            I => \N__3715\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3715\,
            I => \N__3709\
        );

    \I__617\ : InMux
    port map (
            O => \N__3714\,
            I => \N__3706\
        );

    \I__616\ : InMux
    port map (
            O => \N__3713\,
            I => \N__3701\
        );

    \I__615\ : InMux
    port map (
            O => \N__3712\,
            I => \N__3701\
        );

    \I__614\ : Span4Mux_h
    port map (
            O => \N__3709\,
            I => \N__3696\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3706\,
            I => \N__3696\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3701\,
            I => \U400_SDRAM.TA_COUNTER23\
        );

    \I__611\ : Odrv4
    port map (
            O => \N__3696\,
            I => \U400_SDRAM.TA_COUNTER23\
        );

    \I__610\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3688\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3688\,
            I => \N__3682\
        );

    \I__608\ : InMux
    port map (
            O => \N__3687\,
            I => \N__3676\
        );

    \I__607\ : InMux
    port map (
            O => \N__3686\,
            I => \N__3676\
        );

    \I__606\ : InMux
    port map (
            O => \N__3685\,
            I => \N__3672\
        );

    \I__605\ : Span4Mux_h
    port map (
            O => \N__3682\,
            I => \N__3669\
        );

    \I__604\ : InMux
    port map (
            O => \N__3681\,
            I => \N__3666\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3676\,
            I => \N__3663\
        );

    \I__602\ : InMux
    port map (
            O => \N__3675\,
            I => \N__3660\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3672\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__600\ : Odrv4
    port map (
            O => \N__3669\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3666\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__598\ : Odrv4
    port map (
            O => \N__3663\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3660\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__596\ : ClkMux
    port map (
            O => \N__3649\,
            I => \N__3568\
        );

    \I__595\ : ClkMux
    port map (
            O => \N__3648\,
            I => \N__3568\
        );

    \I__594\ : ClkMux
    port map (
            O => \N__3647\,
            I => \N__3568\
        );

    \I__593\ : ClkMux
    port map (
            O => \N__3646\,
            I => \N__3568\
        );

    \I__592\ : ClkMux
    port map (
            O => \N__3645\,
            I => \N__3568\
        );

    \I__591\ : ClkMux
    port map (
            O => \N__3644\,
            I => \N__3568\
        );

    \I__590\ : ClkMux
    port map (
            O => \N__3643\,
            I => \N__3568\
        );

    \I__589\ : ClkMux
    port map (
            O => \N__3642\,
            I => \N__3568\
        );

    \I__588\ : ClkMux
    port map (
            O => \N__3641\,
            I => \N__3568\
        );

    \I__587\ : ClkMux
    port map (
            O => \N__3640\,
            I => \N__3568\
        );

    \I__586\ : ClkMux
    port map (
            O => \N__3639\,
            I => \N__3568\
        );

    \I__585\ : ClkMux
    port map (
            O => \N__3638\,
            I => \N__3568\
        );

    \I__584\ : ClkMux
    port map (
            O => \N__3637\,
            I => \N__3568\
        );

    \I__583\ : ClkMux
    port map (
            O => \N__3636\,
            I => \N__3568\
        );

    \I__582\ : ClkMux
    port map (
            O => \N__3635\,
            I => \N__3568\
        );

    \I__581\ : ClkMux
    port map (
            O => \N__3634\,
            I => \N__3568\
        );

    \I__580\ : ClkMux
    port map (
            O => \N__3633\,
            I => \N__3568\
        );

    \I__579\ : ClkMux
    port map (
            O => \N__3632\,
            I => \N__3568\
        );

    \I__578\ : ClkMux
    port map (
            O => \N__3631\,
            I => \N__3568\
        );

    \I__577\ : ClkMux
    port map (
            O => \N__3630\,
            I => \N__3568\
        );

    \I__576\ : ClkMux
    port map (
            O => \N__3629\,
            I => \N__3568\
        );

    \I__575\ : ClkMux
    port map (
            O => \N__3628\,
            I => \N__3568\
        );

    \I__574\ : ClkMux
    port map (
            O => \N__3627\,
            I => \N__3568\
        );

    \I__573\ : ClkMux
    port map (
            O => \N__3626\,
            I => \N__3568\
        );

    \I__572\ : ClkMux
    port map (
            O => \N__3625\,
            I => \N__3568\
        );

    \I__571\ : ClkMux
    port map (
            O => \N__3624\,
            I => \N__3568\
        );

    \I__570\ : ClkMux
    port map (
            O => \N__3623\,
            I => \N__3568\
        );

    \I__569\ : GlobalMux
    port map (
            O => \N__3568\,
            I => \N__3565\
        );

    \I__568\ : gio2CtrlBuf
    port map (
            O => \N__3565\,
            I => \CLK40_c_g\
        );

    \I__567\ : CEMux
    port map (
            O => \N__3562\,
            I => \N__3559\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3559\,
            I => \N__3556\
        );

    \I__565\ : Odrv12
    port map (
            O => \N__3556\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__3553\,
            I => \U400_SDRAM.N_252_cascade_\
        );

    \I__563\ : CascadeMux
    port map (
            O => \N__3550\,
            I => \N__3547\
        );

    \I__562\ : InMux
    port map (
            O => \N__3547\,
            I => \N__3543\
        );

    \I__561\ : InMux
    port map (
            O => \N__3546\,
            I => \N__3540\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3543\,
            I => \U400_SDRAM.RAM_CYCLEZ0\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3540\,
            I => \U400_SDRAM.RAM_CYCLEZ0\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__3535\,
            I => \U400_SDRAM.N_75_cascade_\
        );

    \I__557\ : InMux
    port map (
            O => \N__3532\,
            I => \N__3529\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3529\,
            I => \U400_SDRAM.CS1_EN_0\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__3526\,
            I => \U400_SDRAM.CS1_EN_7_i_0_o3_0_cascade_\
        );

    \I__554\ : InMux
    port map (
            O => \N__3523\,
            I => \N__3520\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3520\,
            I => \U400_SDRAM.N_159\
        );

    \I__552\ : InMux
    port map (
            O => \N__3517\,
            I => \N__3511\
        );

    \I__551\ : InMux
    port map (
            O => \N__3516\,
            I => \N__3511\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3511\,
            I => \N__3508\
        );

    \I__549\ : Odrv12
    port map (
            O => \N__3508\,
            I => \A_c_23\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__3505\,
            I => \N__3502\
        );

    \I__547\ : InMux
    port map (
            O => \N__3502\,
            I => \N__3498\
        );

    \I__546\ : InMux
    port map (
            O => \N__3501\,
            I => \N__3495\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3498\,
            I => \U400_SDRAM.CS0_ENZ0\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3495\,
            I => \U400_SDRAM.CS0_ENZ0\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__3490\,
            I => \U400_SDRAM.N_159_cascade_\
        );

    \I__542\ : InMux
    port map (
            O => \N__3487\,
            I => \N__3484\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3484\,
            I => \U400_SDRAM.N_75\
        );

    \I__540\ : InMux
    port map (
            O => \N__3481\,
            I => \N__3478\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3478\,
            I => \U400_SDRAM.CS0_EN_0\
        );

    \I__538\ : InMux
    port map (
            O => \N__3475\,
            I => \N__3472\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3472\,
            I => \N__3468\
        );

    \I__536\ : InMux
    port map (
            O => \N__3471\,
            I => \N__3465\
        );

    \I__535\ : Odrv12
    port map (
            O => \N__3468\,
            I => \U400_SDRAM.N_250\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3465\,
            I => \U400_SDRAM.N_250\
        );

    \I__533\ : InMux
    port map (
            O => \N__3460\,
            I => \N__3457\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3457\,
            I => \U400_SDRAM.N_189\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__3454\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_1_32_i_0_i_1_1_cascade_\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__3451\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_1_32_i_0_i_1_cascade_\
        );

    \I__529\ : CascadeMux
    port map (
            O => \N__3448\,
            I => \N__3445\
        );

    \I__528\ : InMux
    port map (
            O => \N__3445\,
            I => \N__3440\
        );

    \I__527\ : InMux
    port map (
            O => \N__3444\,
            I => \N__3435\
        );

    \I__526\ : InMux
    port map (
            O => \N__3443\,
            I => \N__3435\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3440\,
            I => \U400_SDRAM.N_128\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3435\,
            I => \U400_SDRAM.N_128\
        );

    \I__523\ : InMux
    port map (
            O => \N__3430\,
            I => \N__3427\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3427\,
            I => \U400_SDRAM.N_185\
        );

    \I__521\ : SRMux
    port map (
            O => \N__3424\,
            I => \N__3420\
        );

    \I__520\ : SRMux
    port map (
            O => \N__3423\,
            I => \N__3417\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3420\,
            I => \N__3412\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3417\,
            I => \N__3412\
        );

    \I__517\ : Odrv4
    port map (
            O => \N__3412\,
            I => \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1\
        );

    \I__516\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3405\
        );

    \I__515\ : InMux
    port map (
            O => \N__3408\,
            I => \N__3402\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__3405\,
            I => \N__3399\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3402\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__512\ : Odrv4
    port map (
            O => \N__3399\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__511\ : InMux
    port map (
            O => \N__3394\,
            I => \N__3390\
        );

    \I__510\ : InMux
    port map (
            O => \N__3393\,
            I => \N__3387\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3390\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3387\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__507\ : CascadeMux
    port map (
            O => \N__3382\,
            I => \N__3378\
        );

    \I__506\ : InMux
    port map (
            O => \N__3381\,
            I => \N__3375\
        );

    \I__505\ : InMux
    port map (
            O => \N__3378\,
            I => \N__3372\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3375\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3372\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__502\ : InMux
    port map (
            O => \N__3367\,
            I => \N__3362\
        );

    \I__501\ : InMux
    port map (
            O => \N__3366\,
            I => \N__3359\
        );

    \I__500\ : InMux
    port map (
            O => \N__3365\,
            I => \N__3356\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3362\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3359\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3356\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__496\ : InMux
    port map (
            O => \N__3349\,
            I => \N__3346\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3346\,
            I => \N__3336\
        );

    \I__494\ : InMux
    port map (
            O => \N__3345\,
            I => \N__3331\
        );

    \I__493\ : InMux
    port map (
            O => \N__3344\,
            I => \N__3331\
        );

    \I__492\ : InMux
    port map (
            O => \N__3343\,
            I => \N__3328\
        );

    \I__491\ : InMux
    port map (
            O => \N__3342\,
            I => \N__3319\
        );

    \I__490\ : InMux
    port map (
            O => \N__3341\,
            I => \N__3319\
        );

    \I__489\ : InMux
    port map (
            O => \N__3340\,
            I => \N__3319\
        );

    \I__488\ : InMux
    port map (
            O => \N__3339\,
            I => \N__3319\
        );

    \I__487\ : Odrv4
    port map (
            O => \N__3336\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_0\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3331\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_0\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3328\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_0\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3319\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_0\
        );

    \I__483\ : InMux
    port map (
            O => \N__3310\,
            I => \N__3305\
        );

    \I__482\ : InMux
    port map (
            O => \N__3309\,
            I => \N__3300\
        );

    \I__481\ : InMux
    port map (
            O => \N__3308\,
            I => \N__3300\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3305\,
            I => \U400_SDRAM.BURSTZ0\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3300\,
            I => \U400_SDRAM.BURSTZ0\
        );

    \I__478\ : InMux
    port map (
            O => \N__3295\,
            I => \N__3292\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3292\,
            I => \U400_SDRAM.TA_EN11_m\
        );

    \I__476\ : InMux
    port map (
            O => \N__3289\,
            I => \N__3285\
        );

    \I__475\ : InMux
    port map (
            O => \N__3288\,
            I => \N__3282\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3285\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3282\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__472\ : CascadeMux
    port map (
            O => \N__3277\,
            I => \N__3272\
        );

    \I__471\ : InMux
    port map (
            O => \N__3276\,
            I => \N__3266\
        );

    \I__470\ : InMux
    port map (
            O => \N__3275\,
            I => \N__3266\
        );

    \I__469\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3263\
        );

    \I__468\ : InMux
    port map (
            O => \N__3271\,
            I => \N__3260\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__3266\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3263\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3260\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__464\ : CascadeMux
    port map (
            O => \N__3253\,
            I => \N__3249\
        );

    \I__463\ : InMux
    port map (
            O => \N__3252\,
            I => \N__3246\
        );

    \I__462\ : InMux
    port map (
            O => \N__3249\,
            I => \N__3243\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__3246\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__3243\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__459\ : InMux
    port map (
            O => \N__3238\,
            I => \N__3234\
        );

    \I__458\ : InMux
    port map (
            O => \N__3237\,
            I => \N__3231\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3234\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__3231\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__455\ : CascadeMux
    port map (
            O => \N__3226\,
            I => \U400_SDRAM.N_205_cascade_\
        );

    \I__454\ : CascadeMux
    port map (
            O => \N__3223\,
            I => \N__3220\
        );

    \I__453\ : InMux
    port map (
            O => \N__3220\,
            I => \N__3217\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3217\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en\
        );

    \I__451\ : InMux
    port map (
            O => \N__3214\,
            I => \N__3211\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3211\,
            I => \U400_SDRAM.un1_REFRESH_COUNTERlto7_4\
        );

    \I__449\ : InMux
    port map (
            O => \N__3208\,
            I => \N__3204\
        );

    \I__448\ : InMux
    port map (
            O => \N__3207\,
            I => \N__3201\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3204\,
            I => \N__3198\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__3201\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\
        );

    \I__445\ : Odrv4
    port map (
            O => \N__3198\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\
        );

    \I__444\ : InMux
    port map (
            O => \N__3193\,
            I => \N__3190\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__3190\,
            I => \U400_SDRAM.un1_REFRESH_COUNTERlto7_5\
        );

    \I__442\ : InMux
    port map (
            O => \N__3187\,
            I => \N__3183\
        );

    \I__441\ : InMux
    port map (
            O => \N__3186\,
            I => \N__3180\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3183\,
            I => \U400_SDRAM.N_255\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3180\,
            I => \U400_SDRAM.N_255\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__3175\,
            I => \U400_SDRAM.TACK_7_iv_i_i_0_cascade_\
        );

    \I__437\ : InMux
    port map (
            O => \N__3172\,
            I => \N__3169\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3169\,
            I => \U400_SDRAM.TACK_7_iv_i_i_1\
        );

    \I__435\ : InMux
    port map (
            O => \N__3166\,
            I => \N__3163\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3163\,
            I => \U400_SDRAM.N_15\
        );

    \I__433\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3157\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__3157\,
            I => \U400_SDRAM.RAM_CYCLE_e_1\
        );

    \I__431\ : InMux
    port map (
            O => \N__3154\,
            I => \N__3149\
        );

    \I__430\ : InMux
    port map (
            O => \N__3153\,
            I => \N__3144\
        );

    \I__429\ : InMux
    port map (
            O => \N__3152\,
            I => \N__3144\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3149\,
            I => \U400_SDRAM.N_6\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3144\,
            I => \U400_SDRAM.N_6\
        );

    \I__426\ : InMux
    port map (
            O => \N__3139\,
            I => \N__3136\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3136\,
            I => \N__3133\
        );

    \I__424\ : Span4Mux_v
    port map (
            O => \N__3133\,
            I => \N__3130\
        );

    \I__423\ : Span4Mux_h
    port map (
            O => \N__3130\,
            I => \N__3127\
        );

    \I__422\ : Odrv4
    port map (
            O => \N__3127\,
            I => \RnW_c\
        );

    \I__421\ : IoInMux
    port map (
            O => \N__3124\,
            I => \N__3121\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3121\,
            I => \N__3118\
        );

    \I__419\ : IoSpan4Mux
    port map (
            O => \N__3118\,
            I => \N__3115\
        );

    \I__418\ : Span4Mux_s3_h
    port map (
            O => \N__3115\,
            I => \N__3112\
        );

    \I__417\ : Odrv4
    port map (
            O => \N__3112\,
            I => \CS0n_c\
        );

    \I__416\ : CascadeMux
    port map (
            O => \N__3109\,
            I => \N__3106\
        );

    \I__415\ : InMux
    port map (
            O => \N__3106\,
            I => \N__3103\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__3103\,
            I => \N__3100\
        );

    \I__413\ : Span4Mux_v
    port map (
            O => \N__3100\,
            I => \N__3097\
        );

    \I__412\ : Sp12to4
    port map (
            O => \N__3097\,
            I => \N__3094\
        );

    \I__411\ : Odrv12
    port map (
            O => \N__3094\,
            I => \A_c_19\
        );

    \I__410\ : IoInMux
    port map (
            O => \N__3091\,
            I => \N__3088\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3088\,
            I => \N__3085\
        );

    \I__408\ : Odrv12
    port map (
            O => \N__3085\,
            I => \MA_c_9\
        );

    \I__407\ : InMux
    port map (
            O => \N__3082\,
            I => \N__3074\
        );

    \I__406\ : InMux
    port map (
            O => \N__3081\,
            I => \N__3071\
        );

    \I__405\ : InMux
    port map (
            O => \N__3080\,
            I => \N__3062\
        );

    \I__404\ : InMux
    port map (
            O => \N__3079\,
            I => \N__3062\
        );

    \I__403\ : InMux
    port map (
            O => \N__3078\,
            I => \N__3062\
        );

    \I__402\ : InMux
    port map (
            O => \N__3077\,
            I => \N__3062\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__3074\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_1\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3071\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_1\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3062\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_1\
        );

    \I__398\ : CascadeMux
    port map (
            O => \N__3055\,
            I => \N__3050\
        );

    \I__397\ : CascadeMux
    port map (
            O => \N__3054\,
            I => \N__3045\
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__3053\,
            I => \N__3042\
        );

    \I__395\ : InMux
    port map (
            O => \N__3050\,
            I => \N__3039\
        );

    \I__394\ : InMux
    port map (
            O => \N__3049\,
            I => \N__3032\
        );

    \I__393\ : InMux
    port map (
            O => \N__3048\,
            I => \N__3032\
        );

    \I__392\ : InMux
    port map (
            O => \N__3045\,
            I => \N__3032\
        );

    \I__391\ : InMux
    port map (
            O => \N__3042\,
            I => \N__3029\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3039\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_3\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__3032\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_3\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3029\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_3\
        );

    \I__387\ : InMux
    port map (
            O => \N__3022\,
            I => \N__3018\
        );

    \I__386\ : InMux
    port map (
            O => \N__3021\,
            I => \N__3015\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__3018\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3015\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa\
        );

    \I__383\ : InMux
    port map (
            O => \N__3010\,
            I => \N__3006\
        );

    \I__382\ : InMux
    port map (
            O => \N__3009\,
            I => \N__3003\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__3006\,
            I => \U400_SDRAM.TA_COUNTER27\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__3003\,
            I => \U400_SDRAM.TA_COUNTER27\
        );

    \I__379\ : CascadeMux
    port map (
            O => \N__2998\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__2995\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER52_2_0_i_1_cascade_\
        );

    \I__377\ : InMux
    port map (
            O => \N__2992\,
            I => \N__2986\
        );

    \I__376\ : InMux
    port map (
            O => \N__2991\,
            I => \N__2986\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2986\,
            I => \U400_SDRAM.N_23\
        );

    \I__374\ : InMux
    port map (
            O => \N__2983\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_1\
        );

    \I__373\ : InMux
    port map (
            O => \N__2980\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_2\
        );

    \I__372\ : InMux
    port map (
            O => \N__2977\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_3\
        );

    \I__371\ : InMux
    port map (
            O => \N__2974\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_4\
        );

    \I__370\ : InMux
    port map (
            O => \N__2971\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_5\
        );

    \I__369\ : InMux
    port map (
            O => \N__2968\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_6\
        );

    \I__368\ : InMux
    port map (
            O => \N__2965\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_7\
        );

    \I__367\ : CascadeMux
    port map (
            O => \N__2962\,
            I => \N__2955\
        );

    \I__366\ : InMux
    port map (
            O => \N__2961\,
            I => \N__2951\
        );

    \I__365\ : InMux
    port map (
            O => \N__2960\,
            I => \N__2948\
        );

    \I__364\ : InMux
    port map (
            O => \N__2959\,
            I => \N__2939\
        );

    \I__363\ : InMux
    port map (
            O => \N__2958\,
            I => \N__2939\
        );

    \I__362\ : InMux
    port map (
            O => \N__2955\,
            I => \N__2939\
        );

    \I__361\ : InMux
    port map (
            O => \N__2954\,
            I => \N__2939\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2951\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_2\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2948\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_2\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2939\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_2\
        );

    \I__357\ : InMux
    port map (
            O => \N__2932\,
            I => \N__2929\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2929\,
            I => \U400_SDRAM.un1_TA_COUNTER26_2_0\
        );

    \I__355\ : IoInMux
    port map (
            O => \N__2926\,
            I => \N__2923\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2923\,
            I => \N__2919\
        );

    \I__353\ : CascadeMux
    port map (
            O => \N__2922\,
            I => \N__2916\
        );

    \I__352\ : Span12Mux_s7_h
    port map (
            O => \N__2919\,
            I => \N__2913\
        );

    \I__351\ : InMux
    port map (
            O => \N__2916\,
            I => \N__2910\
        );

    \I__350\ : Odrv12
    port map (
            O => \N__2913\,
            I => \TA_OUT\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2910\,
            I => \TA_OUT\
        );

    \I__348\ : CascadeMux
    port map (
            O => \N__2905\,
            I => \U400_SDRAM.N_208_cascade_\
        );

    \I__347\ : CascadeMux
    port map (
            O => \N__2902\,
            I => \N__2899\
        );

    \I__346\ : InMux
    port map (
            O => \N__2899\,
            I => \N__2896\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__2896\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_2\
        );

    \I__344\ : IoInMux
    port map (
            O => \N__2893\,
            I => \N__2890\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2890\,
            I => \N__2887\
        );

    \I__342\ : Span4Mux_s3_h
    port map (
            O => \N__2887\,
            I => \N__2884\
        );

    \I__341\ : Odrv4
    port map (
            O => \N__2884\,
            I => \RASn_c\
        );

    \I__340\ : IoInMux
    port map (
            O => \N__2881\,
            I => \N__2878\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__2878\,
            I => \N__2875\
        );

    \I__338\ : Odrv12
    port map (
            O => \N__2875\,
            I => \CASn_c\
        );

    \I__337\ : IoInMux
    port map (
            O => \N__2872\,
            I => \N__2869\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2869\,
            I => \N__2866\
        );

    \I__335\ : Odrv12
    port map (
            O => \N__2866\,
            I => \WEn_c\
        );

    \I__334\ : InMux
    port map (
            O => \N__2863\,
            I => \N__2860\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2860\,
            I => \N__2857\
        );

    \I__332\ : Span4Mux_h
    port map (
            O => \N__2857\,
            I => \N__2854\
        );

    \I__331\ : Sp12to4
    port map (
            O => \N__2854\,
            I => \N__2851\
        );

    \I__330\ : Span12Mux_v
    port map (
            O => \N__2851\,
            I => \N__2848\
        );

    \I__329\ : Odrv12
    port map (
            O => \N__2848\,
            I => \A_c_24\
        );

    \I__328\ : CascadeMux
    port map (
            O => \N__2845\,
            I => \N__2842\
        );

    \I__327\ : InMux
    port map (
            O => \N__2842\,
            I => \N__2839\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2839\,
            I => \N__2836\
        );

    \I__325\ : Span12Mux_s10_v
    port map (
            O => \N__2836\,
            I => \N__2833\
        );

    \I__324\ : Odrv12
    port map (
            O => \N__2833\,
            I => \A_c_18\
        );

    \I__323\ : IoInMux
    port map (
            O => \N__2830\,
            I => \N__2827\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__2827\,
            I => \N__2824\
        );

    \I__321\ : Span4Mux_s1_v
    port map (
            O => \N__2824\,
            I => \N__2821\
        );

    \I__320\ : Odrv4
    port map (
            O => \N__2821\,
            I => \MA_c_8\
        );

    \I__319\ : InMux
    port map (
            O => \N__2818\,
            I => \N__2815\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2815\,
            I => \N__2812\
        );

    \I__317\ : Span4Mux_v
    port map (
            O => \N__2812\,
            I => \N__2809\
        );

    \I__316\ : Odrv4
    port map (
            O => \N__2809\,
            I => \A_c_17\
        );

    \I__315\ : InMux
    port map (
            O => \N__2806\,
            I => \N__2803\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2803\,
            I => \N__2800\
        );

    \I__313\ : Odrv12
    port map (
            O => \N__2800\,
            I => \A_c_9\
        );

    \I__312\ : IoInMux
    port map (
            O => \N__2797\,
            I => \N__2794\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2794\,
            I => \N__2791\
        );

    \I__310\ : Odrv12
    port map (
            O => \N__2791\,
            I => \MA_c_7\
        );

    \I__309\ : InMux
    port map (
            O => \N__2788\,
            I => \N__2785\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2785\,
            I => \N__2782\
        );

    \I__307\ : Odrv12
    port map (
            O => \N__2782\,
            I => \A_c_8\
        );

    \I__306\ : CascadeMux
    port map (
            O => \N__2779\,
            I => \N__2776\
        );

    \I__305\ : InMux
    port map (
            O => \N__2776\,
            I => \N__2773\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2773\,
            I => \N__2770\
        );

    \I__303\ : Span4Mux_v
    port map (
            O => \N__2770\,
            I => \N__2767\
        );

    \I__302\ : Span4Mux_v
    port map (
            O => \N__2767\,
            I => \N__2764\
        );

    \I__301\ : Odrv4
    port map (
            O => \N__2764\,
            I => \A_c_16\
        );

    \I__300\ : IoInMux
    port map (
            O => \N__2761\,
            I => \N__2758\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2758\,
            I => \N__2755\
        );

    \I__298\ : Odrv12
    port map (
            O => \N__2755\,
            I => \MA_c_6\
        );

    \I__297\ : CascadeMux
    port map (
            O => \N__2752\,
            I => \U400_SDRAM.TA_COUNTER23_cascade_\
        );

    \I__296\ : InMux
    port map (
            O => \N__2749\,
            I => \N__2746\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2746\,
            I => \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0\
        );

    \I__294\ : CascadeMux
    port map (
            O => \N__2743\,
            I => \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_\
        );

    \I__293\ : InMux
    port map (
            O => \N__2740\,
            I => \N__2737\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2737\,
            I => \U400_SDRAM.CO1\
        );

    \I__291\ : CascadeMux
    port map (
            O => \N__2734\,
            I => \U400_SDRAM.CO1_cascade_\
        );

    \I__290\ : CascadeMux
    port map (
            O => \N__2731\,
            I => \N__2728\
        );

    \I__289\ : InMux
    port map (
            O => \N__2728\,
            I => \N__2725\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2725\,
            I => \N__2722\
        );

    \I__287\ : Span4Mux_v
    port map (
            O => \N__2722\,
            I => \N__2719\
        );

    \I__286\ : Odrv4
    port map (
            O => \N__2719\,
            I => \A_c_21\
        );

    \I__285\ : IoInMux
    port map (
            O => \N__2716\,
            I => \N__2713\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2713\,
            I => \N__2710\
        );

    \I__283\ : Span4Mux_s3_h
    port map (
            O => \N__2710\,
            I => \N__2707\
        );

    \I__282\ : Span4Mux_v
    port map (
            O => \N__2707\,
            I => \N__2703\
        );

    \I__281\ : InMux
    port map (
            O => \N__2706\,
            I => \N__2700\
        );

    \I__280\ : Odrv4
    port map (
            O => \N__2703\,
            I => \BANK0_c\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2700\,
            I => \BANK0_c\
        );

    \I__278\ : CascadeMux
    port map (
            O => \N__2695\,
            I => \N__2692\
        );

    \I__277\ : InMux
    port map (
            O => \N__2692\,
            I => \N__2689\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2689\,
            I => \N__2686\
        );

    \I__275\ : Span4Mux_h
    port map (
            O => \N__2686\,
            I => \N__2683\
        );

    \I__274\ : Span4Mux_v
    port map (
            O => \N__2683\,
            I => \N__2680\
        );

    \I__273\ : Odrv4
    port map (
            O => \N__2680\,
            I => \A_c_22\
        );

    \I__272\ : IoInMux
    port map (
            O => \N__2677\,
            I => \N__2674\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2674\,
            I => \N__2671\
        );

    \I__270\ : Span4Mux_s3_h
    port map (
            O => \N__2671\,
            I => \N__2668\
        );

    \I__269\ : Span4Mux_v
    port map (
            O => \N__2668\,
            I => \N__2664\
        );

    \I__268\ : InMux
    port map (
            O => \N__2667\,
            I => \N__2661\
        );

    \I__267\ : Odrv4
    port map (
            O => \N__2664\,
            I => \BANK1_c\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2661\,
            I => \BANK1_c\
        );

    \I__265\ : CascadeMux
    port map (
            O => \N__2656\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_a3_0_cascade_\
        );

    \I__264\ : InMux
    port map (
            O => \N__2653\,
            I => \N__2650\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__2650\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_1\
        );

    \I__262\ : IoInMux
    port map (
            O => \N__2647\,
            I => \N__2644\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2644\,
            I => \N__2641\
        );

    \I__260\ : Odrv4
    port map (
            O => \N__2641\,
            I => \RESETn_c_i\
        );

    \I__259\ : InMux
    port map (
            O => \N__2638\,
            I => \N__2635\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__2635\,
            I => \N__2632\
        );

    \I__257\ : Span4Mux_h
    port map (
            O => \N__2632\,
            I => \N__2629\
        );

    \I__256\ : Odrv4
    port map (
            O => \N__2629\,
            I => \A_c_30\
        );

    \I__255\ : InMux
    port map (
            O => \N__2626\,
            I => \N__2623\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2623\,
            I => \N__2620\
        );

    \I__253\ : Span12Mux_s10_h
    port map (
            O => \N__2620\,
            I => \N__2617\
        );

    \I__252\ : Odrv12
    port map (
            O => \N__2617\,
            I => \A_c_29\
        );

    \I__251\ : CascadeMux
    port map (
            O => \N__2614\,
            I => \N__2611\
        );

    \I__250\ : InMux
    port map (
            O => \N__2611\,
            I => \N__2608\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__2608\,
            I => \A_c_28\
        );

    \I__248\ : InMux
    port map (
            O => \N__2605\,
            I => \N__2602\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__2602\,
            I => \N__2599\
        );

    \I__246\ : Span4Mux_s1_v
    port map (
            O => \N__2599\,
            I => \N__2596\
        );

    \I__245\ : Odrv4
    port map (
            O => \N__2596\,
            I => \A_c_27\
        );

    \I__244\ : CascadeMux
    port map (
            O => \N__2593\,
            I => \U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_\
        );

    \I__243\ : CascadeMux
    port map (
            O => \N__2590\,
            I => \U400_SDRAM.un1_TA_COUNTER26_0_cascade_\
        );

    \I__242\ : IoInMux
    port map (
            O => \N__2587\,
            I => \N__2584\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__2584\,
            I => \N__2581\
        );

    \I__240\ : IoSpan4Mux
    port map (
            O => \N__2581\,
            I => \N__2578\
        );

    \I__239\ : IoSpan4Mux
    port map (
            O => \N__2578\,
            I => \N__2575\
        );

    \I__238\ : Span4Mux_s2_h
    port map (
            O => \N__2575\,
            I => \N__2572\
        );

    \I__237\ : Sp12to4
    port map (
            O => \N__2572\,
            I => \N__2569\
        );

    \I__236\ : Odrv12
    port map (
            O => \N__2569\,
            I => \CLK40_ibuf_gb_io_gb_input\
        );

    \INVU400_SDRAM.MA_2C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_2C_net\,
            I => \N__3649\
        );

    \INVU400_SDRAM.MA_3C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_3C_net\,
            I => \N__3646\
        );

    \INVU400_SDRAM.MA_0C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_0C_net\,
            I => \N__3648\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_2C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            I => \N__3638\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_1C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_1C_net\,
            I => \N__3642\
        );

    \INVU400_SDRAM.MA_4C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_4C_net\,
            I => \N__3647\
        );

    \INVU400_SDRAM.MA_11C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_11C_net\,
            I => \N__3632\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_0C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_0C_net\,
            I => \N__3625\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_3C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_3C_net\,
            I => \N__3637\
        );

    \INVU400_SDRAM.SDRAM_CMD_2C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CMD_2C_net\,
            I => \N__3641\
        );

    \INVU400_SDRAM.CS1nC\ : INV
    port map (
            O => \INVU400_SDRAM.CS1nC_net\,
            I => \N__3629\
        );

    \INVU400_SDRAM.SDRAM_CMD_0C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CMD_0C_net\,
            I => \N__3636\
        );

    \INVU400_SDRAM.SDRAM_CMD_1C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CMD_1C_net\,
            I => \N__3640\
        );

    \INVU400_SDRAM.REFRESH_COUNTER_0C\ : INV
    port map (
            O => \INVU400_SDRAM.REFRESH_COUNTER_0C_net\,
            I => \N__3645\
        );

    \INVU400_SDRAM.CS0_ENC\ : INV
    port map (
            O => \INVU400_SDRAM.CS0_ENC_net\,
            I => \N__3624\
        );

    \INVU400_SDRAM.RAM_CYCLEC\ : INV
    port map (
            O => \INVU400_SDRAM.RAM_CYCLEC_net\,
            I => \N__3628\
        );

    \INVU400_SDRAM.BURSTC\ : INV
    port map (
            O => \INVU400_SDRAM.BURSTC_net\,
            I => \N__3635\
        );

    \INVU400_SDRAM.REFRESH_COUNTER_2C\ : INV
    port map (
            O => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            I => \N__3643\
        );

    \INVU400_SDRAM.MA_6C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_6C_net\,
            I => \N__3633\
        );

    \INVU400_SDRAM.MA_8C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_8C_net\,
            I => \N__3626\
        );

    \INVU400_SDRAM.RASnC\ : INV
    port map (
            O => \INVU400_SDRAM.RASnC_net\,
            I => \N__3623\
        );

    \INVU400_SDRAM.BANK0C\ : INV
    port map (
            O => \INVU400_SDRAM.BANK0C_net\,
            I => \N__3627\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_3_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \CLK40_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2587\,
            GLOBALBUFFEROUTPUT => \CLK40_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2647\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5555\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.RAM_SPACE_0_a3_3_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__2638\,
            in1 => \N__2626\,
            in2 => \N__2614\,
            in3 => \N__2605\,
            lcout => \U400_ADDRESS_DECODE_RAM_SPACE_0_a3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__3345\,
            in1 => \N__3712\,
            in2 => \_gnd_net_\,
            in3 => \N__3686\,
            lcout => OPEN,
            ltout => \U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_0_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__5522\,
            in1 => \_gnd_net_\,
            in2 => \N__2593\,
            in3 => \N__3022\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3634\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_OUT_RNO_2_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__2960\,
            in1 => \N__3082\,
            in2 => \N__3055\,
            in3 => \N__3344\,
            lcout => OPEN,
            ltout => \U400_SDRAM.un1_TA_COUNTER26_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_OUT_RNO_1_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3713\,
            in2 => \N__2590\,
            in3 => \N__3687\,
            lcout => \U400_SDRAM.un1_TA_COUNTER26_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__3339\,
            in1 => \N__2954\,
            in2 => \N__3054\,
            in3 => \N__3077\,
            lcout => \U400_SDRAM.TA_COUNTER27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_1_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__3342\,
            in1 => \N__3080\,
            in2 => \N__5557\,
            in3 => \N__2749\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3630\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3078\,
            in1 => \N__3048\,
            in2 => \N__2962\,
            in3 => \N__3340\,
            lcout => \U400_SDRAM.TA_COUNTER23\,
            ltout => \U400_SDRAM.TA_COUNTER23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNI0LUG4_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__3010\,
            in1 => \N__3681\,
            in2 => \N__2752\,
            in3 => \N__3021\,
            lcout => \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0\,
            ltout => \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_2_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__2958\,
            in1 => \N__5551\,
            in2 => \N__2743\,
            in3 => \N__2740\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3630\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3341\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3079\,
            lcout => \U400_SDRAM.CO1\,
            ltout => \U400_SDRAM.CO1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_3_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110010000000"
        )
    port map (
            in0 => \N__2959\,
            in1 => \N__5552\,
            in2 => \N__2734\,
            in3 => \N__3049\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3630\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.BANK0_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__2991\,
            in1 => \N__2706\,
            in2 => \N__2731\,
            in3 => \N__3967\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK0C_net\,
            ce => 'H',
            sr => \N__5922\
        );

    \U400_SDRAM.BANK1_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__3966\,
            in1 => \N__2667\,
            in2 => \N__2695\,
            in3 => \N__2992\,
            lcout => \BANK1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK0C_net\,
            ce => 'H',
            sr => \N__5922\
        );

    \U400_SDRAM.TACK_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100000001"
        )
    port map (
            in0 => \N__3166\,
            in1 => \N__2653\,
            in2 => \N__2902\,
            in3 => \N__3685\,
            lcout => \U400_SDRAM.TACKZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK0C_net\,
            ce => 'H',
            sr => \N__5922\
        );

    \U400_SDRAM.TACK_RNO_6_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__5079\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4959\,
            lcout => OPEN,
            ltout => \U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_1_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100000"
        )
    port map (
            in0 => \N__5149\,
            in1 => \N__5269\,
            in2 => \N__2656\,
            in3 => \N__4741\,
            lcout => \U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_7_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__4960\,
            in1 => \N__5078\,
            in2 => \N__5159\,
            in3 => \N__4827\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_208_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_2_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111111"
        )
    port map (
            in0 => \N__5080\,
            in1 => \N__3187\,
            in2 => \N__2905\,
            in3 => \N__4712\,
            lcout => \U400_SDRAM.un1_SDRAM_COUNTER52_4_0_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RASn_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6049\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.RASnC_net\,
            ce => 'H',
            sr => \N__5921\
        );

    \U400_SDRAM.CASn_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6299\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.RASnC_net\,
            ce => 'H',
            sr => \N__5921\
        );

    \U400_SDRAM.WEn_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6198\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.RASnC_net\,
            ce => 'H',
            sr => \N__5921\
        );

    \U400_SDRAM.MA_8_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__2863\,
            in1 => \N__6113\,
            in2 => \N__2845\,
            in3 => \N__6360\,
            lcout => \MA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_8C_net\,
            ce => 'H',
            sr => \N__5924\
        );

    \U400_SDRAM.MA_7_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__2818\,
            in1 => \N__2806\,
            in2 => \N__6115\,
            in3 => \N__6359\,
            lcout => \MA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_8C_net\,
            ce => 'H',
            sr => \N__5924\
        );

    \U400_SDRAM.MA_6_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__2788\,
            in1 => \N__6109\,
            in2 => \N__2779\,
            in3 => \N__6376\,
            lcout => \MA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_6C_net\,
            ce => 'H',
            sr => \N__5932\
        );

    \U400_SDRAM.un2_REFRESH_COUNTER_cry_1_c_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3366\,
            in2 => \N__3277\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_2_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3394\,
            in2 => \_gnd_net_\,
            in3 => \N__2983\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un2_REFRESH_COUNTER_cry_1\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_2\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3424\
        );

    \U400_SDRAM.REFRESH_COUNTER_3_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3408\,
            in2 => \_gnd_net_\,
            in3 => \N__2980\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un2_REFRESH_COUNTER_cry_2\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_3\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3424\
        );

    \U400_SDRAM.REFRESH_COUNTER_4_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3381\,
            in2 => \_gnd_net_\,
            in3 => \N__2977\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un2_REFRESH_COUNTER_cry_3\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_4\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3424\
        );

    \U400_SDRAM.REFRESH_COUNTER_5_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3238\,
            in2 => \_gnd_net_\,
            in3 => \N__2974\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un2_REFRESH_COUNTER_cry_4\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_5\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3424\
        );

    \U400_SDRAM.REFRESH_COUNTER_6_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3289\,
            in2 => \_gnd_net_\,
            in3 => \N__2971\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un2_REFRESH_COUNTER_cry_5\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_6\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3424\
        );

    \U400_SDRAM.REFRESH_COUNTER_7_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3252\,
            in2 => \_gnd_net_\,
            in3 => \N__2968\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un2_REFRESH_COUNTER_cry_6\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_7\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3424\
        );

    \U400_SDRAM.REFRESH_COUNTER_8_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3207\,
            in2 => \_gnd_net_\,
            in3 => \N__2965\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3424\
        );

    \U400_SDRAM.TA_OUT_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__2961\,
            in1 => \N__2932\,
            in2 => \N__2922\,
            in3 => \N__3295\,
            lcout => \TA_OUT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3639\,
            ce => 'H',
            sr => \N__5927\
        );

    \U400_SDRAM.BURST_RNISKH51_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__3081\,
            in1 => \N__3343\,
            in2 => \N__3053\,
            in3 => \N__3308\,
            lcout => \U400_SDRAM.TA_COUNTER_0_sqmuxa\,
            ltout => \U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__3714\,
            in1 => \N__3009\,
            in2 => \N__2998\,
            in3 => \N__3675\,
            lcout => \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.BURST_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__3309\,
            in1 => \N__5751\,
            in2 => \N__5686\,
            in3 => \N__3154\,
            lcout => \U400_SDRAM.BURSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BURSTC_net\,
            ce => 'H',
            sr => \N__5925\
        );

    \U400_SDRAM.RAM_CYCLE_RNO_1_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111001111"
        )
    port map (
            in0 => \N__4963\,
            in1 => \N__5272\,
            in2 => \N__4709\,
            in3 => \N__5077\,
            lcout => OPEN,
            ltout => \U400_SDRAM.un1_SDRAM_COUNTER52_2_0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_RNO_0_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001100"
        )
    port map (
            in0 => \N__4015\,
            in1 => \N__3444\,
            in2 => \N__2995\,
            in3 => \N__3950\,
            lcout => \U400_SDRAM.RAM_CYCLE_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNISAQQ4_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4014\,
            in2 => \N__4711\,
            in3 => \N__4067\,
            lcout => \U400_SDRAM.N_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_5_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110001"
        )
    port map (
            in0 => \N__5271\,
            in1 => \N__3443\,
            in2 => \N__5152\,
            in3 => \N__4867\,
            lcout => \U400_SDRAM.TACK_7_iv_i_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNI58I35_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__3951\,
            in1 => \N__4066\,
            in2 => \N__4710\,
            in3 => \N__4013\,
            lcout => \U400_SDRAM.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.WRITE_CYCLE_RNI18LH_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__5270\,
            in1 => \N__5127\,
            in2 => \_gnd_net_\,
            in3 => \N__4961\,
            lcout => \U400_SDRAM.N_255\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_4_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011011100"
        )
    port map (
            in0 => \N__4962\,
            in1 => \N__4159\,
            in2 => \N__5150\,
            in3 => \N__5273\,
            lcout => OPEN,
            ltout => \U400_SDRAM.TACK_7_iv_i_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_0_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3186\,
            in1 => \N__3460\,
            in2 => \N__3175\,
            in3 => \N__3172\,
            lcout => \U400_SDRAM.N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001110010"
        )
    port map (
            in0 => \N__3160\,
            in1 => \N__3152\,
            in2 => \N__3550\,
            in3 => \N__4441\,
            lcout => \U400_SDRAM.RAM_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.RAM_CYCLEC_net\,
            ce => 'H',
            sr => \N__5923\
        );

    \U400_SDRAM.WRITE_CYCLE_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__3153\,
            in1 => \N__3139\,
            in2 => \_gnd_net_\,
            in3 => \N__5142\,
            lcout => \U400_SDRAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.RAM_CYCLEC_net\,
            ce => 'H',
            sr => \N__5923\
        );

    \U400_SDRAM.CS0_EN_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010011"
        )
    port map (
            in0 => \N__4029\,
            in1 => \N__4073\,
            in2 => \N__4713\,
            in3 => \N__3481\,
            lcout => \U400_SDRAM.CS0_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0_ENC_net\,
            ce => 'H',
            sr => \N__5920\
        );

    \U400_SDRAM.CS0n_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__6297\,
            in1 => \N__6055\,
            in2 => \N__3505\,
            in3 => \N__6188\,
            lcout => \CS0n_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0_ENC_net\,
            ce => 'H',
            sr => \N__5920\
        );

    \U400_SDRAM.MA_9_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6189\,
            in1 => \N__6056\,
            in2 => \N__3109\,
            in3 => \N__6298\,
            lcout => \MA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0_ENC_net\,
            ce => 'H',
            sr => \N__5920\
        );

    \U400_SDRAM.CS1_EN_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010101"
        )
    port map (
            in0 => \N__4074\,
            in1 => \N__4030\,
            in2 => \N__4714\,
            in3 => \N__3532\,
            lcout => \U400_SDRAM.CS1_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0_ENC_net\,
            ce => 'H',
            sr => \N__5920\
        );

    \U400_SDRAM.REFRESH_COUNTER_0_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3275\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__3423\
        );

    \U400_SDRAM.REFRESH_COUNTER_1_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3276\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3367\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__3423\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_1_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__5556\,
            in1 => \N__5276\,
            in2 => \_gnd_net_\,
            in3 => \N__3475\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNIMIPA1_1_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3409\,
            in1 => \N__3393\,
            in2 => \N__3382\,
            in3 => \N__3365\,
            lcout => \U400_SDRAM.un1_REFRESH_COUNTERlto7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_OUT_RNO_0_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3349\,
            in2 => \_gnd_net_\,
            in3 => \N__3310\,
            lcout => \U400_SDRAM.TA_EN11_m\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNIUQPA1_5_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3288\,
            in1 => \N__3271\,
            in2 => \N__3253\,
            in3 => \N__3237\,
            lcout => \U400_SDRAM.un1_REFRESH_COUNTERlto7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3846\,
            in1 => \N__4016\,
            in2 => \_gnd_net_\,
            in3 => \N__4825\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_205_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_1_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001011"
        )
    port map (
            in0 => \N__6255\,
            in1 => \N__3874\,
            in2 => \N__3226\,
            in3 => \N__3853\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__5941\,
            in1 => \_gnd_net_\,
            in2 => \N__3223\,
            in3 => \_gnd_net_\,
            lcout => \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNIVV903_8_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__3214\,
            in1 => \N__3208\,
            in2 => \_gnd_net_\,
            in3 => \N__3193\,
            lcout => \U400_SDRAM.REFRESH_COUNTER_RNIVV903Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__4012\,
            in1 => \N__4577\,
            in2 => \N__3448\,
            in3 => \N__3949\,
            lcout => \U400_SDRAM.N_199\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_3_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001100"
        )
    port map (
            in0 => \N__5274\,
            in1 => \N__5076\,
            in2 => \N__4828\,
            in3 => \N__5131\,
            lcout => \U400_SDRAM.N_189\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011101110111"
        )
    port map (
            in0 => \N__4824\,
            in1 => \N__3845\,
            in2 => \N__5151\,
            in3 => \N__4947\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_0_1_32_i_0_i_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__5275\,
            in1 => \N__4581\,
            in2 => \N__3454\,
            in3 => \N__5135\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_0_1_32_i_0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_0_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001011"
        )
    port map (
            in0 => \N__6161\,
            in1 => \N__3869\,
            in2 => \N__3451\,
            in3 => \N__3430\,
            lcout => \U400_SDRAM.SDRAM_CMDZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIP3PD_0_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__4939\,
            in1 => \_gnd_net_\,
            in2 => \N__5075\,
            in3 => \_gnd_net_\,
            lcout => \U400_SDRAM.N_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNITTDH4_0_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__5541\,
            in1 => \N__3820\,
            in2 => \_gnd_net_\,
            in3 => \N__4242\,
            lcout => \U400_SDRAM.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_0_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4938\,
            in1 => \N__5242\,
            in2 => \N__5074\,
            in3 => \N__4433\,
            lcout => \U400_SDRAM.N_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4147\,
            in2 => \_gnd_net_\,
            in3 => \N__4093\,
            lcout => \U400_SDRAM.N_185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__5764\,
            in1 => \N__3546\,
            in2 => \N__5554\,
            in3 => \N__3958\,
            lcout => \U400_SDRAM.RAM_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3631\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIPOT15_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101111111011"
        )
    port map (
            in0 => \N__4240\,
            in1 => \N__4065\,
            in2 => \N__4707\,
            in3 => \N__4092\,
            lcout => \U400_SDRAM.N_75\,
            ltout => \U400_SDRAM.N_75_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS1_EN_RNO_0_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001011100"
        )
    port map (
            in0 => \N__3517\,
            in1 => \N__3804\,
            in2 => \N__3535\,
            in3 => \N__3523\,
            lcout => \U400_SDRAM.CS1_EN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIHALH3_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__4091\,
            in1 => \N__4680\,
            in2 => \N__5281\,
            in3 => \N__4239\,
            lcout => OPEN,
            ltout => \U400_SDRAM.CS1_EN_7_i_0_o3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNIA1BE8_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__4019\,
            in1 => \N__3471\,
            in2 => \N__3526\,
            in3 => \N__3948\,
            lcout => \U400_SDRAM.N_159\,
            ltout => \U400_SDRAM.N_159_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS0_EN_RNO_0_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__3516\,
            in1 => \N__3501\,
            in2 => \N__3490\,
            in3 => \N__3487\,
            lcout => \U400_SDRAM.CS0_EN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIHPJJ1_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5039\,
            in1 => \N__4940\,
            in2 => \N__4706\,
            in3 => \N__4434\,
            lcout => \U400_SDRAM.N_250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__5043\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3744\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001000100010"
        )
    port map (
            in0 => \N__5280\,
            in1 => \N__5042\,
            in2 => \N__5160\,
            in3 => \N__4826\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_176_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__4640\,
            in1 => \N__4862\,
            in2 => \N__3814\,
            in3 => \N__4099\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS1n_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__6047\,
            in1 => \N__6190\,
            in2 => \N__3811\,
            in3 => \N__6301\,
            lcout => \CS1n_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS1nC_net\,
            ce => 'H',
            sr => \N__5926\
        );

    \U400_SDRAM.MA_12_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6048\,
            in1 => \N__6191\,
            in2 => \N__3784\,
            in3 => \N__6302\,
            lcout => \MA_c_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS1nC_net\,
            ce => 'H',
            sr => \N__5926\
        );

    \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101101010101"
        )
    port map (
            in0 => \N__6042\,
            in1 => \N__6162\,
            in2 => \_gnd_net_\,
            in3 => \N__6256\,
            lcout => \U400_SDRAM.MAc_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_UUBEn_0_a3_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011100000"
        )
    port map (
            in0 => \N__5841\,
            in1 => \N__5812\,
            in2 => \N__5752\,
            in3 => \N__5685\,
            lcout => \UUBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_EN_i_ess_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__5523\,
            in1 => \N__3718\,
            in2 => \_gnd_net_\,
            in3 => \N__3691\,
            lcout => \TA_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3644\,
            ce => \N__3562\,
            sr => \N__5933\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_0_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__5527\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4684\,
            lcout => \U400_SDRAM.N_252\,
            ltout => \U400_SDRAM.N_252_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__5241\,
            in1 => \N__4405\,
            in2 => \N__3553\,
            in3 => \N__4948\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_200_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__4132\,
            in1 => \N__3847\,
            in2 => \N__3889\,
            in3 => \N__4805\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_0_61_i_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_2_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000011"
        )
    port map (
            in0 => \N__6029\,
            in1 => \N__3886\,
            in2 => \N__3877\,
            in3 => \N__3873\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_2C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__4131\,
            in1 => \N__5240\,
            in2 => \N__4582\,
            in3 => \N__3826\,
            lcout => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIA54Q_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__5073\,
            in1 => \_gnd_net_\,
            in2 => \N__4708\,
            in3 => \N__5526\,
            lcout => \U400_SDRAM.N_228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__4565\,
            in1 => \N__3944\,
            in2 => \N__4075\,
            in3 => \N__4017\,
            lcout => \U400_SDRAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_0_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__4018\,
            in1 => \N__4069\,
            in2 => \N__3959\,
            in3 => \N__4566\,
            lcout => \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5Z0Z_0\,
            ltout => \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_3_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__5617\,
            in1 => \N__4372\,
            in2 => \N__3829\,
            in3 => \N__4314\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_3C_net\,
            ce => \N__5315\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__5236\,
            in1 => \N__4946\,
            in2 => \N__5553\,
            in3 => \N__4400\,
            lcout => \U400_SDRAM.N_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_0_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001110"
        )
    port map (
            in0 => \N__4734\,
            in1 => \N__5232\,
            in2 => \N__4576\,
            in3 => \N__5041\,
            lcout => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4332\,
            in1 => \N__4347\,
            in2 => \N__5335\,
            in3 => \N__4362\,
            lcout => \U400_SDRAM.N_126\,
            ltout => \U400_SDRAM.N_126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIFAF21_2_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4108\,
            in3 => \N__4778\,
            lcout => \U400_SDRAM.N_129\,
            ltout => \U400_SDRAM.N_129_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_0_0_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4927\,
            in1 => \N__5225\,
            in2 => \N__4105\,
            in3 => \N__5021\,
            lcout => \U400_SDRAM.N_257\,
            ltout => \U400_SDRAM.N_257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_5_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__5525\,
            in1 => \N__4660\,
            in2 => \N__4102\,
            in3 => \N__4928\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4926\,
            in1 => \N__5022\,
            in2 => \_gnd_net_\,
            in3 => \N__4431\,
            lcout => \U400_SDRAM.N_133\,
            ltout => \U400_SDRAM.N_133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4659\,
            in2 => \N__4078\,
            in3 => \N__4241\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_141_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIJG6G7_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__4068\,
            in1 => \N__5524\,
            in2 => \N__4033\,
            in3 => \N__4969\,
            lcout => \U400_SDRAM.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4028\,
            in1 => \N__4404\,
            in2 => \N__4723\,
            in3 => \N__3965\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_181_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_0_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__3904\,
            in1 => \N__3898\,
            in2 => \N__3892\,
            in3 => \N__4306\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_0C_net\,
            ce => \N__5319\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_11_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6046\,
            in1 => \N__6203\,
            in2 => \N__4273\,
            in3 => \N__6300\,
            lcout => \MA_c_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_11C_net\,
            ce => 'H',
            sr => \N__5928\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4641\,
            in2 => \_gnd_net_\,
            in3 => \N__4246\,
            lcout => \U400_SDRAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_11C_net\,
            ce => 'H',
            sr => \N__5928\
        );

    \U400_SDRAM.MA_4_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__4216\,
            in1 => \N__6090\,
            in2 => \N__4201\,
            in3 => \N__6384\,
            lcout => \MA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_4C_net\,
            ce => 'H',
            sr => \N__5935\
        );

    \U400_SDRAM.MA_5_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000110001"
        )
    port map (
            in0 => \N__6204\,
            in1 => \N__4501\,
            in2 => \N__6108\,
            in3 => \N__6318\,
            lcout => \MA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_4C_net\,
            ce => 'H',
            sr => \N__5935\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI6MLK_2_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__5072\,
            in1 => \N__4929\,
            in2 => \_gnd_net_\,
            in3 => \N__4803\,
            lcout => \U400_SDRAM.N_150\,
            ltout => \U400_SDRAM.N_150_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIVPE21_2_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__4804\,
            in1 => \_gnd_net_\,
            in2 => \N__4150\,
            in3 => \N__5268\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_0_61_i_i_a3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI079H2_2_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4146\,
            in2 => \N__4135\,
            in3 => \N__4866\,
            lcout => \U400_SDRAM.N_201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TAn_obuft_RNO_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4123\,
            lcout => \N_529_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_1_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__4384\,
            in1 => \N__4447\,
            in2 => \N__5613\,
            in3 => \N__4315\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_1C_net\,
            ce => \N__5314\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5040\,
            in2 => \_gnd_net_\,
            in3 => \N__4432\,
            lcout => \U400_SDRAM.N_260\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5267\,
            in2 => \_gnd_net_\,
            in3 => \N__4378\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_1\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_0\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_2_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4316\,
            in1 => \N__4802\,
            in2 => \_gnd_net_\,
            in3 => \N__4375\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_1\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_2\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__5320\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4949\,
            in2 => \_gnd_net_\,
            in3 => \N__4366\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_3\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_2\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_4_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4317\,
            in1 => \N__4363\,
            in2 => \_gnd_net_\,
            in3 => \N__4351\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_3\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_4\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__5320\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_5_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4304\,
            in1 => \N__4348\,
            in2 => \_gnd_net_\,
            in3 => \N__4336\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_4\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_5\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__5320\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_6_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4318\,
            in1 => \N__4333\,
            in2 => \_gnd_net_\,
            in3 => \N__4321\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_5\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_6\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__5320\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_7_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4305\,
            in1 => \N__5334\,
            in2 => \_gnd_net_\,
            in3 => \N__4276\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__5320\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011001100110"
        )
    port map (
            in0 => \N__4951\,
            in1 => \N__5266\,
            in2 => \N__5161\,
            in3 => \N__5038\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_161_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI4ECU1_2_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4780\,
            in1 => \N__4628\,
            in2 => \N__4972\,
            in3 => \N__4855\,
            lcout => \U400_SDRAM.N_183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNITTB91_2_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__4950\,
            in1 => \N__4854\,
            in2 => \_gnd_net_\,
            in3 => \N__4779\,
            lcout => \U400_SDRAM.N_138\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4629\,
            in1 => \N__5741\,
            in2 => \_gnd_net_\,
            in3 => \N__5675\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a3_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5488\,
            in2 => \_gnd_net_\,
            in3 => \N__4627\,
            lcout => \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_RNO_0_5_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000100"
        )
    port map (
            in0 => \N__4528\,
            in1 => \N__6087\,
            in2 => \N__4516\,
            in3 => \N__6303\,
            lcout => \U400_SDRAM.MAc_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_0_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__4495\,
            in1 => \N__6089\,
            in2 => \N__4483\,
            in3 => \N__6385\,
            lcout => \MA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_0C_net\,
            ce => 'H',
            sr => \N__5936\
        );

    \U400_SDRAM.MA_10_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000011010"
        )
    port map (
            in0 => \N__6088\,
            in1 => \N__6199\,
            in2 => \N__6319\,
            in3 => \N__4462\,
            lcout => \MA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_0C_net\,
            ce => 'H',
            sr => \N__5936\
        );

    \U400_BYTE_ENABLE.un1_UMBEn_0_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000001100100"
        )
    port map (
            in0 => \N__5744\,
            in1 => \N__5681\,
            in2 => \N__5857\,
            in3 => \N__5817\,
            lcout => \UMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_LLBEn_0_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100101010"
        )
    port map (
            in0 => \N__5679\,
            in1 => \N__5849\,
            in2 => \N__5818\,
            in3 => \N__5742\,
            lcout => \LLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_LMBEn_0_a3_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000110"
        )
    port map (
            in0 => \N__5743\,
            in1 => \N__5680\,
            in2 => \N__5856\,
            in3 => \N__5816\,
            lcout => \LMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5490\,
            in1 => \N__5596\,
            in2 => \N__5575\,
            in3 => \N__5776\,
            lcout => \U400_SDRAM.N_220\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.BURST8_0_a2_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5724\,
            in2 => \_gnd_net_\,
            in3 => \N__5664\,
            lcout => \U400_SDRAM.BURST8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.N_220_3_i_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__5595\,
            in1 => \N__5571\,
            in2 => \_gnd_net_\,
            in3 => \N__5489\,
            lcout => \N_220_3_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_3_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__5395\,
            in1 => \N__6078\,
            in2 => \N__5386\,
            in3 => \N__6375\,
            lcout => \MA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_3C_net\,
            ce => 'H',
            sr => \N__5934\
        );

    \U400_SDRAM.MA_RNO_0_1_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000100"
        )
    port map (
            in0 => \N__5359\,
            in1 => \N__6103\,
            in2 => \N__5347\,
            in3 => \N__6304\,
            lcout => \U400_SDRAM.MAc_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_2_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__6104\,
            in1 => \N__6409\,
            in2 => \N__6394\,
            in3 => \N__6383\,
            lcout => \MA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_2C_net\,
            ce => 'H',
            sr => \N__5937\
        );

    \U400_SDRAM.MA_1_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011001"
        )
    port map (
            in0 => \N__6314\,
            in1 => \N__6208\,
            in2 => \N__6114\,
            in3 => \N__5953\,
            lcout => \MA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_2C_net\,
            ce => 'H',
            sr => \N__5937\
        );
end \INTERFACE\;

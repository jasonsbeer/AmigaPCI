-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 15 2024 12:53:28

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RAMENn : out std_logic;
    RASn : out std_logic;
    TACKn : out std_logic;
    CLKEN : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__10331\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_OUT_i_i\ : std_logic;
signal \CLK40_OUT_i_i\ : std_logic;
signal \U712_REG_SM.N_120\ : std_logic;
signal \C3_c\ : std_logic;
signal \N_677_i\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \U712_REG_SM.N_86\ : std_logic;
signal \U712_REG_SM.N_68_cascade_\ : std_logic;
signal \U712_REG_SM.N_73_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \C1_c\ : std_logic;
signal \CLK40_OUT_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.N_45_0_0_en_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_45_0_0_en_0\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_REG_SM.N_73\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_5_0_1_cascade_\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_5\ : std_logic;
signal \U712_REG_SM.N_173_0_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.N_54_cascade_\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_5_0_1\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_REG_SM.N_162_0_cascade_\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_165_0_cascade_\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_6\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_a3_0\ : std_logic;
signal \U712_REG_SM.DS_EN_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_REG_SM.N_68\ : std_logic;
signal \U712_REG_SM.N_188_cascade_\ : std_logic;
signal \U712_REG_SM.N_162_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \ASn_c\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.DS_EN_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \U712_REG_SM.N_171_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U712_REG_SM.LDS_OUT_2_0_0\ : std_logic;
signal \U712_REG_SM.UDS_OUT_2_0_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.N_33\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.N_34\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_14\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_6_cascade_\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_167_0\ : std_logic;
signal \U712_REG_SM.N_117\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.RnW_m\ : std_logic;
signal \U712_REG_SM.un1_LDS_OUT_0_sqmuxa_1_0\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_0\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_1\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \U712_REG_SM.UDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_UDSn_i\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.N_32\ : std_logic;
signal \U712_CHIP_RAM.N_37\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_5\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.N_35\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.N_36_cascade_\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_ns_1_2\ : std_logic;
signal \U712_CHIP_RAM.N_61_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_65_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_104_1\ : std_logic;
signal \U712_CHIP_RAM.N_51\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER16_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_99_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_67_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER18_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_m2_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_7\ : std_logic;
signal \U712_BYTE_ENABLE.un2_CUMBEnZ0_cascade_\ : std_logic;
signal \CUMBEn_c\ : std_logic;
signal \U712_BYTE_ENABLE.LLBE_0_0_tz\ : std_logic;
signal \U712_BYTE_ENABLE.un2_CLLBEnZ0_cascade_\ : std_logic;
signal \CLLBEn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un2_CLMBEnZ0_cascade_\ : std_logic;
signal \CLMBEn_c\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \U712_BYTE_ENABLE.LW_TRANS_0\ : std_logic;
signal \U712_BYTE_ENABLE.un2_CUUBEnZ0_cascade_\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \CUUBEn_c\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \bfn_14_4_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8_cascade_\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.N_38\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER18_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_158_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_ns_1_1\ : std_logic;
signal \U712_CHIP_RAM.N_132\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_i\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER18_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0\ : std_logic;
signal \U712_REG_SM.DS_ENZ0\ : std_logic;
signal \U712_REG_SM.LDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_LDSn_i\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.N_39\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_1_a3_0\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6\ : std_logic;
signal \U712_REG_SM.N_173_0\ : std_logic;
signal \U712_REG_SM.N_183_1\ : std_logic;
signal \U712_REG_SM.N_165_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.un1_DBR_SYNC\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_2_1\ : std_logic;
signal \U712_CHIP_RAM.N_108\ : std_logic;
signal \U712_CHIP_RAM.N_77_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4\ : std_logic;
signal \U712_CHIP_RAM.N_80\ : std_logic;
signal \U712_CHIP_RAM.N_77\ : std_logic;
signal \U712_CHIP_RAM.N_80_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_50_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.N_60\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER39_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER39_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_50\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \DRDDIR_0_i\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i_0\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.N_65\ : std_logic;
signal \U712_CHIP_RAM.N_78\ : std_logic;
signal \U712_CHIP_RAM.N_67\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_135\ : std_logic;
signal \U712_CHIP_RAM.N_122\ : std_logic;
signal \U712_CHIP_RAM.N_135_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_121\ : std_logic;
signal \U712_CHIP_RAM.N_66\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_61\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \RnW_c\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_47\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_63\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_63_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER46\ : std_logic;
signal \U712_CHIP_RAM.N_127\ : std_logic;
signal \U712_CHIP_RAM.N_124\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_107\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \CLKEN_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    CLKEN <= \CLKEN_wire\;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    LDSn <= \LDSn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_OUT_i\,
            REFERENCECLK => \N__3610\,
            RESETB => \N__9217\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_OUT\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10331\,
            DIN => \N__10330\,
            DOUT => \N__10329\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10331\,
            PADOUT => \N__10330\,
            PADIN => \N__10329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5788\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10322\,
            DIN => \N__10321\,
            DOUT => \N__10320\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10322\,
            PADOUT => \N__10321\,
            PADIN => \N__10320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10313\,
            DIN => \N__10312\,
            DOUT => \N__10311\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10313\,
            PADOUT => \N__10312\,
            PADIN => \N__10311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8566\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10304\,
            DIN => \N__10303\,
            DOUT => \N__10302\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10304\,
            PADOUT => \N__10303\,
            PADIN => \N__10302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7435\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10295\,
            DIN => \N__10294\,
            DOUT => \N__10293\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10295\,
            PADOUT => \N__10294\,
            PADIN => \N__10293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKEN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10286\,
            DIN => \N__10285\,
            DOUT => \N__10284\,
            PACKAGEPIN => \CLKEN_wire\
        );

    \CLKEN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10286\,
            PADOUT => \N__10285\,
            PADIN => \N__10284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9213\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10277\,
            DIN => \N__10276\,
            DOUT => \N__10275\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10277\,
            PADOUT => \N__10276\,
            PADIN => \N__10275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10268\,
            DIN => \N__10267\,
            DOUT => \N__10266\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10268\,
            PADOUT => \N__10267\,
            PADIN => \N__10266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10259\,
            DIN => \N__10258\,
            DOUT => \N__10257\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10259\,
            PADOUT => \N__10258\,
            PADIN => \N__10257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10250\,
            DIN => \N__10249\,
            DOUT => \N__10248\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10250\,
            PADOUT => \N__10249\,
            PADIN => \N__10248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10241\,
            DIN => \N__10240\,
            DOUT => \N__10239\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10241\,
            PADOUT => \N__10240\,
            PADIN => \N__10239\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10232\,
            DIN => \N__10231\,
            DOUT => \N__10230\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10232\,
            PADOUT => \N__10231\,
            PADIN => \N__10230\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6205\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10223\,
            DIN => \N__10222\,
            DOUT => \N__10221\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10223\,
            PADOUT => \N__10222\,
            PADIN => \N__10221\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4290\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10214\,
            DIN => \N__10213\,
            DOUT => \N__10212\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10214\,
            PADOUT => \N__10213\,
            PADIN => \N__10212\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10205\,
            DIN => \N__10204\,
            DOUT => \N__10203\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10205\,
            PADOUT => \N__10204\,
            PADIN => \N__10203\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10196\,
            DIN => \N__10195\,
            DOUT => \N__10194\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10196\,
            PADOUT => \N__10195\,
            PADIN => \N__10194\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3799\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10187\,
            DIN => \N__10186\,
            DOUT => \N__10185\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10187\,
            PADOUT => \N__10186\,
            PADIN => \N__10185\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10178\,
            DIN => \N__10177\,
            DOUT => \N__10176\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10178\,
            PADOUT => \N__10177\,
            PADIN => \N__10176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10169\,
            DIN => \N__10168\,
            DOUT => \N__10167\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10169\,
            PADOUT => \N__10168\,
            PADIN => \N__10167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4615\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10160\,
            DIN => \N__10159\,
            DOUT => \N__10158\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10160\,
            PADOUT => \N__10159\,
            PADIN => \N__10158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10151\,
            DIN => \N__10150\,
            DOUT => \N__10149\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10151\,
            PADOUT => \N__10150\,
            PADIN => \N__10149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8839\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10142\,
            DIN => \N__10141\,
            DOUT => \N__10140\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10142\,
            PADOUT => \N__10141\,
            PADIN => \N__10140\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10133\,
            DIN => \N__10132\,
            DOUT => \N__10131\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10133\,
            PADOUT => \N__10132\,
            PADIN => \N__10131\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10124\,
            DIN => \N__10123\,
            DOUT => \N__10122\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10124\,
            PADOUT => \N__10123\,
            PADIN => \N__10122\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10115\,
            DIN => \N__10114\,
            DOUT => \N__10113\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10115\,
            PADOUT => \N__10114\,
            PADIN => \N__10113\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10106\,
            DIN => \N__10105\,
            DOUT => \N__10104\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10106\,
            PADOUT => \N__10105\,
            PADIN => \N__10104\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10097\,
            DIN => \N__10096\,
            DOUT => \N__10095\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10097\,
            PADOUT => \N__10096\,
            PADIN => \N__10095\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10088\,
            DIN => \N__10087\,
            DOUT => \N__10086\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10088\,
            PADOUT => \N__10087\,
            PADIN => \N__10086\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10079\,
            DIN => \N__10078\,
            DOUT => \N__10077\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10079\,
            PADOUT => \N__10078\,
            PADIN => \N__10077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10070\,
            DIN => \N__10069\,
            DOUT => \N__10068\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10070\,
            PADOUT => \N__10069\,
            PADIN => \N__10068\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10061\,
            DIN => \N__10060\,
            DOUT => \N__10059\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10061\,
            PADOUT => \N__10060\,
            PADIN => \N__10059\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10052\,
            DIN => \N__10051\,
            DOUT => \N__10050\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10052\,
            PADOUT => \N__10051\,
            PADIN => \N__10050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5932\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10043\,
            DIN => \N__10042\,
            DOUT => \N__10041\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10043\,
            PADOUT => \N__10042\,
            PADIN => \N__10041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10034\,
            DIN => \N__10033\,
            DOUT => \N__10032\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10034\,
            PADOUT => \N__10033\,
            PADIN => \N__10032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10025\,
            DIN => \N__10024\,
            DOUT => \N__10023\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10025\,
            PADOUT => \N__10024\,
            PADIN => \N__10023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10016\,
            DIN => \N__10015\,
            DOUT => \N__10014\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10016\,
            PADOUT => \N__10015\,
            PADIN => \N__10014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10007\,
            DIN => \N__10006\,
            DOUT => \N__10005\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10007\,
            PADOUT => \N__10006\,
            PADIN => \N__10005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3685\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9998\,
            DIN => \N__9997\,
            DOUT => \N__9996\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9998\,
            PADOUT => \N__9997\,
            PADIN => \N__9996\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6271\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9989\,
            DIN => \N__9988\,
            DOUT => \N__9987\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9989\,
            PADOUT => \N__9988\,
            PADIN => \N__9987\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9980\,
            DIN => \N__9979\,
            DOUT => \N__9978\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9980\,
            PADOUT => \N__9979\,
            PADIN => \N__9978\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8722\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9971\,
            DIN => \N__9970\,
            DOUT => \N__9969\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9971\,
            PADOUT => \N__9970\,
            PADIN => \N__9969\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9962\,
            DIN => \N__9961\,
            DOUT => \N__9960\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9962\,
            PADOUT => \N__9961\,
            PADIN => \N__9960\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9953\,
            DIN => \N__9952\,
            DOUT => \N__9951\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9953\,
            PADOUT => \N__9952\,
            PADIN => \N__9951\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3625\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9944\,
            DIN => \N__9943\,
            DOUT => \N__9942\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9944\,
            PADOUT => \N__9943\,
            PADIN => \N__9942\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9935\,
            DIN => \N__9934\,
            DOUT => \N__9933\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9935\,
            PADOUT => \N__9934\,
            PADIN => \N__9933\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4429\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9926\,
            DIN => \N__9925\,
            DOUT => \N__9924\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9926\,
            PADOUT => \N__9925\,
            PADIN => \N__9924\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5368\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9917\,
            DIN => \N__9916\,
            DOUT => \N__9915\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9917\,
            PADOUT => \N__9916\,
            PADIN => \N__9915\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9908\,
            DIN => \N__9907\,
            DOUT => \N__9906\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9908\,
            PADOUT => \N__9907\,
            PADIN => \N__9906\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9899\,
            DIN => \N__9898\,
            DOUT => \N__9897\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9899\,
            PADOUT => \N__9898\,
            PADIN => \N__9897\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9890\,
            DIN => \N__9889\,
            DOUT => \N__9888\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9890\,
            PADOUT => \N__9889\,
            PADIN => \N__9888\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7414\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9881\,
            DIN => \N__9880\,
            DOUT => \N__9879\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9881\,
            PADOUT => \N__9880\,
            PADIN => \N__9879\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9872\,
            DIN => \N__9871\,
            DOUT => \N__9870\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9872\,
            PADOUT => \N__9871\,
            PADIN => \N__9870\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5302\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9863\,
            DIN => \N__9862\,
            DOUT => \N__9861\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9863\,
            PADOUT => \N__9862\,
            PADIN => \N__9861\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9085\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9854\,
            DIN => \N__9853\,
            DOUT => \N__9852\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9854\,
            PADOUT => \N__9853\,
            PADIN => \N__9852\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5554\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9845\,
            DIN => \N__9844\,
            DOUT => \N__9843\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9845\,
            PADOUT => \N__9844\,
            PADIN => \N__9843\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5881\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9836\,
            DIN => \N__9835\,
            DOUT => \N__9834\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9836\,
            PADOUT => \N__9835\,
            PADIN => \N__9834\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4428\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9827\,
            DIN => \N__9826\,
            DOUT => \N__9825\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9827\,
            PADOUT => \N__9826\,
            PADIN => \N__9825\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9818\,
            DIN => \N__9817\,
            DOUT => \N__9816\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9818\,
            PADOUT => \N__9817\,
            PADIN => \N__9816\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9809\,
            DIN => \N__9808\,
            DOUT => \N__9807\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9809\,
            PADOUT => \N__9808\,
            PADIN => \N__9807\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5530\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9800\,
            DIN => \N__9799\,
            DOUT => \N__9798\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9800\,
            PADOUT => \N__9799\,
            PADIN => \N__9798\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8431\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9791\,
            DIN => \N__9790\,
            DOUT => \N__9789\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9791\,
            PADOUT => \N__9790\,
            PADIN => \N__9789\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7477\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9782\,
            DIN => \N__9781\,
            DOUT => \N__9780\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9782\,
            PADOUT => \N__9781\,
            PADIN => \N__9780\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5590\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9773\,
            DIN => \N__9772\,
            DOUT => \N__9771\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9773\,
            PADOUT => \N__9772\,
            PADIN => \N__9771\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9764\,
            DIN => \N__9763\,
            DOUT => \N__9762\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9764\,
            PADOUT => \N__9763\,
            PADIN => \N__9762\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9755\,
            DIN => \N__9754\,
            DOUT => \N__9753\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9755\,
            PADOUT => \N__9754\,
            PADIN => \N__9753\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9746\,
            DIN => \N__9745\,
            DOUT => \N__9744\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9746\,
            PADOUT => \N__9745\,
            PADIN => \N__9744\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9737\,
            DIN => \N__9736\,
            DOUT => \N__9735\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9737\,
            PADOUT => \N__9736\,
            PADIN => \N__9735\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4594\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9728\,
            DIN => \N__9727\,
            DOUT => \N__9726\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9728\,
            PADOUT => \N__9727\,
            PADIN => \N__9726\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9719\,
            DIN => \N__9718\,
            DOUT => \N__9717\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9719\,
            PADOUT => \N__9718\,
            PADIN => \N__9717\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5746\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9710\,
            DIN => \N__9709\,
            DOUT => \N__9708\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9710\,
            PADOUT => \N__9709\,
            PADIN => \N__9708\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3649\,
            DIN0 => OPEN,
            DOUT0 => \N__3736\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9701\,
            DIN => \N__9700\,
            DOUT => \N__9699\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9701\,
            PADOUT => \N__9700\,
            PADIN => \N__9699\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4582\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9692\,
            DIN => \N__9691\,
            DOUT => \N__9690\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9692\,
            PADOUT => \N__9691\,
            PADIN => \N__9690\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9683\,
            DIN => \N__9682\,
            DOUT => \N__9681\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9683\,
            PADOUT => \N__9682\,
            PADIN => \N__9681\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9674\,
            DIN => \N__9673\,
            DOUT => \N__9672\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9674\,
            PADOUT => \N__9673\,
            PADIN => \N__9672\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5962\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9665\,
            DIN => \N__9664\,
            DOUT => \N__9663\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9665\,
            PADOUT => \N__9664\,
            PADIN => \N__9663\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9656\,
            DIN => \N__9655\,
            DOUT => \N__9654\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9656\,
            PADOUT => \N__9655\,
            PADIN => \N__9654\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9647\,
            DIN => \N__9646\,
            DOUT => \N__9645\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9647\,
            PADOUT => \N__9646\,
            PADIN => \N__9645\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9638\,
            DIN => \N__9637\,
            DOUT => \N__9636\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9638\,
            PADOUT => \N__9637\,
            PADIN => \N__9636\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9629\,
            DIN => \N__9628\,
            DOUT => \N__9627\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9629\,
            PADOUT => \N__9628\,
            PADIN => \N__9627\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5206\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9620\,
            DIN => \N__9619\,
            DOUT => \N__9618\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9620\,
            PADOUT => \N__9619\,
            PADIN => \N__9618\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4852\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2307\ : InMux
    port map (
            O => \N__9601\,
            I => \N__9598\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__9598\,
            I => \N__9595\
        );

    \I__2305\ : Odrv12
    port map (
            O => \N__9595\,
            I => \RAS1n_c\
        );

    \I__2304\ : InMux
    port map (
            O => \N__9592\,
            I => \N__9588\
        );

    \I__2303\ : InMux
    port map (
            O => \N__9591\,
            I => \N__9585\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__9588\,
            I => \N__9582\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__9585\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2300\ : Odrv4
    port map (
            O => \N__9582\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2299\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9574\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__9574\,
            I => \N__9535\
        );

    \I__2297\ : ClkMux
    port map (
            O => \N__9573\,
            I => \N__9421\
        );

    \I__2296\ : ClkMux
    port map (
            O => \N__9572\,
            I => \N__9421\
        );

    \I__2295\ : ClkMux
    port map (
            O => \N__9571\,
            I => \N__9421\
        );

    \I__2294\ : ClkMux
    port map (
            O => \N__9570\,
            I => \N__9421\
        );

    \I__2293\ : ClkMux
    port map (
            O => \N__9569\,
            I => \N__9421\
        );

    \I__2292\ : ClkMux
    port map (
            O => \N__9568\,
            I => \N__9421\
        );

    \I__2291\ : ClkMux
    port map (
            O => \N__9567\,
            I => \N__9421\
        );

    \I__2290\ : ClkMux
    port map (
            O => \N__9566\,
            I => \N__9421\
        );

    \I__2289\ : ClkMux
    port map (
            O => \N__9565\,
            I => \N__9421\
        );

    \I__2288\ : ClkMux
    port map (
            O => \N__9564\,
            I => \N__9421\
        );

    \I__2287\ : ClkMux
    port map (
            O => \N__9563\,
            I => \N__9421\
        );

    \I__2286\ : ClkMux
    port map (
            O => \N__9562\,
            I => \N__9421\
        );

    \I__2285\ : ClkMux
    port map (
            O => \N__9561\,
            I => \N__9421\
        );

    \I__2284\ : ClkMux
    port map (
            O => \N__9560\,
            I => \N__9421\
        );

    \I__2283\ : ClkMux
    port map (
            O => \N__9559\,
            I => \N__9421\
        );

    \I__2282\ : ClkMux
    port map (
            O => \N__9558\,
            I => \N__9421\
        );

    \I__2281\ : ClkMux
    port map (
            O => \N__9557\,
            I => \N__9421\
        );

    \I__2280\ : ClkMux
    port map (
            O => \N__9556\,
            I => \N__9421\
        );

    \I__2279\ : ClkMux
    port map (
            O => \N__9555\,
            I => \N__9421\
        );

    \I__2278\ : ClkMux
    port map (
            O => \N__9554\,
            I => \N__9421\
        );

    \I__2277\ : ClkMux
    port map (
            O => \N__9553\,
            I => \N__9421\
        );

    \I__2276\ : ClkMux
    port map (
            O => \N__9552\,
            I => \N__9421\
        );

    \I__2275\ : ClkMux
    port map (
            O => \N__9551\,
            I => \N__9421\
        );

    \I__2274\ : ClkMux
    port map (
            O => \N__9550\,
            I => \N__9421\
        );

    \I__2273\ : ClkMux
    port map (
            O => \N__9549\,
            I => \N__9421\
        );

    \I__2272\ : ClkMux
    port map (
            O => \N__9548\,
            I => \N__9421\
        );

    \I__2271\ : ClkMux
    port map (
            O => \N__9547\,
            I => \N__9421\
        );

    \I__2270\ : ClkMux
    port map (
            O => \N__9546\,
            I => \N__9421\
        );

    \I__2269\ : ClkMux
    port map (
            O => \N__9545\,
            I => \N__9421\
        );

    \I__2268\ : ClkMux
    port map (
            O => \N__9544\,
            I => \N__9421\
        );

    \I__2267\ : ClkMux
    port map (
            O => \N__9543\,
            I => \N__9421\
        );

    \I__2266\ : ClkMux
    port map (
            O => \N__9542\,
            I => \N__9421\
        );

    \I__2265\ : ClkMux
    port map (
            O => \N__9541\,
            I => \N__9421\
        );

    \I__2264\ : ClkMux
    port map (
            O => \N__9540\,
            I => \N__9421\
        );

    \I__2263\ : ClkMux
    port map (
            O => \N__9539\,
            I => \N__9421\
        );

    \I__2262\ : ClkMux
    port map (
            O => \N__9538\,
            I => \N__9421\
        );

    \I__2261\ : Glb2LocalMux
    port map (
            O => \N__9535\,
            I => \N__9421\
        );

    \I__2260\ : ClkMux
    port map (
            O => \N__9534\,
            I => \N__9421\
        );

    \I__2259\ : ClkMux
    port map (
            O => \N__9533\,
            I => \N__9421\
        );

    \I__2258\ : ClkMux
    port map (
            O => \N__9532\,
            I => \N__9421\
        );

    \I__2257\ : ClkMux
    port map (
            O => \N__9531\,
            I => \N__9421\
        );

    \I__2256\ : ClkMux
    port map (
            O => \N__9530\,
            I => \N__9421\
        );

    \I__2255\ : ClkMux
    port map (
            O => \N__9529\,
            I => \N__9421\
        );

    \I__2254\ : ClkMux
    port map (
            O => \N__9528\,
            I => \N__9421\
        );

    \I__2253\ : ClkMux
    port map (
            O => \N__9527\,
            I => \N__9421\
        );

    \I__2252\ : ClkMux
    port map (
            O => \N__9526\,
            I => \N__9421\
        );

    \I__2251\ : ClkMux
    port map (
            O => \N__9525\,
            I => \N__9421\
        );

    \I__2250\ : ClkMux
    port map (
            O => \N__9524\,
            I => \N__9421\
        );

    \I__2249\ : ClkMux
    port map (
            O => \N__9523\,
            I => \N__9421\
        );

    \I__2248\ : ClkMux
    port map (
            O => \N__9522\,
            I => \N__9421\
        );

    \I__2247\ : GlobalMux
    port map (
            O => \N__9421\,
            I => \CLK80_OUT\
        );

    \I__2246\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9406\
        );

    \I__2245\ : InMux
    port map (
            O => \N__9417\,
            I => \N__9403\
        );

    \I__2244\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9400\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9391\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9391\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9391\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9391\
        );

    \I__2239\ : InMux
    port map (
            O => \N__9411\,
            I => \N__9388\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9385\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9382\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__9406\,
            I => \N__9371\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__9403\,
            I => \N__9360\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__9400\,
            I => \N__9346\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__9391\,
            I => \N__9341\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__9388\,
            I => \N__9335\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9385\,
            I => \N__9332\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__9382\,
            I => \N__9325\
        );

    \I__2229\ : SRMux
    port map (
            O => \N__9381\,
            I => \N__9223\
        );

    \I__2228\ : SRMux
    port map (
            O => \N__9380\,
            I => \N__9223\
        );

    \I__2227\ : SRMux
    port map (
            O => \N__9379\,
            I => \N__9223\
        );

    \I__2226\ : SRMux
    port map (
            O => \N__9378\,
            I => \N__9223\
        );

    \I__2225\ : SRMux
    port map (
            O => \N__9377\,
            I => \N__9223\
        );

    \I__2224\ : SRMux
    port map (
            O => \N__9376\,
            I => \N__9223\
        );

    \I__2223\ : SRMux
    port map (
            O => \N__9375\,
            I => \N__9223\
        );

    \I__2222\ : SRMux
    port map (
            O => \N__9374\,
            I => \N__9223\
        );

    \I__2221\ : Glb2LocalMux
    port map (
            O => \N__9371\,
            I => \N__9223\
        );

    \I__2220\ : SRMux
    port map (
            O => \N__9370\,
            I => \N__9223\
        );

    \I__2219\ : SRMux
    port map (
            O => \N__9369\,
            I => \N__9223\
        );

    \I__2218\ : SRMux
    port map (
            O => \N__9368\,
            I => \N__9223\
        );

    \I__2217\ : SRMux
    port map (
            O => \N__9367\,
            I => \N__9223\
        );

    \I__2216\ : SRMux
    port map (
            O => \N__9366\,
            I => \N__9223\
        );

    \I__2215\ : SRMux
    port map (
            O => \N__9365\,
            I => \N__9223\
        );

    \I__2214\ : SRMux
    port map (
            O => \N__9364\,
            I => \N__9223\
        );

    \I__2213\ : SRMux
    port map (
            O => \N__9363\,
            I => \N__9223\
        );

    \I__2212\ : Glb2LocalMux
    port map (
            O => \N__9360\,
            I => \N__9223\
        );

    \I__2211\ : SRMux
    port map (
            O => \N__9359\,
            I => \N__9223\
        );

    \I__2210\ : SRMux
    port map (
            O => \N__9358\,
            I => \N__9223\
        );

    \I__2209\ : SRMux
    port map (
            O => \N__9357\,
            I => \N__9223\
        );

    \I__2208\ : SRMux
    port map (
            O => \N__9356\,
            I => \N__9223\
        );

    \I__2207\ : SRMux
    port map (
            O => \N__9355\,
            I => \N__9223\
        );

    \I__2206\ : SRMux
    port map (
            O => \N__9354\,
            I => \N__9223\
        );

    \I__2205\ : SRMux
    port map (
            O => \N__9353\,
            I => \N__9223\
        );

    \I__2204\ : SRMux
    port map (
            O => \N__9352\,
            I => \N__9223\
        );

    \I__2203\ : SRMux
    port map (
            O => \N__9351\,
            I => \N__9223\
        );

    \I__2202\ : SRMux
    port map (
            O => \N__9350\,
            I => \N__9223\
        );

    \I__2201\ : SRMux
    port map (
            O => \N__9349\,
            I => \N__9223\
        );

    \I__2200\ : Glb2LocalMux
    port map (
            O => \N__9346\,
            I => \N__9223\
        );

    \I__2199\ : SRMux
    port map (
            O => \N__9345\,
            I => \N__9223\
        );

    \I__2198\ : SRMux
    port map (
            O => \N__9344\,
            I => \N__9223\
        );

    \I__2197\ : Glb2LocalMux
    port map (
            O => \N__9341\,
            I => \N__9223\
        );

    \I__2196\ : SRMux
    port map (
            O => \N__9340\,
            I => \N__9223\
        );

    \I__2195\ : SRMux
    port map (
            O => \N__9339\,
            I => \N__9223\
        );

    \I__2194\ : SRMux
    port map (
            O => \N__9338\,
            I => \N__9223\
        );

    \I__2193\ : Glb2LocalMux
    port map (
            O => \N__9335\,
            I => \N__9223\
        );

    \I__2192\ : Glb2LocalMux
    port map (
            O => \N__9332\,
            I => \N__9223\
        );

    \I__2191\ : SRMux
    port map (
            O => \N__9331\,
            I => \N__9223\
        );

    \I__2190\ : SRMux
    port map (
            O => \N__9330\,
            I => \N__9223\
        );

    \I__2189\ : SRMux
    port map (
            O => \N__9329\,
            I => \N__9223\
        );

    \I__2188\ : SRMux
    port map (
            O => \N__9328\,
            I => \N__9223\
        );

    \I__2187\ : Glb2LocalMux
    port map (
            O => \N__9325\,
            I => \N__9223\
        );

    \I__2186\ : SRMux
    port map (
            O => \N__9324\,
            I => \N__9223\
        );

    \I__2185\ : SRMux
    port map (
            O => \N__9323\,
            I => \N__9223\
        );

    \I__2184\ : SRMux
    port map (
            O => \N__9322\,
            I => \N__9223\
        );

    \I__2183\ : SRMux
    port map (
            O => \N__9321\,
            I => \N__9223\
        );

    \I__2182\ : SRMux
    port map (
            O => \N__9320\,
            I => \N__9223\
        );

    \I__2181\ : GlobalMux
    port map (
            O => \N__9223\,
            I => \N__9220\
        );

    \I__2180\ : gio2CtrlBuf
    port map (
            O => \N__9220\,
            I => \RESETn_c_i_g\
        );

    \I__2179\ : IoInMux
    port map (
            O => \N__9217\,
            I => \N__9214\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9214\,
            I => \N__9210\
        );

    \I__2177\ : IoInMux
    port map (
            O => \N__9213\,
            I => \N__9207\
        );

    \I__2176\ : Span4Mux_s3_v
    port map (
            O => \N__9210\,
            I => \N__9204\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__9207\,
            I => \N__9201\
        );

    \I__2174\ : Span4Mux_v
    port map (
            O => \N__9204\,
            I => \N__9198\
        );

    \I__2173\ : Span4Mux_s3_h
    port map (
            O => \N__9201\,
            I => \N__9195\
        );

    \I__2172\ : Span4Mux_h
    port map (
            O => \N__9198\,
            I => \N__9192\
        );

    \I__2171\ : Span4Mux_h
    port map (
            O => \N__9195\,
            I => \N__9189\
        );

    \I__2170\ : Odrv4
    port map (
            O => \N__9192\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__9189\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9184\,
            I => \N__9181\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9181\,
            I => \N__9177\
        );

    \I__2166\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9174\
        );

    \I__2165\ : Span4Mux_h
    port map (
            O => \N__9177\,
            I => \N__9168\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9174\,
            I => \N__9168\
        );

    \I__2163\ : InMux
    port map (
            O => \N__9173\,
            I => \N__9165\
        );

    \I__2162\ : Span4Mux_v
    port map (
            O => \N__9168\,
            I => \N__9162\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__9165\,
            I => \N__9159\
        );

    \I__2160\ : Sp12to4
    port map (
            O => \N__9162\,
            I => \N__9155\
        );

    \I__2159\ : Span4Mux_v
    port map (
            O => \N__9159\,
            I => \N__9152\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9149\
        );

    \I__2157\ : Odrv12
    port map (
            O => \N__9155\,
            I => \REG_CYCLEm\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__9152\,
            I => \REG_CYCLEm\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9149\,
            I => \REG_CYCLEm\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9142\,
            I => \N__9136\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9141\,
            I => \N__9133\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9140\,
            I => \N__9130\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9139\,
            I => \N__9127\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__9136\,
            I => \N__9119\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__9133\,
            I => \N__9114\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9130\,
            I => \N__9114\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__9127\,
            I => \N__9111\
        );

    \I__2146\ : InMux
    port map (
            O => \N__9126\,
            I => \N__9102\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9125\,
            I => \N__9102\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9124\,
            I => \N__9102\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9102\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9099\
        );

    \I__2141\ : Span4Mux_v
    port map (
            O => \N__9119\,
            I => \N__9094\
        );

    \I__2140\ : Span4Mux_v
    port map (
            O => \N__9114\,
            I => \N__9094\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__9111\,
            I => \DMA_CYCLEm\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9102\,
            I => \DMA_CYCLEm\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9099\,
            I => \DMA_CYCLEm\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__9094\,
            I => \DMA_CYCLEm\
        );

    \I__2135\ : IoInMux
    port map (
            O => \N__9085\,
            I => \N__9082\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9082\,
            I => \N__9079\
        );

    \I__2133\ : IoSpan4Mux
    port map (
            O => \N__9079\,
            I => \N__9076\
        );

    \I__2132\ : Sp12to4
    port map (
            O => \N__9076\,
            I => \N__9073\
        );

    \I__2131\ : Span12Mux_v
    port map (
            O => \N__9073\,
            I => \N__9070\
        );

    \I__2130\ : Span12Mux_h
    port map (
            O => \N__9070\,
            I => \N__9067\
        );

    \I__2129\ : Odrv12
    port map (
            O => \N__9067\,
            I => \DRDENn_c\
        );

    \I__2128\ : CEMux
    port map (
            O => \N__9064\,
            I => \N__9060\
        );

    \I__2127\ : CEMux
    port map (
            O => \N__9063\,
            I => \N__9055\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__9060\,
            I => \N__9052\
        );

    \I__2125\ : CEMux
    port map (
            O => \N__9059\,
            I => \N__9049\
        );

    \I__2124\ : CEMux
    port map (
            O => \N__9058\,
            I => \N__9046\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__9055\,
            I => \N__9042\
        );

    \I__2122\ : Span4Mux_h
    port map (
            O => \N__9052\,
            I => \N__9037\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__9049\,
            I => \N__9037\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9046\,
            I => \N__9034\
        );

    \I__2119\ : CEMux
    port map (
            O => \N__9045\,
            I => \N__9031\
        );

    \I__2118\ : Span4Mux_v
    port map (
            O => \N__9042\,
            I => \N__9028\
        );

    \I__2117\ : Span4Mux_v
    port map (
            O => \N__9037\,
            I => \N__9023\
        );

    \I__2116\ : Span4Mux_v
    port map (
            O => \N__9034\,
            I => \N__9023\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9031\,
            I => \N__9020\
        );

    \I__2114\ : Span4Mux_h
    port map (
            O => \N__9028\,
            I => \N__9017\
        );

    \I__2113\ : Span4Mux_h
    port map (
            O => \N__9023\,
            I => \N__9012\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__9020\,
            I => \N__9012\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__9017\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__9012\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__2109\ : InMux
    port map (
            O => \N__9007\,
            I => \N__9004\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__9004\,
            I => \N__9000\
        );

    \I__2107\ : InMux
    port map (
            O => \N__9003\,
            I => \N__8997\
        );

    \I__2106\ : Span4Mux_v
    port map (
            O => \N__9000\,
            I => \N__8994\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__8997\,
            I => \N__8991\
        );

    \I__2104\ : Sp12to4
    port map (
            O => \N__8994\,
            I => \N__8988\
        );

    \I__2103\ : Span4Mux_h
    port map (
            O => \N__8991\,
            I => \N__8985\
        );

    \I__2102\ : Span12Mux_h
    port map (
            O => \N__8988\,
            I => \N__8982\
        );

    \I__2101\ : Sp12to4
    port map (
            O => \N__8985\,
            I => \N__8979\
        );

    \I__2100\ : Span12Mux_v
    port map (
            O => \N__8982\,
            I => \N__8976\
        );

    \I__2099\ : Span12Mux_v
    port map (
            O => \N__8979\,
            I => \N__8973\
        );

    \I__2098\ : Odrv12
    port map (
            O => \N__8976\,
            I => \DRA_c_0\
        );

    \I__2097\ : Odrv12
    port map (
            O => \N__8973\,
            I => \DRA_c_0\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__8968\,
            I => \N__8965\
        );

    \I__2095\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8962\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__8962\,
            I => \N__8959\
        );

    \I__2093\ : Span12Mux_v
    port map (
            O => \N__8959\,
            I => \N__8956\
        );

    \I__2092\ : Odrv12
    port map (
            O => \N__8956\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2091\ : CEMux
    port map (
            O => \N__8953\,
            I => \N__8949\
        );

    \I__2090\ : CEMux
    port map (
            O => \N__8952\,
            I => \N__8946\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__8949\,
            I => \N__8942\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__8946\,
            I => \N__8939\
        );

    \I__2087\ : CEMux
    port map (
            O => \N__8945\,
            I => \N__8936\
        );

    \I__2086\ : Span4Mux_h
    port map (
            O => \N__8942\,
            I => \N__8927\
        );

    \I__2085\ : Span4Mux_h
    port map (
            O => \N__8939\,
            I => \N__8927\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__8936\,
            I => \N__8927\
        );

    \I__2083\ : CEMux
    port map (
            O => \N__8935\,
            I => \N__8924\
        );

    \I__2082\ : CEMux
    port map (
            O => \N__8934\,
            I => \N__8921\
        );

    \I__2081\ : Span4Mux_v
    port map (
            O => \N__8927\,
            I => \N__8917\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__8924\,
            I => \N__8914\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__8921\,
            I => \N__8911\
        );

    \I__2078\ : CEMux
    port map (
            O => \N__8920\,
            I => \N__8908\
        );

    \I__2077\ : Span4Mux_h
    port map (
            O => \N__8917\,
            I => \N__8905\
        );

    \I__2076\ : Span4Mux_h
    port map (
            O => \N__8914\,
            I => \N__8902\
        );

    \I__2075\ : Span4Mux_h
    port map (
            O => \N__8911\,
            I => \N__8899\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__8908\,
            I => \N__8896\
        );

    \I__2073\ : Odrv4
    port map (
            O => \N__8905\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__8902\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__2071\ : Odrv4
    port map (
            O => \N__8899\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__2070\ : Odrv12
    port map (
            O => \N__8896\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__2069\ : InMux
    port map (
            O => \N__8887\,
            I => \N__8883\
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__8886\,
            I => \N__8880\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__8883\,
            I => \N__8876\
        );

    \I__2066\ : InMux
    port map (
            O => \N__8880\,
            I => \N__8873\
        );

    \I__2065\ : InMux
    port map (
            O => \N__8879\,
            I => \N__8870\
        );

    \I__2064\ : Span4Mux_v
    port map (
            O => \N__8876\,
            I => \N__8867\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__8873\,
            I => \N__8861\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__8870\,
            I => \N__8861\
        );

    \I__2061\ : Span4Mux_v
    port map (
            O => \N__8867\,
            I => \N__8858\
        );

    \I__2060\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8855\
        );

    \I__2059\ : Span4Mux_h
    port map (
            O => \N__8861\,
            I => \N__8852\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__8858\,
            I => \N__8847\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__8855\,
            I => \N__8847\
        );

    \I__2056\ : Span4Mux_v
    port map (
            O => \N__8852\,
            I => \N__8844\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__8847\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__8844\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2053\ : IoInMux
    port map (
            O => \N__8839\,
            I => \N__8836\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__8836\,
            I => \N__8833\
        );

    \I__2051\ : Span4Mux_s1_v
    port map (
            O => \N__8833\,
            I => \N__8830\
        );

    \I__2050\ : Span4Mux_v
    port map (
            O => \N__8830\,
            I => \N__8827\
        );

    \I__2049\ : Span4Mux_v
    port map (
            O => \N__8827\,
            I => \N__8824\
        );

    \I__2048\ : Odrv4
    port map (
            O => \N__8824\,
            I => \CRCSn_c\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__8821\,
            I => \N__8813\
        );

    \I__2046\ : InMux
    port map (
            O => \N__8820\,
            I => \N__8808\
        );

    \I__2045\ : InMux
    port map (
            O => \N__8819\,
            I => \N__8805\
        );

    \I__2044\ : InMux
    port map (
            O => \N__8818\,
            I => \N__8802\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__8817\,
            I => \N__8797\
        );

    \I__2042\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8794\
        );

    \I__2041\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8787\
        );

    \I__2040\ : InMux
    port map (
            O => \N__8812\,
            I => \N__8787\
        );

    \I__2039\ : InMux
    port map (
            O => \N__8811\,
            I => \N__8787\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__8808\,
            I => \N__8782\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__8805\,
            I => \N__8782\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__8802\,
            I => \N__8778\
        );

    \I__2035\ : InMux
    port map (
            O => \N__8801\,
            I => \N__8773\
        );

    \I__2034\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8773\
        );

    \I__2033\ : InMux
    port map (
            O => \N__8797\,
            I => \N__8770\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__8794\,
            I => \N__8761\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__8787\,
            I => \N__8761\
        );

    \I__2030\ : Span4Mux_h
    port map (
            O => \N__8782\,
            I => \N__8761\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__8781\,
            I => \N__8758\
        );

    \I__2028\ : Span4Mux_v
    port map (
            O => \N__8778\,
            I => \N__8755\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__8773\,
            I => \N__8750\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__8770\,
            I => \N__8750\
        );

    \I__2025\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8747\
        );

    \I__2024\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8744\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__8761\,
            I => \N__8741\
        );

    \I__2022\ : InMux
    port map (
            O => \N__8758\,
            I => \N__8738\
        );

    \I__2021\ : Span4Mux_h
    port map (
            O => \N__8755\,
            I => \N__8733\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__8750\,
            I => \N__8733\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__8747\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__8744\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__8741\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__8738\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__8733\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2014\ : IoInMux
    port map (
            O => \N__8722\,
            I => \N__8719\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__8719\,
            I => \N__8716\
        );

    \I__2012\ : Span4Mux_s2_v
    port map (
            O => \N__8716\,
            I => \N__8713\
        );

    \I__2011\ : Span4Mux_v
    port map (
            O => \N__8713\,
            I => \N__8710\
        );

    \I__2010\ : Span4Mux_v
    port map (
            O => \N__8710\,
            I => \N__8707\
        );

    \I__2009\ : Odrv4
    port map (
            O => \N__8707\,
            I => \RASn_c\
        );

    \I__2008\ : InMux
    port map (
            O => \N__8704\,
            I => \N__8696\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__8703\,
            I => \N__8692\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__8702\,
            I => \N__8687\
        );

    \I__2005\ : InMux
    port map (
            O => \N__8701\,
            I => \N__8684\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__8700\,
            I => \N__8681\
        );

    \I__2003\ : CascadeMux
    port map (
            O => \N__8699\,
            I => \N__8677\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__8696\,
            I => \N__8673\
        );

    \I__2001\ : InMux
    port map (
            O => \N__8695\,
            I => \N__8670\
        );

    \I__2000\ : InMux
    port map (
            O => \N__8692\,
            I => \N__8667\
        );

    \I__1999\ : InMux
    port map (
            O => \N__8691\,
            I => \N__8664\
        );

    \I__1998\ : InMux
    port map (
            O => \N__8690\,
            I => \N__8660\
        );

    \I__1997\ : InMux
    port map (
            O => \N__8687\,
            I => \N__8657\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__8684\,
            I => \N__8654\
        );

    \I__1995\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8651\
        );

    \I__1994\ : InMux
    port map (
            O => \N__8680\,
            I => \N__8648\
        );

    \I__1993\ : InMux
    port map (
            O => \N__8677\,
            I => \N__8645\
        );

    \I__1992\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8641\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__8673\,
            I => \N__8638\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__8670\,
            I => \N__8633\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__8667\,
            I => \N__8633\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__8664\,
            I => \N__8630\
        );

    \I__1987\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8627\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__8660\,
            I => \N__8622\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__8657\,
            I => \N__8622\
        );

    \I__1984\ : Span4Mux_v
    port map (
            O => \N__8654\,
            I => \N__8617\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__8651\,
            I => \N__8617\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__8648\,
            I => \N__8612\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__8645\,
            I => \N__8609\
        );

    \I__1980\ : InMux
    port map (
            O => \N__8644\,
            I => \N__8606\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__8641\,
            I => \N__8603\
        );

    \I__1978\ : Span4Mux_v
    port map (
            O => \N__8638\,
            I => \N__8598\
        );

    \I__1977\ : Span4Mux_v
    port map (
            O => \N__8633\,
            I => \N__8598\
        );

    \I__1976\ : Span4Mux_h
    port map (
            O => \N__8630\,
            I => \N__8589\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__8627\,
            I => \N__8589\
        );

    \I__1974\ : Span4Mux_h
    port map (
            O => \N__8622\,
            I => \N__8589\
        );

    \I__1973\ : Span4Mux_h
    port map (
            O => \N__8617\,
            I => \N__8589\
        );

    \I__1972\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8584\
        );

    \I__1971\ : InMux
    port map (
            O => \N__8615\,
            I => \N__8584\
        );

    \I__1970\ : Span4Mux_v
    port map (
            O => \N__8612\,
            I => \N__8575\
        );

    \I__1969\ : Span4Mux_h
    port map (
            O => \N__8609\,
            I => \N__8575\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__8606\,
            I => \N__8575\
        );

    \I__1967\ : Span4Mux_v
    port map (
            O => \N__8603\,
            I => \N__8575\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__8598\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1965\ : Odrv4
    port map (
            O => \N__8589\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__8584\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__8575\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1962\ : IoInMux
    port map (
            O => \N__8566\,
            I => \N__8563\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__8563\,
            I => \N__8560\
        );

    \I__1960\ : Span4Mux_s3_v
    port map (
            O => \N__8560\,
            I => \N__8557\
        );

    \I__1959\ : Sp12to4
    port map (
            O => \N__8557\,
            I => \N__8554\
        );

    \I__1958\ : Span12Mux_s10_h
    port map (
            O => \N__8554\,
            I => \N__8551\
        );

    \I__1957\ : Odrv12
    port map (
            O => \N__8551\,
            I => \CASn_c\
        );

    \I__1956\ : InMux
    port map (
            O => \N__8548\,
            I => \N__8545\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__8545\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8542\,
            I => \N__8535\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__8541\,
            I => \N__8531\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__8540\,
            I => \N__8527\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__8539\,
            I => \N__8524\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8538\,
            I => \N__8521\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__8535\,
            I => \N__8518\
        );

    \I__1948\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8512\
        );

    \I__1947\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8507\
        );

    \I__1946\ : InMux
    port map (
            O => \N__8530\,
            I => \N__8500\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8527\,
            I => \N__8500\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8500\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__8521\,
            I => \N__8497\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__8518\,
            I => \N__8494\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8489\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8489\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8515\,
            I => \N__8486\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__8512\,
            I => \N__8483\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8511\,
            I => \N__8480\
        );

    \I__1936\ : InMux
    port map (
            O => \N__8510\,
            I => \N__8477\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__8507\,
            I => \N__8472\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__8500\,
            I => \N__8472\
        );

    \I__1933\ : Span4Mux_v
    port map (
            O => \N__8497\,
            I => \N__8469\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__8494\,
            I => \N__8460\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__8489\,
            I => \N__8460\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__8486\,
            I => \N__8460\
        );

    \I__1929\ : Span4Mux_v
    port map (
            O => \N__8483\,
            I => \N__8457\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__8480\,
            I => \N__8448\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__8477\,
            I => \N__8448\
        );

    \I__1926\ : Span4Mux_v
    port map (
            O => \N__8472\,
            I => \N__8448\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__8469\,
            I => \N__8448\
        );

    \I__1924\ : InMux
    port map (
            O => \N__8468\,
            I => \N__8443\
        );

    \I__1923\ : InMux
    port map (
            O => \N__8467\,
            I => \N__8443\
        );

    \I__1922\ : Span4Mux_v
    port map (
            O => \N__8460\,
            I => \N__8440\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__8457\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1920\ : Odrv4
    port map (
            O => \N__8448\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__8443\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__8440\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1917\ : IoInMux
    port map (
            O => \N__8431\,
            I => \N__8428\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__8428\,
            I => \N__8425\
        );

    \I__1915\ : IoSpan4Mux
    port map (
            O => \N__8425\,
            I => \N__8422\
        );

    \I__1914\ : Span4Mux_s1_h
    port map (
            O => \N__8422\,
            I => \N__8419\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__8419\,
            I => \N__8416\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__8416\,
            I => \N__8413\
        );

    \I__1911\ : Span4Mux_h
    port map (
            O => \N__8413\,
            I => \N__8410\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__8410\,
            I => \WEn_c\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8407\,
            I => \N__8404\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8404\,
            I => \N__8400\
        );

    \I__1907\ : InMux
    port map (
            O => \N__8403\,
            I => \N__8397\
        );

    \I__1906\ : Span4Mux_v
    port map (
            O => \N__8400\,
            I => \N__8394\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__8397\,
            I => \N__8391\
        );

    \I__1904\ : Span4Mux_h
    port map (
            O => \N__8394\,
            I => \N__8388\
        );

    \I__1903\ : Sp12to4
    port map (
            O => \N__8391\,
            I => \N__8385\
        );

    \I__1902\ : Sp12to4
    port map (
            O => \N__8388\,
            I => \N__8380\
        );

    \I__1901\ : Span12Mux_v
    port map (
            O => \N__8385\,
            I => \N__8380\
        );

    \I__1900\ : Odrv12
    port map (
            O => \N__8380\,
            I => \RAS0n_c\
        );

    \I__1899\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8373\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8370\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__8373\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__8370\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8358\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8358\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8363\,
            I => \N__8355\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__8358\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__8355\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8345\
        );

    \I__1889\ : InMux
    port map (
            O => \N__8349\,
            I => \N__8342\
        );

    \I__1888\ : InMux
    port map (
            O => \N__8348\,
            I => \N__8339\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8345\,
            I => \N__8336\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__8342\,
            I => \N__8333\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8339\,
            I => \N__8328\
        );

    \I__1884\ : Span4Mux_v
    port map (
            O => \N__8336\,
            I => \N__8328\
        );

    \I__1883\ : Odrv12
    port map (
            O => \N__8333\,
            I => \U712_CHIP_RAM.N_135\
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__8328\,
            I => \U712_CHIP_RAM.N_135\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8323\,
            I => \N__8317\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8322\,
            I => \N__8314\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8309\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8320\,
            I => \N__8309\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8317\,
            I => \U712_CHIP_RAM.N_122\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8314\,
            I => \U712_CHIP_RAM.N_122\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8309\,
            I => \U712_CHIP_RAM.N_122\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__8302\,
            I => \U712_CHIP_RAM.N_135_cascade_\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8299\,
            I => \N__8294\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8298\,
            I => \N__8291\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8297\,
            I => \N__8288\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8294\,
            I => \U712_CHIP_RAM.N_121\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__8291\,
            I => \U712_CHIP_RAM.N_121\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8288\,
            I => \U712_CHIP_RAM.N_121\
        );

    \I__1867\ : InMux
    port map (
            O => \N__8281\,
            I => \N__8278\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__8278\,
            I => \U712_CHIP_RAM.N_66\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__8275\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_2_cascade_\
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__8272\,
            I => \N__8268\
        );

    \I__1863\ : InMux
    port map (
            O => \N__8271\,
            I => \N__8264\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8268\,
            I => \N__8261\
        );

    \I__1861\ : InMux
    port map (
            O => \N__8267\,
            I => \N__8258\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8264\,
            I => \N__8255\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__8261\,
            I => \N__8252\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__8258\,
            I => \N__8245\
        );

    \I__1857\ : Span4Mux_h
    port map (
            O => \N__8255\,
            I => \N__8240\
        );

    \I__1856\ : Span4Mux_h
    port map (
            O => \N__8252\,
            I => \N__8240\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8251\,
            I => \N__8235\
        );

    \I__1854\ : InMux
    port map (
            O => \N__8250\,
            I => \N__8235\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8249\,
            I => \N__8232\
        );

    \I__1852\ : InMux
    port map (
            O => \N__8248\,
            I => \N__8229\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__8245\,
            I => \U712_CHIP_RAM.N_61\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__8240\,
            I => \U712_CHIP_RAM.N_61\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8235\,
            I => \U712_CHIP_RAM.N_61\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8232\,
            I => \U712_CHIP_RAM.N_61\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__8229\,
            I => \U712_CHIP_RAM.N_61\
        );

    \I__1846\ : InMux
    port map (
            O => \N__8218\,
            I => \N__8215\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8215\,
            I => \N__8211\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8208\
        );

    \I__1843\ : Span4Mux_h
    port map (
            O => \N__8211\,
            I => \N__8205\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__8208\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1841\ : Odrv4
    port map (
            O => \N__8205\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8196\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8199\,
            I => \N__8193\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8196\,
            I => \N__8190\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__8193\,
            I => \N__8186\
        );

    \I__1836\ : Span4Mux_v
    port map (
            O => \N__8190\,
            I => \N__8183\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8189\,
            I => \N__8180\
        );

    \I__1834\ : Span4Mux_v
    port map (
            O => \N__8186\,
            I => \N__8175\
        );

    \I__1833\ : Span4Mux_h
    port map (
            O => \N__8183\,
            I => \N__8170\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8180\,
            I => \N__8170\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8179\,
            I => \N__8167\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__8178\,
            I => \N__8164\
        );

    \I__1829\ : Sp12to4
    port map (
            O => \N__8175\,
            I => \N__8160\
        );

    \I__1828\ : Span4Mux_h
    port map (
            O => \N__8170\,
            I => \N__8155\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8167\,
            I => \N__8155\
        );

    \I__1826\ : InMux
    port map (
            O => \N__8164\,
            I => \N__8150\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8150\
        );

    \I__1824\ : Span12Mux_h
    port map (
            O => \N__8160\,
            I => \N__8147\
        );

    \I__1823\ : Sp12to4
    port map (
            O => \N__8155\,
            I => \N__8142\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__8150\,
            I => \N__8142\
        );

    \I__1821\ : Span12Mux_h
    port map (
            O => \N__8147\,
            I => \N__8139\
        );

    \I__1820\ : Span12Mux_v
    port map (
            O => \N__8142\,
            I => \N__8136\
        );

    \I__1819\ : Span12Mux_v
    port map (
            O => \N__8139\,
            I => \N__8131\
        );

    \I__1818\ : Span12Mux_h
    port map (
            O => \N__8136\,
            I => \N__8131\
        );

    \I__1817\ : Odrv12
    port map (
            O => \N__8131\,
            I => \RnW_c\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__8128\,
            I => \N__8124\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8127\,
            I => \N__8113\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8110\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8123\,
            I => \N__8106\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__8122\,
            I => \N__8100\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__8121\,
            I => \N__8093\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8120\,
            I => \N__8079\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8119\,
            I => \N__8079\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8118\,
            I => \N__8079\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8117\,
            I => \N__8079\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8116\,
            I => \N__8076\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__8113\,
            I => \N__8070\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__8110\,
            I => \N__8070\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8067\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8106\,
            I => \N__8062\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8105\,
            I => \N__8057\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8104\,
            I => \N__8057\
        );

    \I__1799\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8054\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8100\,
            I => \N__8051\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8048\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8098\,
            I => \N__8043\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8043\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8096\,
            I => \N__8040\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8093\,
            I => \N__8037\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8092\,
            I => \N__8028\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8028\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8090\,
            I => \N__8028\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8028\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__8088\,
            I => \N__8025\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__8079\,
            I => \N__8020\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8076\,
            I => \N__8017\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8075\,
            I => \N__8014\
        );

    \I__1784\ : Span4Mux_v
    port map (
            O => \N__8070\,
            I => \N__8009\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8067\,
            I => \N__8009\
        );

    \I__1782\ : InMux
    port map (
            O => \N__8066\,
            I => \N__8004\
        );

    \I__1781\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8004\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__8062\,
            I => \N__8001\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8057\,
            I => \N__7998\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__8054\,
            I => \N__7991\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__8051\,
            I => \N__7991\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__8048\,
            I => \N__7991\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__8043\,
            I => \N__7988\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__8040\,
            I => \N__7985\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__8037\,
            I => \N__7980\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8028\,
            I => \N__7980\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8025\,
            I => \N__7977\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8024\,
            I => \N__7974\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8023\,
            I => \N__7971\
        );

    \I__1768\ : Span4Mux_h
    port map (
            O => \N__8020\,
            I => \N__7962\
        );

    \I__1767\ : Span4Mux_h
    port map (
            O => \N__8017\,
            I => \N__7962\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__8014\,
            I => \N__7962\
        );

    \I__1765\ : Span4Mux_h
    port map (
            O => \N__8009\,
            I => \N__7962\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8004\,
            I => \N__7953\
        );

    \I__1763\ : Span4Mux_h
    port map (
            O => \N__8001\,
            I => \N__7953\
        );

    \I__1762\ : Span4Mux_h
    port map (
            O => \N__7998\,
            I => \N__7953\
        );

    \I__1761\ : Span4Mux_h
    port map (
            O => \N__7991\,
            I => \N__7953\
        );

    \I__1760\ : Span4Mux_h
    port map (
            O => \N__7988\,
            I => \N__7944\
        );

    \I__1759\ : Span4Mux_h
    port map (
            O => \N__7985\,
            I => \N__7944\
        );

    \I__1758\ : Span4Mux_h
    port map (
            O => \N__7980\,
            I => \N__7944\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__7977\,
            I => \N__7944\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__7974\,
            I => \CPU_CYCLEm\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__7971\,
            I => \CPU_CYCLEm\
        );

    \I__1754\ : Odrv4
    port map (
            O => \N__7962\,
            I => \CPU_CYCLEm\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__7953\,
            I => \CPU_CYCLEm\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__7944\,
            I => \CPU_CYCLEm\
        );

    \I__1751\ : InMux
    port map (
            O => \N__7933\,
            I => \N__7930\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__7930\,
            I => \N__7926\
        );

    \I__1749\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7923\
        );

    \I__1748\ : Sp12to4
    port map (
            O => \N__7926\,
            I => \N__7920\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__7923\,
            I => \N__7917\
        );

    \I__1746\ : Span12Mux_v
    port map (
            O => \N__7920\,
            I => \N__7914\
        );

    \I__1745\ : Span12Mux_v
    port map (
            O => \N__7917\,
            I => \N__7911\
        );

    \I__1744\ : Span12Mux_h
    port map (
            O => \N__7914\,
            I => \N__7908\
        );

    \I__1743\ : Span12Mux_h
    port map (
            O => \N__7911\,
            I => \N__7905\
        );

    \I__1742\ : Odrv12
    port map (
            O => \N__7908\,
            I => \AWEn_c\
        );

    \I__1741\ : Odrv12
    port map (
            O => \N__7905\,
            I => \AWEn_c\
        );

    \I__1740\ : InMux
    port map (
            O => \N__7900\,
            I => \N__7897\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__7897\,
            I => \U712_CHIP_RAM.N_47\
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__7894\,
            I => \N__7891\
        );

    \I__1737\ : InMux
    port map (
            O => \N__7891\,
            I => \N__7888\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__7888\,
            I => \N__7884\
        );

    \I__1735\ : InMux
    port map (
            O => \N__7887\,
            I => \N__7877\
        );

    \I__1734\ : Span4Mux_v
    port map (
            O => \N__7884\,
            I => \N__7874\
        );

    \I__1733\ : InMux
    port map (
            O => \N__7883\,
            I => \N__7867\
        );

    \I__1732\ : InMux
    port map (
            O => \N__7882\,
            I => \N__7867\
        );

    \I__1731\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7867\
        );

    \I__1730\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7864\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__7877\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1728\ : Odrv4
    port map (
            O => \N__7874\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__7867\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__7864\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1725\ : InMux
    port map (
            O => \N__7855\,
            I => \N__7850\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__7854\,
            I => \N__7847\
        );

    \I__1723\ : InMux
    port map (
            O => \N__7853\,
            I => \N__7844\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__7850\,
            I => \N__7841\
        );

    \I__1721\ : InMux
    port map (
            O => \N__7847\,
            I => \N__7836\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__7844\,
            I => \N__7833\
        );

    \I__1719\ : Span4Mux_h
    port map (
            O => \N__7841\,
            I => \N__7830\
        );

    \I__1718\ : InMux
    port map (
            O => \N__7840\,
            I => \N__7825\
        );

    \I__1717\ : InMux
    port map (
            O => \N__7839\,
            I => \N__7825\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__7836\,
            I => \U712_CHIP_RAM.N_63\
        );

    \I__1715\ : Odrv4
    port map (
            O => \N__7833\,
            I => \U712_CHIP_RAM.N_63\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__7830\,
            I => \U712_CHIP_RAM.N_63\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__7825\,
            I => \U712_CHIP_RAM.N_63\
        );

    \I__1712\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7812\
        );

    \I__1711\ : InMux
    port map (
            O => \N__7815\,
            I => \N__7809\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__7812\,
            I => \N__7803\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__7809\,
            I => \N__7803\
        );

    \I__1708\ : InMux
    port map (
            O => \N__7808\,
            I => \N__7800\
        );

    \I__1707\ : Span4Mux_v
    port map (
            O => \N__7803\,
            I => \N__7792\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__7800\,
            I => \N__7789\
        );

    \I__1705\ : InMux
    port map (
            O => \N__7799\,
            I => \N__7784\
        );

    \I__1704\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7784\
        );

    \I__1703\ : InMux
    port map (
            O => \N__7797\,
            I => \N__7781\
        );

    \I__1702\ : InMux
    port map (
            O => \N__7796\,
            I => \N__7777\
        );

    \I__1701\ : InMux
    port map (
            O => \N__7795\,
            I => \N__7774\
        );

    \I__1700\ : Span4Mux_h
    port map (
            O => \N__7792\,
            I => \N__7767\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__7789\,
            I => \N__7767\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__7784\,
            I => \N__7767\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__7781\,
            I => \N__7764\
        );

    \I__1696\ : InMux
    port map (
            O => \N__7780\,
            I => \N__7761\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__7777\,
            I => \N__7758\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__7774\,
            I => \N__7755\
        );

    \I__1693\ : Span4Mux_h
    port map (
            O => \N__7767\,
            I => \N__7747\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__7764\,
            I => \N__7747\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__7761\,
            I => \N__7744\
        );

    \I__1690\ : Span4Mux_v
    port map (
            O => \N__7758\,
            I => \N__7739\
        );

    \I__1689\ : Span4Mux_v
    port map (
            O => \N__7755\,
            I => \N__7739\
        );

    \I__1688\ : InMux
    port map (
            O => \N__7754\,
            I => \N__7734\
        );

    \I__1687\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7734\
        );

    \I__1686\ : InMux
    port map (
            O => \N__7752\,
            I => \N__7731\
        );

    \I__1685\ : Span4Mux_h
    port map (
            O => \N__7747\,
            I => \N__7728\
        );

    \I__1684\ : Span12Mux_v
    port map (
            O => \N__7744\,
            I => \N__7719\
        );

    \I__1683\ : Sp12to4
    port map (
            O => \N__7739\,
            I => \N__7719\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__7734\,
            I => \N__7719\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__7731\,
            I => \N__7719\
        );

    \I__1680\ : Span4Mux_h
    port map (
            O => \N__7728\,
            I => \N__7716\
        );

    \I__1679\ : Span12Mux_h
    port map (
            O => \N__7719\,
            I => \N__7713\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__7716\,
            I => \RESETn_c\
        );

    \I__1677\ : Odrv12
    port map (
            O => \N__7713\,
            I => \RESETn_c\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__7708\,
            I => \N__7703\
        );

    \I__1675\ : InMux
    port map (
            O => \N__7707\,
            I => \N__7696\
        );

    \I__1674\ : InMux
    port map (
            O => \N__7706\,
            I => \N__7696\
        );

    \I__1673\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7693\
        );

    \I__1672\ : InMux
    port map (
            O => \N__7702\,
            I => \N__7688\
        );

    \I__1671\ : InMux
    port map (
            O => \N__7701\,
            I => \N__7688\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__7696\,
            I => \N__7685\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__7693\,
            I => \N__7674\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__7688\,
            I => \N__7669\
        );

    \I__1667\ : Span4Mux_v
    port map (
            O => \N__7685\,
            I => \N__7669\
        );

    \I__1666\ : InMux
    port map (
            O => \N__7684\,
            I => \N__7664\
        );

    \I__1665\ : InMux
    port map (
            O => \N__7683\,
            I => \N__7664\
        );

    \I__1664\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7661\
        );

    \I__1663\ : InMux
    port map (
            O => \N__7681\,
            I => \N__7654\
        );

    \I__1662\ : InMux
    port map (
            O => \N__7680\,
            I => \N__7654\
        );

    \I__1661\ : InMux
    port map (
            O => \N__7679\,
            I => \N__7654\
        );

    \I__1660\ : InMux
    port map (
            O => \N__7678\,
            I => \N__7649\
        );

    \I__1659\ : InMux
    port map (
            O => \N__7677\,
            I => \N__7649\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__7674\,
            I => \N__7646\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__7669\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__7664\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__7661\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__7654\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__7649\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1652\ : Odrv4
    port map (
            O => \N__7646\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1651\ : CascadeMux
    port map (
            O => \N__7633\,
            I => \U712_CHIP_RAM.N_63_cascade_\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__7630\,
            I => \N__7625\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__7629\,
            I => \N__7621\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7628\,
            I => \N__7616\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7625\,
            I => \N__7616\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__7624\,
            I => \N__7612\
        );

    \I__1645\ : InMux
    port map (
            O => \N__7621\,
            I => \N__7606\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7616\,
            I => \N__7603\
        );

    \I__1643\ : InMux
    port map (
            O => \N__7615\,
            I => \N__7600\
        );

    \I__1642\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7597\
        );

    \I__1641\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7592\
        );

    \I__1640\ : InMux
    port map (
            O => \N__7610\,
            I => \N__7592\
        );

    \I__1639\ : InMux
    port map (
            O => \N__7609\,
            I => \N__7589\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__7606\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46\
        );

    \I__1637\ : Odrv12
    port map (
            O => \N__7603\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__7600\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__7597\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__7592\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7589\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER46\
        );

    \I__1632\ : InMux
    port map (
            O => \N__7576\,
            I => \N__7572\
        );

    \I__1631\ : InMux
    port map (
            O => \N__7575\,
            I => \N__7566\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__7572\,
            I => \N__7563\
        );

    \I__1629\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7560\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7557\
        );

    \I__1627\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7554\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__7566\,
            I => \U712_CHIP_RAM.N_127\
        );

    \I__1625\ : Odrv12
    port map (
            O => \N__7563\,
            I => \U712_CHIP_RAM.N_127\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7560\,
            I => \U712_CHIP_RAM.N_127\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7557\,
            I => \U712_CHIP_RAM.N_127\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__7554\,
            I => \U712_CHIP_RAM.N_127\
        );

    \I__1621\ : InMux
    port map (
            O => \N__7543\,
            I => \N__7537\
        );

    \I__1620\ : InMux
    port map (
            O => \N__7542\,
            I => \N__7537\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7537\,
            I => \N__7534\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__7534\,
            I => \N__7531\
        );

    \I__1617\ : Odrv4
    port map (
            O => \N__7531\,
            I => \U712_CHIP_RAM.N_124\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__7528\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_cascade_\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__7525\,
            I => \N__7518\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__7524\,
            I => \N__7515\
        );

    \I__1613\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7510\
        );

    \I__1612\ : InMux
    port map (
            O => \N__7522\,
            I => \N__7507\
        );

    \I__1611\ : InMux
    port map (
            O => \N__7521\,
            I => \N__7502\
        );

    \I__1610\ : InMux
    port map (
            O => \N__7518\,
            I => \N__7502\
        );

    \I__1609\ : InMux
    port map (
            O => \N__7515\,
            I => \N__7499\
        );

    \I__1608\ : InMux
    port map (
            O => \N__7514\,
            I => \N__7494\
        );

    \I__1607\ : InMux
    port map (
            O => \N__7513\,
            I => \N__7494\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__7510\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__7507\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__7502\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__7499\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__7494\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7483\,
            I => \N__7480\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7480\,
            I => \U712_CHIP_RAM.N_107\
        );

    \I__1599\ : IoInMux
    port map (
            O => \N__7477\,
            I => \N__7474\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__7474\,
            I => \N__7471\
        );

    \I__1597\ : Span4Mux_s3_v
    port map (
            O => \N__7471\,
            I => \N__7468\
        );

    \I__1596\ : Span4Mux_h
    port map (
            O => \N__7468\,
            I => \N__7464\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__7467\,
            I => \N__7461\
        );

    \I__1594\ : Sp12to4
    port map (
            O => \N__7464\,
            I => \N__7457\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7461\,
            I => \N__7454\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__7460\,
            I => \N__7451\
        );

    \I__1591\ : Span12Mux_v
    port map (
            O => \N__7457\,
            I => \N__7448\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__7454\,
            I => \N__7445\
        );

    \I__1589\ : InMux
    port map (
            O => \N__7451\,
            I => \N__7442\
        );

    \I__1588\ : Odrv12
    port map (
            O => \N__7448\,
            I => \DBDIR_c\
        );

    \I__1587\ : Odrv12
    port map (
            O => \N__7445\,
            I => \DBDIR_c\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__7442\,
            I => \DBDIR_c\
        );

    \I__1585\ : IoInMux
    port map (
            O => \N__7435\,
            I => \N__7432\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7432\,
            I => \N__7429\
        );

    \I__1583\ : Span4Mux_s1_h
    port map (
            O => \N__7429\,
            I => \N__7426\
        );

    \I__1582\ : Sp12to4
    port map (
            O => \N__7426\,
            I => \N__7423\
        );

    \I__1581\ : Span12Mux_v
    port map (
            O => \N__7423\,
            I => \N__7420\
        );

    \I__1580\ : Span12Mux_h
    port map (
            O => \N__7420\,
            I => \N__7417\
        );

    \I__1579\ : Odrv12
    port map (
            O => \N__7417\,
            I => \DRDDIR_0_i\
        );

    \I__1578\ : IoInMux
    port map (
            O => \N__7414\,
            I => \N__7411\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7411\,
            I => \N__7408\
        );

    \I__1576\ : Span4Mux_s2_v
    port map (
            O => \N__7408\,
            I => \N__7405\
        );

    \I__1575\ : Span4Mux_v
    port map (
            O => \N__7405\,
            I => \N__7402\
        );

    \I__1574\ : Span4Mux_v
    port map (
            O => \N__7402\,
            I => \N__7399\
        );

    \I__1573\ : Odrv4
    port map (
            O => \N__7399\,
            I => \CMA_c_10\
        );

    \I__1572\ : CEMux
    port map (
            O => \N__7396\,
            I => \N__7389\
        );

    \I__1571\ : CEMux
    port map (
            O => \N__7395\,
            I => \N__7386\
        );

    \I__1570\ : CEMux
    port map (
            O => \N__7394\,
            I => \N__7383\
        );

    \I__1569\ : CEMux
    port map (
            O => \N__7393\,
            I => \N__7380\
        );

    \I__1568\ : CEMux
    port map (
            O => \N__7392\,
            I => \N__7376\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__7389\,
            I => \N__7373\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7386\,
            I => \N__7368\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__7383\,
            I => \N__7368\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__7380\,
            I => \N__7365\
        );

    \I__1563\ : CEMux
    port map (
            O => \N__7379\,
            I => \N__7362\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__7376\,
            I => \N__7359\
        );

    \I__1561\ : Span4Mux_h
    port map (
            O => \N__7373\,
            I => \N__7354\
        );

    \I__1560\ : Span4Mux_v
    port map (
            O => \N__7368\,
            I => \N__7354\
        );

    \I__1559\ : Span4Mux_v
    port map (
            O => \N__7365\,
            I => \N__7351\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7362\,
            I => \N__7348\
        );

    \I__1557\ : Span4Mux_h
    port map (
            O => \N__7359\,
            I => \N__7345\
        );

    \I__1556\ : Span4Mux_h
    port map (
            O => \N__7354\,
            I => \N__7342\
        );

    \I__1555\ : Span4Mux_v
    port map (
            O => \N__7351\,
            I => \N__7339\
        );

    \I__1554\ : Odrv12
    port map (
            O => \N__7348\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__7345\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__7342\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__7339\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7330\,
            I => \N__7326\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7329\,
            I => \N__7323\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7326\,
            I => \N__7320\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7323\,
            I => \N__7317\
        );

    \I__1546\ : Span4Mux_v
    port map (
            O => \N__7320\,
            I => \N__7314\
        );

    \I__1545\ : Span12Mux_v
    port map (
            O => \N__7317\,
            I => \N__7309\
        );

    \I__1544\ : Sp12to4
    port map (
            O => \N__7314\,
            I => \N__7309\
        );

    \I__1543\ : Span12Mux_h
    port map (
            O => \N__7309\,
            I => \N__7306\
        );

    \I__1542\ : Odrv12
    port map (
            O => \N__7306\,
            I => \DRA_c_7\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7303\,
            I => \N__7300\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7300\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7297\,
            I => \N__7294\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7294\,
            I => \N__7290\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7293\,
            I => \N__7287\
        );

    \I__1536\ : Span4Mux_v
    port map (
            O => \N__7290\,
            I => \N__7284\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__7287\,
            I => \N__7281\
        );

    \I__1534\ : Sp12to4
    port map (
            O => \N__7284\,
            I => \N__7278\
        );

    \I__1533\ : Span4Mux_v
    port map (
            O => \N__7281\,
            I => \N__7275\
        );

    \I__1532\ : Span12Mux_h
    port map (
            O => \N__7278\,
            I => \N__7272\
        );

    \I__1531\ : Sp12to4
    port map (
            O => \N__7275\,
            I => \N__7269\
        );

    \I__1530\ : Odrv12
    port map (
            O => \N__7272\,
            I => \DRA_c_8\
        );

    \I__1529\ : Odrv12
    port map (
            O => \N__7269\,
            I => \DRA_c_8\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7264\,
            I => \N__7261\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7261\,
            I => \N__7258\
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__7258\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1525\ : InMux
    port map (
            O => \N__7255\,
            I => \N__7252\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7252\,
            I => \N__7248\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7251\,
            I => \N__7245\
        );

    \I__1522\ : Odrv4
    port map (
            O => \N__7248\,
            I => \U712_CHIP_RAM.N_65\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7245\,
            I => \U712_CHIP_RAM.N_65\
        );

    \I__1520\ : InMux
    port map (
            O => \N__7240\,
            I => \N__7237\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7237\,
            I => \N__7232\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7236\,
            I => \N__7229\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7235\,
            I => \N__7226\
        );

    \I__1516\ : Odrv12
    port map (
            O => \N__7232\,
            I => \U712_CHIP_RAM.N_78\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__7229\,
            I => \U712_CHIP_RAM.N_78\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__7226\,
            I => \U712_CHIP_RAM.N_78\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7219\,
            I => \N__7214\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7218\,
            I => \N__7211\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7217\,
            I => \N__7208\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7214\,
            I => \N__7204\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__7211\,
            I => \N__7199\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7208\,
            I => \N__7199\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7207\,
            I => \N__7194\
        );

    \I__1506\ : Span4Mux_h
    port map (
            O => \N__7204\,
            I => \N__7189\
        );

    \I__1505\ : Span4Mux_h
    port map (
            O => \N__7199\,
            I => \N__7186\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7198\,
            I => \N__7181\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7197\,
            I => \N__7181\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7194\,
            I => \N__7178\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7173\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7173\
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__7189\,
            I => \U712_CHIP_RAM.N_67\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__7186\,
            I => \U712_CHIP_RAM.N_67\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7181\,
            I => \U712_CHIP_RAM.N_67\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__7178\,
            I => \U712_CHIP_RAM.N_67\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7173\,
            I => \U712_CHIP_RAM.N_67\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__7162\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_cascade_\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7159\,
            I => \N__7156\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7156\,
            I => \N__7153\
        );

    \I__1491\ : Span4Mux_v
    port map (
            O => \N__7153\,
            I => \N__7150\
        );

    \I__1490\ : Odrv4
    port map (
            O => \N__7150\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7147\,
            I => \N__7144\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7144\,
            I => \N__7141\
        );

    \I__1487\ : Span4Mux_v
    port map (
            O => \N__7141\,
            I => \N__7138\
        );

    \I__1486\ : Odrv4
    port map (
            O => \N__7138\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_5\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7131\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7134\,
            I => \N__7128\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7131\,
            I => \U712_CHIP_RAM.N_77\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7128\,
            I => \U712_CHIP_RAM.N_77\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__7123\,
            I => \U712_CHIP_RAM.N_80_cascade_\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__7120\,
            I => \U712_CHIP_RAM.N_50_cascade_\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7117\,
            I => \N__7113\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7116\,
            I => \N__7108\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__7113\,
            I => \N__7105\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7112\,
            I => \N__7102\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7111\,
            I => \N__7099\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7108\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__7105\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__7102\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7099\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7090\,
            I => \N__7085\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__7089\,
            I => \N__7082\
        );

    \I__1468\ : InMux
    port map (
            O => \N__7088\,
            I => \N__7079\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__7085\,
            I => \N__7076\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7082\,
            I => \N__7073\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7079\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1464\ : Odrv4
    port map (
            O => \N__7076\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7073\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__7066\,
            I => \N__7062\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7065\,
            I => \N__7055\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7062\,
            I => \N__7055\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7061\,
            I => \N__7052\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7060\,
            I => \N__7049\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7055\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7052\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7049\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7042\,
            I => \N__7036\
        );

    \I__1453\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7036\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__7036\,
            I => \U712_CHIP_RAM.N_60\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7033\,
            I => \N__7030\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7030\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER39_0\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__7027\,
            I => \N__7022\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__7026\,
            I => \N__7019\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7025\,
            I => \N__7016\
        );

    \I__1446\ : InMux
    port map (
            O => \N__7022\,
            I => \N__7009\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7019\,
            I => \N__7009\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__7016\,
            I => \N__7006\
        );

    \I__1443\ : InMux
    port map (
            O => \N__7015\,
            I => \N__7003\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7014\,
            I => \N__7000\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7009\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1440\ : Odrv4
    port map (
            O => \N__7006\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__7003\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__7000\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1437\ : InMux
    port map (
            O => \N__6991\,
            I => \N__6985\
        );

    \I__1436\ : InMux
    port map (
            O => \N__6990\,
            I => \N__6985\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__6985\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER39_2\
        );

    \I__1434\ : InMux
    port map (
            O => \N__6982\,
            I => \N__6978\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6981\,
            I => \N__6969\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__6978\,
            I => \N__6966\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__6977\,
            I => \N__6963\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__6976\,
            I => \N__6960\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__6975\,
            I => \N__6951\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__6974\,
            I => \N__6948\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6973\,
            I => \N__6944\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6972\,
            I => \N__6941\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__6969\,
            I => \N__6938\
        );

    \I__1424\ : Span4Mux_h
    port map (
            O => \N__6966\,
            I => \N__6935\
        );

    \I__1423\ : InMux
    port map (
            O => \N__6963\,
            I => \N__6932\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6960\,
            I => \N__6929\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6959\,
            I => \N__6926\
        );

    \I__1420\ : InMux
    port map (
            O => \N__6958\,
            I => \N__6921\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6957\,
            I => \N__6921\
        );

    \I__1418\ : InMux
    port map (
            O => \N__6956\,
            I => \N__6916\
        );

    \I__1417\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6916\
        );

    \I__1416\ : InMux
    port map (
            O => \N__6954\,
            I => \N__6907\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6951\,
            I => \N__6907\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6948\,
            I => \N__6907\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6947\,
            I => \N__6907\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6944\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6941\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1410\ : Odrv12
    port map (
            O => \N__6938\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1409\ : Odrv4
    port map (
            O => \N__6935\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__6932\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__6929\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__6926\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__6921\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__6916\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__6907\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6886\,
            I => \N__6882\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6885\,
            I => \N__6879\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__6882\,
            I => \U712_CHIP_RAM.N_50\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__6879\,
            I => \U712_CHIP_RAM.N_50\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__6874\,
            I => \N__6869\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__6873\,
            I => \N__6865\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__6872\,
            I => \N__6858\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6869\,
            I => \N__6848\
        );

    \I__1394\ : InMux
    port map (
            O => \N__6868\,
            I => \N__6848\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6865\,
            I => \N__6843\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6864\,
            I => \N__6838\
        );

    \I__1391\ : InMux
    port map (
            O => \N__6863\,
            I => \N__6838\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__6862\,
            I => \N__6834\
        );

    \I__1389\ : InMux
    port map (
            O => \N__6861\,
            I => \N__6830\
        );

    \I__1388\ : InMux
    port map (
            O => \N__6858\,
            I => \N__6827\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6857\,
            I => \N__6820\
        );

    \I__1386\ : InMux
    port map (
            O => \N__6856\,
            I => \N__6820\
        );

    \I__1385\ : InMux
    port map (
            O => \N__6855\,
            I => \N__6820\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__6854\,
            I => \N__6817\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__6853\,
            I => \N__6814\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__6848\,
            I => \N__6811\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6847\,
            I => \N__6808\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6801\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6843\,
            I => \N__6796\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6838\,
            I => \N__6796\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6837\,
            I => \N__6791\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6834\,
            I => \N__6791\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6833\,
            I => \N__6788\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__6830\,
            I => \N__6781\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__6827\,
            I => \N__6781\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__6820\,
            I => \N__6781\
        );

    \I__1371\ : InMux
    port map (
            O => \N__6817\,
            I => \N__6776\
        );

    \I__1370\ : InMux
    port map (
            O => \N__6814\,
            I => \N__6776\
        );

    \I__1369\ : Span12Mux_v
    port map (
            O => \N__6811\,
            I => \N__6771\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__6808\,
            I => \N__6771\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6807\,
            I => \N__6762\
        );

    \I__1366\ : InMux
    port map (
            O => \N__6806\,
            I => \N__6762\
        );

    \I__1365\ : InMux
    port map (
            O => \N__6805\,
            I => \N__6762\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6804\,
            I => \N__6762\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__6801\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1362\ : Odrv12
    port map (
            O => \N__6796\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6791\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__6788\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1359\ : Odrv4
    port map (
            O => \N__6781\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__6776\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1357\ : Odrv12
    port map (
            O => \N__6771\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__6762\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6740\
        );

    \I__1354\ : InMux
    port map (
            O => \N__6744\,
            I => \N__6735\
        );

    \I__1353\ : InMux
    port map (
            O => \N__6743\,
            I => \N__6735\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__6740\,
            I => \N__6732\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6735\,
            I => \N__6729\
        );

    \I__1350\ : Span4Mux_v
    port map (
            O => \N__6732\,
            I => \N__6726\
        );

    \I__1349\ : Sp12to4
    port map (
            O => \N__6729\,
            I => \N__6723\
        );

    \I__1348\ : Sp12to4
    port map (
            O => \N__6726\,
            I => \N__6720\
        );

    \I__1347\ : Span12Mux_v
    port map (
            O => \N__6723\,
            I => \N__6717\
        );

    \I__1346\ : Span12Mux_h
    port map (
            O => \N__6720\,
            I => \N__6714\
        );

    \I__1345\ : Span12Mux_h
    port map (
            O => \N__6717\,
            I => \N__6711\
        );

    \I__1344\ : Span12Mux_v
    port map (
            O => \N__6714\,
            I => \N__6708\
        );

    \I__1343\ : Odrv12
    port map (
            O => \N__6711\,
            I => \CASLn_c\
        );

    \I__1342\ : Odrv12
    port map (
            O => \N__6708\,
            I => \CASLn_c\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6703\,
            I => \N__6697\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6702\,
            I => \N__6697\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__6697\,
            I => \N__6693\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6696\,
            I => \N__6690\
        );

    \I__1337\ : Span4Mux_h
    port map (
            O => \N__6693\,
            I => \N__6687\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__6690\,
            I => \N__6684\
        );

    \I__1335\ : Sp12to4
    port map (
            O => \N__6687\,
            I => \N__6679\
        );

    \I__1334\ : Sp12to4
    port map (
            O => \N__6684\,
            I => \N__6679\
        );

    \I__1333\ : Span12Mux_v
    port map (
            O => \N__6679\,
            I => \N__6676\
        );

    \I__1332\ : Span12Mux_h
    port map (
            O => \N__6676\,
            I => \N__6673\
        );

    \I__1331\ : Odrv12
    port map (
            O => \N__6673\,
            I => \CASUn_c\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__6670\,
            I => \N__6666\
        );

    \I__1329\ : InMux
    port map (
            O => \N__6669\,
            I => \N__6662\
        );

    \I__1328\ : InMux
    port map (
            O => \N__6666\,
            I => \N__6657\
        );

    \I__1327\ : InMux
    port map (
            O => \N__6665\,
            I => \N__6657\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__6662\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__6657\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6652\,
            I => \N__6646\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6646\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6646\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6643\,
            I => \N__6640\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6640\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_2_1\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6637\,
            I => \N__6634\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__6634\,
            I => \N__6631\
        );

    \I__1317\ : Odrv4
    port map (
            O => \N__6631\,
            I => \U712_CHIP_RAM.N_108\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__6628\,
            I => \U712_CHIP_RAM.N_77_cascade_\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6625\,
            I => \N__6622\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__6622\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6616\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6616\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_0\
        );

    \I__1311\ : CascadeMux
    port map (
            O => \N__6613\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_\
        );

    \I__1310\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6607\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6607\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__1308\ : CascadeMux
    port map (
            O => \N__6604\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_\
        );

    \I__1307\ : CEMux
    port map (
            O => \N__6601\,
            I => \N__6598\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__6598\,
            I => \N__6595\
        );

    \I__1305\ : Span4Mux_h
    port map (
            O => \N__6595\,
            I => \N__6592\
        );

    \I__1304\ : Span4Mux_h
    port map (
            O => \N__6592\,
            I => \N__6589\
        );

    \I__1303\ : Odrv4
    port map (
            O => \N__6589\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6579\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6585\,
            I => \N__6579\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6584\,
            I => \N__6576\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6579\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6576\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6568\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__6568\,
            I => \U712_CHIP_RAM.N_80\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6565\,
            I => \N__6562\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6562\,
            I => \N__6559\
        );

    \I__1293\ : Odrv12
    port map (
            O => \N__6559\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6553\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__6553\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6546\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6549\,
            I => \N__6543\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6546\,
            I => \N__6540\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__6543\,
            I => \N__6537\
        );

    \I__1286\ : Sp12to4
    port map (
            O => \N__6540\,
            I => \N__6534\
        );

    \I__1285\ : Span12Mux_v
    port map (
            O => \N__6537\,
            I => \N__6531\
        );

    \I__1284\ : Span12Mux_v
    port map (
            O => \N__6534\,
            I => \N__6528\
        );

    \I__1283\ : Span12Mux_h
    port map (
            O => \N__6531\,
            I => \N__6525\
        );

    \I__1282\ : Span12Mux_h
    port map (
            O => \N__6528\,
            I => \N__6522\
        );

    \I__1281\ : Odrv12
    port map (
            O => \N__6525\,
            I => \DRA_c_4\
        );

    \I__1280\ : Odrv12
    port map (
            O => \N__6522\,
            I => \DRA_c_4\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6517\,
            I => \N__6514\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__6514\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__1277\ : InMux
    port map (
            O => \N__6511\,
            I => \N__6508\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__6508\,
            I => \N__6505\
        );

    \I__1275\ : Span4Mux_v
    port map (
            O => \N__6505\,
            I => \N__6501\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6504\,
            I => \N__6498\
        );

    \I__1273\ : Odrv4
    port map (
            O => \N__6501\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_1_a3_0\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6498\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_1_a3_0\
        );

    \I__1271\ : InMux
    port map (
            O => \N__6493\,
            I => \N__6490\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__6490\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6481\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6481\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__6481\,
            I => \N__6478\
        );

    \I__1266\ : Odrv4
    port map (
            O => \N__6478\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6472\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6472\,
            I => \N__6469\
        );

    \I__1263\ : Span4Mux_h
    port map (
            O => \N__6469\,
            I => \N__6466\
        );

    \I__1262\ : Span4Mux_h
    port map (
            O => \N__6466\,
            I => \N__6463\
        );

    \I__1261\ : Odrv4
    port map (
            O => \N__6463\,
            I => \U712_REG_SM.N_173_0\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6460\,
            I => \N__6457\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6457\,
            I => \N__6454\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__6454\,
            I => \N__6451\
        );

    \I__1257\ : Span4Mux_h
    port map (
            O => \N__6451\,
            I => \N__6447\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6450\,
            I => \N__6444\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__6447\,
            I => \U712_REG_SM.N_183_1\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6444\,
            I => \U712_REG_SM.N_183_1\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__6439\,
            I => \N__6436\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6436\,
            I => \N__6433\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__6433\,
            I => \N__6430\
        );

    \I__1250\ : Span4Mux_h
    port map (
            O => \N__6430\,
            I => \N__6427\
        );

    \I__1249\ : Span4Mux_h
    port map (
            O => \N__6427\,
            I => \N__6423\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6426\,
            I => \N__6420\
        );

    \I__1247\ : Odrv4
    port map (
            O => \N__6423\,
            I => \U712_REG_SM.N_165_0\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6420\,
            I => \U712_REG_SM.N_165_0\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6415\,
            I => \N__6412\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6412\,
            I => \N__6408\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6411\,
            I => \N__6405\
        );

    \I__1242\ : Span4Mux_h
    port map (
            O => \N__6408\,
            I => \N__6399\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6405\,
            I => \N__6399\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6404\,
            I => \N__6396\
        );

    \I__1239\ : Span4Mux_h
    port map (
            O => \N__6399\,
            I => \N__6393\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6396\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__6393\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6384\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6387\,
            I => \N__6381\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6384\,
            I => \N__6372\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6381\,
            I => \N__6372\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6380\,
            I => \N__6369\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6379\,
            I => \N__6366\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6378\,
            I => \N__6363\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6377\,
            I => \N__6360\
        );

    \I__1228\ : Span4Mux_h
    port map (
            O => \N__6372\,
            I => \N__6355\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6369\,
            I => \N__6355\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6366\,
            I => \N__6352\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6363\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6360\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__6355\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__6352\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__6343\,
            I => \N__6340\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6340\,
            I => \N__6337\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6337\,
            I => \N__6333\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6330\
        );

    \I__1217\ : Span4Mux_h
    port map (
            O => \N__6333\,
            I => \N__6327\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__6330\,
            I => \U712_CHIP_RAM.un1_DBR_SYNC\
        );

    \I__1215\ : Odrv4
    port map (
            O => \N__6327\,
            I => \U712_CHIP_RAM.un1_DBR_SYNC\
        );

    \I__1214\ : CEMux
    port map (
            O => \N__6322\,
            I => \N__6319\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__6319\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6313\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6313\,
            I => \N__6309\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6306\
        );

    \I__1209\ : Span4Mux_h
    port map (
            O => \N__6309\,
            I => \N__6300\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__6306\,
            I => \N__6300\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6297\
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__6300\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6297\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6292\,
            I => \N__6289\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6289\,
            I => \N__6285\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__6288\,
            I => \N__6282\
        );

    \I__1201\ : Span4Mux_v
    port map (
            O => \N__6285\,
            I => \N__6279\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6282\,
            I => \N__6276\
        );

    \I__1199\ : Odrv4
    port map (
            O => \N__6279\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6276\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__1197\ : IoInMux
    port map (
            O => \N__6271\,
            I => \N__6268\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__6268\,
            I => \N__6265\
        );

    \I__1195\ : IoSpan4Mux
    port map (
            O => \N__6265\,
            I => \N__6262\
        );

    \I__1194\ : Span4Mux_s3_v
    port map (
            O => \N__6262\,
            I => \N__6259\
        );

    \I__1193\ : Sp12to4
    port map (
            O => \N__6259\,
            I => \N__6256\
        );

    \I__1192\ : Span12Mux_s11_v
    port map (
            O => \N__6256\,
            I => \N__6253\
        );

    \I__1191\ : Odrv12
    port map (
            O => \N__6253\,
            I => \U712_REG_SM_un1_LDSn_i\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6250\,
            I => \N__6247\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__6247\,
            I => \N__6244\
        );

    \I__1188\ : Odrv4
    port map (
            O => \N__6244\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6237\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6240\,
            I => \N__6234\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6237\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6234\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__6229\,
            I => \N__6225\
        );

    \I__1182\ : InMux
    port map (
            O => \N__6228\,
            I => \N__6222\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6219\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6222\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6219\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6211\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6211\,
            I => \N__6208\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__6208\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__1175\ : IoInMux
    port map (
            O => \N__6205\,
            I => \N__6202\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6202\,
            I => \N__6199\
        );

    \I__1173\ : IoSpan4Mux
    port map (
            O => \N__6199\,
            I => \N__6196\
        );

    \I__1172\ : IoSpan4Mux
    port map (
            O => \N__6196\,
            I => \N__6193\
        );

    \I__1171\ : Span4Mux_s2_h
    port map (
            O => \N__6193\,
            I => \N__6190\
        );

    \I__1170\ : Sp12to4
    port map (
            O => \N__6190\,
            I => \N__6187\
        );

    \I__1169\ : Odrv12
    port map (
            O => \N__6187\,
            I => \CMA_c_7\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6181\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__6181\,
            I => \N__6178\
        );

    \I__1166\ : Span4Mux_v
    port map (
            O => \N__6178\,
            I => \N__6175\
        );

    \I__1165\ : Span4Mux_v
    port map (
            O => \N__6175\,
            I => \N__6172\
        );

    \I__1164\ : Sp12to4
    port map (
            O => \N__6172\,
            I => \N__6169\
        );

    \I__1163\ : Span12Mux_h
    port map (
            O => \N__6169\,
            I => \N__6166\
        );

    \I__1162\ : Odrv12
    port map (
            O => \N__6166\,
            I => \A_c_18\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__6163\,
            I => \N__6160\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6160\,
            I => \N__6157\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6157\,
            I => \N__6154\
        );

    \I__1158\ : Span4Mux_v
    port map (
            O => \N__6154\,
            I => \N__6151\
        );

    \I__1157\ : Span4Mux_v
    port map (
            O => \N__6151\,
            I => \N__6148\
        );

    \I__1156\ : Sp12to4
    port map (
            O => \N__6148\,
            I => \N__6145\
        );

    \I__1155\ : Span12Mux_h
    port map (
            O => \N__6145\,
            I => \N__6142\
        );

    \I__1154\ : Odrv12
    port map (
            O => \N__6142\,
            I => \A_c_16\
        );

    \I__1153\ : InMux
    port map (
            O => \N__6139\,
            I => \N__6136\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6136\,
            I => \U712_CHIP_RAM.N_39\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6130\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6130\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_7\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__6127\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_0_cascade_\
        );

    \I__1148\ : CEMux
    port map (
            O => \N__6124\,
            I => \N__6120\
        );

    \I__1147\ : CEMux
    port map (
            O => \N__6123\,
            I => \N__6117\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6120\,
            I => \N__6114\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6117\,
            I => \N__6111\
        );

    \I__1144\ : Odrv4
    port map (
            O => \N__6114\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_i\
        );

    \I__1143\ : Odrv4
    port map (
            O => \N__6111\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_i\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__6106\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_5_cascade_\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6103\,
            I => \N__6100\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__6100\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER18_0\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__6097\,
            I => \N__6094\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6091\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6091\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6085\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6085\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_4\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6078\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6075\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6078\,
            I => \U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6075\,
            I => \U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6070\,
            I => \N__6066\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6069\,
            I => \N__6063\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6066\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER18_0\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__6063\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER18_0\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__6058\,
            I => \U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa_cascade_\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__6055\,
            I => \N__6050\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__6054\,
            I => \N__6046\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6053\,
            I => \N__6043\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6050\,
            I => \N__6040\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6037\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6046\,
            I => \N__6034\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6043\,
            I => \U712_CHIP_RAM.N_158_0\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6040\,
            I => \U712_CHIP_RAM.N_158_0\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__6037\,
            I => \U712_CHIP_RAM.N_158_0\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6034\,
            I => \U712_CHIP_RAM.N_158_0\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6025\,
            I => \N__6022\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6022\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_ns_1_1\
        );

    \I__1113\ : CascadeMux
    port map (
            O => \N__6019\,
            I => \N__6016\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6016\,
            I => \N__6013\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__6013\,
            I => \U712_CHIP_RAM.N_132\
        );

    \I__1110\ : SRMux
    port map (
            O => \N__6010\,
            I => \N__6007\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6007\,
            I => \N__6004\
        );

    \I__1108\ : Odrv4
    port map (
            O => \N__6004\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5998\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__5998\,
            I => \N__5995\
        );

    \I__1105\ : Odrv12
    port map (
            O => \N__5995\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1104\ : InMux
    port map (
            O => \N__5992\,
            I => \N__5989\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5989\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1102\ : InMux
    port map (
            O => \N__5986\,
            I => \N__5983\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5983\,
            I => \N__5980\
        );

    \I__1100\ : Span4Mux_v
    port map (
            O => \N__5980\,
            I => \N__5977\
        );

    \I__1099\ : Sp12to4
    port map (
            O => \N__5977\,
            I => \N__5974\
        );

    \I__1098\ : Span12Mux_h
    port map (
            O => \N__5974\,
            I => \N__5971\
        );

    \I__1097\ : Span12Mux_v
    port map (
            O => \N__5971\,
            I => \N__5968\
        );

    \I__1096\ : Odrv12
    port map (
            O => \N__5968\,
            I => \A_c_17\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__5965\,
            I => \U712_CHIP_RAM.CMA_5_0_8_cascade_\
        );

    \I__1094\ : IoInMux
    port map (
            O => \N__5962\,
            I => \N__5959\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5959\,
            I => \N__5956\
        );

    \I__1092\ : IoSpan4Mux
    port map (
            O => \N__5956\,
            I => \N__5953\
        );

    \I__1091\ : Span4Mux_s3_h
    port map (
            O => \N__5953\,
            I => \N__5950\
        );

    \I__1090\ : Sp12to4
    port map (
            O => \N__5950\,
            I => \N__5947\
        );

    \I__1089\ : Span12Mux_h
    port map (
            O => \N__5947\,
            I => \N__5944\
        );

    \I__1088\ : Odrv12
    port map (
            O => \N__5944\,
            I => \CMA_c_8\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5938\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5938\,
            I => \N__5935\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__5935\,
            I => \U712_CHIP_RAM.N_38\
        );

    \I__1084\ : IoInMux
    port map (
            O => \N__5932\,
            I => \N__5929\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__5929\,
            I => \N__5926\
        );

    \I__1082\ : Span4Mux_s2_h
    port map (
            O => \N__5926\,
            I => \N__5923\
        );

    \I__1081\ : Sp12to4
    port map (
            O => \N__5923\,
            I => \N__5920\
        );

    \I__1080\ : Span12Mux_s6_v
    port map (
            O => \N__5920\,
            I => \N__5917\
        );

    \I__1079\ : Span12Mux_h
    port map (
            O => \N__5917\,
            I => \N__5914\
        );

    \I__1078\ : Odrv12
    port map (
            O => \N__5914\,
            I => \CMA_c_6\
        );

    \I__1077\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5908\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5908\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__5905\,
            I => \N__5902\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5899\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__5899\,
            I => \N__5896\
        );

    \I__1072\ : Span4Mux_h
    port map (
            O => \N__5896\,
            I => \N__5893\
        );

    \I__1071\ : Sp12to4
    port map (
            O => \N__5893\,
            I => \N__5890\
        );

    \I__1070\ : Span12Mux_v
    port map (
            O => \N__5890\,
            I => \N__5887\
        );

    \I__1069\ : Span12Mux_h
    port map (
            O => \N__5887\,
            I => \N__5884\
        );

    \I__1068\ : Odrv12
    port map (
            O => \N__5884\,
            I => \A_c_19\
        );

    \I__1067\ : IoInMux
    port map (
            O => \N__5881\,
            I => \N__5878\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5878\,
            I => \N__5875\
        );

    \I__1065\ : Span4Mux_s3_h
    port map (
            O => \N__5875\,
            I => \N__5872\
        );

    \I__1064\ : Span4Mux_v
    port map (
            O => \N__5872\,
            I => \N__5869\
        );

    \I__1063\ : Span4Mux_v
    port map (
            O => \N__5869\,
            I => \N__5866\
        );

    \I__1062\ : Sp12to4
    port map (
            O => \N__5866\,
            I => \N__5863\
        );

    \I__1061\ : Odrv12
    port map (
            O => \N__5863\,
            I => \CMA_c_9\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5857\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5857\,
            I => \N__5853\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5856\,
            I => \N__5850\
        );

    \I__1057\ : Span12Mux_v
    port map (
            O => \N__5853\,
            I => \N__5847\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__5850\,
            I => \N__5844\
        );

    \I__1055\ : Span12Mux_v
    port map (
            O => \N__5847\,
            I => \N__5841\
        );

    \I__1054\ : Span12Mux_h
    port map (
            O => \N__5844\,
            I => \N__5838\
        );

    \I__1053\ : Span12Mux_h
    port map (
            O => \N__5841\,
            I => \N__5835\
        );

    \I__1052\ : Span12Mux_v
    port map (
            O => \N__5838\,
            I => \N__5832\
        );

    \I__1051\ : Odrv12
    port map (
            O => \N__5835\,
            I => \DRA_c_1\
        );

    \I__1050\ : Odrv12
    port map (
            O => \N__5832\,
            I => \DRA_c_1\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5827\,
            I => \N__5824\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5824\,
            I => \N__5821\
        );

    \I__1047\ : Odrv4
    port map (
            O => \N__5821\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5815\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5815\,
            I => \N__5811\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5814\,
            I => \N__5808\
        );

    \I__1043\ : Sp12to4
    port map (
            O => \N__5811\,
            I => \N__5803\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5808\,
            I => \N__5803\
        );

    \I__1041\ : Span12Mux_v
    port map (
            O => \N__5803\,
            I => \N__5800\
        );

    \I__1040\ : Span12Mux_h
    port map (
            O => \N__5800\,
            I => \N__5797\
        );

    \I__1039\ : Odrv12
    port map (
            O => \N__5797\,
            I => \DRA_c_6\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5794\,
            I => \N__5791\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__5791\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1036\ : IoInMux
    port map (
            O => \N__5788\,
            I => \N__5785\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5785\,
            I => \N__5782\
        );

    \I__1034\ : Span4Mux_s0_v
    port map (
            O => \N__5782\,
            I => \N__5779\
        );

    \I__1033\ : Sp12to4
    port map (
            O => \N__5779\,
            I => \N__5776\
        );

    \I__1032\ : Span12Mux_h
    port map (
            O => \N__5776\,
            I => \N__5773\
        );

    \I__1031\ : Span12Mux_v
    port map (
            O => \N__5773\,
            I => \N__5765\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5756\
        );

    \I__1029\ : InMux
    port map (
            O => \N__5771\,
            I => \N__5756\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5770\,
            I => \N__5756\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5769\,
            I => \N__5756\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5768\,
            I => \N__5753\
        );

    \I__1025\ : Odrv12
    port map (
            O => \N__5765\,
            I => \DBENn_c\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__5756\,
            I => \DBENn_c\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__5753\,
            I => \DBENn_c\
        );

    \I__1022\ : IoInMux
    port map (
            O => \N__5746\,
            I => \N__5743\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__5743\,
            I => \N__5740\
        );

    \I__1020\ : Span4Mux_s3_h
    port map (
            O => \N__5740\,
            I => \N__5737\
        );

    \I__1019\ : Sp12to4
    port map (
            O => \N__5737\,
            I => \N__5734\
        );

    \I__1018\ : Span12Mux_v
    port map (
            O => \N__5734\,
            I => \N__5731\
        );

    \I__1017\ : Span12Mux_h
    port map (
            O => \N__5731\,
            I => \N__5728\
        );

    \I__1016\ : Odrv12
    port map (
            O => \N__5728\,
            I => \CUUBEn_c\
        );

    \I__1015\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5721\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5718\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__5721\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5718\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5713\,
            I => \bfn_14_4_0_\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5710\,
            I => \N__5706\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5709\,
            I => \N__5703\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5706\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__5703\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5698\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5695\,
            I => \N__5691\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5694\,
            I => \N__5688\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5691\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__5688\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5683\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5680\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__5677\,
            I => \N__5673\
        );

    \I__998\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5670\
        );

    \I__997\ : InMux
    port map (
            O => \N__5673\,
            I => \N__5667\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5670\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5667\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__994\ : InMux
    port map (
            O => \N__5662\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__993\ : InMux
    port map (
            O => \N__5659\,
            I => \N__5655\
        );

    \I__992\ : InMux
    port map (
            O => \N__5658\,
            I => \N__5652\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5655\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__5652\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__989\ : InMux
    port map (
            O => \N__5647\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__988\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5640\
        );

    \I__987\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5637\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5640\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__5637\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__984\ : InMux
    port map (
            O => \N__5632\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__983\ : InMux
    port map (
            O => \N__5629\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__982\ : ClkMux
    port map (
            O => \N__5626\,
            I => \N__5623\
        );

    \I__981\ : GlobalMux
    port map (
            O => \N__5623\,
            I => \N__5620\
        );

    \I__980\ : gio2CtrlBuf
    port map (
            O => \N__5620\,
            I => \C1_c_g\
        );

    \I__979\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5613\
        );

    \I__978\ : InMux
    port map (
            O => \N__5616\,
            I => \N__5610\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5613\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5610\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0\
        );

    \I__975\ : InMux
    port map (
            O => \N__5605\,
            I => \N__5602\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__5602\,
            I => \N__5599\
        );

    \I__973\ : Span4Mux_h
    port map (
            O => \N__5599\,
            I => \N__5596\
        );

    \I__972\ : Odrv4
    port map (
            O => \N__5596\,
            I => \U712_CHIP_RAM.DMA_CYCLE_7\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__5593\,
            I => \U712_BYTE_ENABLE.un2_CUMBEnZ0_cascade_\
        );

    \I__970\ : IoInMux
    port map (
            O => \N__5590\,
            I => \N__5587\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__5587\,
            I => \N__5584\
        );

    \I__968\ : Span4Mux_s3_h
    port map (
            O => \N__5584\,
            I => \N__5581\
        );

    \I__967\ : Span4Mux_v
    port map (
            O => \N__5581\,
            I => \N__5578\
        );

    \I__966\ : Sp12to4
    port map (
            O => \N__5578\,
            I => \N__5575\
        );

    \I__965\ : Span12Mux_h
    port map (
            O => \N__5575\,
            I => \N__5572\
        );

    \I__964\ : Span12Mux_v
    port map (
            O => \N__5572\,
            I => \N__5569\
        );

    \I__963\ : Odrv12
    port map (
            O => \N__5569\,
            I => \CUMBEn_c\
        );

    \I__962\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5560\
        );

    \I__961\ : InMux
    port map (
            O => \N__5565\,
            I => \N__5560\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__5560\,
            I => \U712_BYTE_ENABLE.LLBE_0_0_tz\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__5557\,
            I => \U712_BYTE_ENABLE.un2_CLLBEnZ0_cascade_\
        );

    \I__958\ : IoInMux
    port map (
            O => \N__5554\,
            I => \N__5551\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__5551\,
            I => \N__5548\
        );

    \I__956\ : IoSpan4Mux
    port map (
            O => \N__5548\,
            I => \N__5545\
        );

    \I__955\ : Sp12to4
    port map (
            O => \N__5545\,
            I => \N__5542\
        );

    \I__954\ : Span12Mux_s7_v
    port map (
            O => \N__5542\,
            I => \N__5539\
        );

    \I__953\ : Span12Mux_v
    port map (
            O => \N__5539\,
            I => \N__5536\
        );

    \I__952\ : Odrv12
    port map (
            O => \N__5536\,
            I => \CLLBEn_c\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__5533\,
            I => \U712_BYTE_ENABLE.un2_CLMBEnZ0_cascade_\
        );

    \I__950\ : IoInMux
    port map (
            O => \N__5530\,
            I => \N__5527\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5527\,
            I => \N__5524\
        );

    \I__948\ : Span4Mux_s3_h
    port map (
            O => \N__5524\,
            I => \N__5521\
        );

    \I__947\ : Sp12to4
    port map (
            O => \N__5521\,
            I => \N__5518\
        );

    \I__946\ : Span12Mux_v
    port map (
            O => \N__5518\,
            I => \N__5515\
        );

    \I__945\ : Span12Mux_h
    port map (
            O => \N__5515\,
            I => \N__5512\
        );

    \I__944\ : Odrv12
    port map (
            O => \N__5512\,
            I => \CLMBEn_c\
        );

    \I__943\ : InMux
    port map (
            O => \N__5509\,
            I => \N__5497\
        );

    \I__942\ : InMux
    port map (
            O => \N__5508\,
            I => \N__5497\
        );

    \I__941\ : InMux
    port map (
            O => \N__5507\,
            I => \N__5497\
        );

    \I__940\ : InMux
    port map (
            O => \N__5506\,
            I => \N__5497\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5497\,
            I => \N__5494\
        );

    \I__938\ : Span4Mux_v
    port map (
            O => \N__5494\,
            I => \N__5491\
        );

    \I__937\ : Span4Mux_v
    port map (
            O => \N__5491\,
            I => \N__5488\
        );

    \I__936\ : Sp12to4
    port map (
            O => \N__5488\,
            I => \N__5485\
        );

    \I__935\ : Span12Mux_h
    port map (
            O => \N__5485\,
            I => \N__5482\
        );

    \I__934\ : Odrv12
    port map (
            O => \N__5482\,
            I => \A_c_1\
        );

    \I__933\ : InMux
    port map (
            O => \N__5479\,
            I => \N__5470\
        );

    \I__932\ : InMux
    port map (
            O => \N__5478\,
            I => \N__5470\
        );

    \I__931\ : InMux
    port map (
            O => \N__5477\,
            I => \N__5467\
        );

    \I__930\ : InMux
    port map (
            O => \N__5476\,
            I => \N__5462\
        );

    \I__929\ : InMux
    port map (
            O => \N__5475\,
            I => \N__5462\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5470\,
            I => \N__5457\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__5467\,
            I => \N__5457\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5462\,
            I => \N__5454\
        );

    \I__925\ : Span4Mux_v
    port map (
            O => \N__5457\,
            I => \N__5451\
        );

    \I__924\ : Span4Mux_v
    port map (
            O => \N__5454\,
            I => \N__5448\
        );

    \I__923\ : Sp12to4
    port map (
            O => \N__5451\,
            I => \N__5443\
        );

    \I__922\ : Sp12to4
    port map (
            O => \N__5448\,
            I => \N__5443\
        );

    \I__921\ : Span12Mux_h
    port map (
            O => \N__5443\,
            I => \N__5440\
        );

    \I__920\ : Odrv12
    port map (
            O => \N__5440\,
            I => \A_c_0\
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__5437\,
            I => \N__5431\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__5436\,
            I => \N__5428\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__5435\,
            I => \N__5425\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__5434\,
            I => \N__5422\
        );

    \I__915\ : InMux
    port map (
            O => \N__5431\,
            I => \N__5413\
        );

    \I__914\ : InMux
    port map (
            O => \N__5428\,
            I => \N__5413\
        );

    \I__913\ : InMux
    port map (
            O => \N__5425\,
            I => \N__5413\
        );

    \I__912\ : InMux
    port map (
            O => \N__5422\,
            I => \N__5413\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__5413\,
            I => \N__5410\
        );

    \I__910\ : Odrv4
    port map (
            O => \N__5410\,
            I => \U712_BYTE_ENABLE.LW_TRANS_0\
        );

    \I__909\ : CascadeMux
    port map (
            O => \N__5407\,
            I => \U712_BYTE_ENABLE.un2_CUUBEnZ0_cascade_\
        );

    \I__908\ : InMux
    port map (
            O => \N__5404\,
            I => \N__5398\
        );

    \I__907\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5398\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5398\,
            I => \N__5395\
        );

    \I__905\ : Odrv4
    port map (
            O => \N__5395\,
            I => \U712_CHIP_RAM.N_51\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__5392\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER16_2_0_cascade_\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__5389\,
            I => \U712_CHIP_RAM.N_99_cascade_\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__5386\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_cascade_\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__5383\,
            I => \U712_CHIP_RAM.N_67_cascade_\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__5380\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER18_0_cascade_\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__5377\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_m2_3_cascade_\
        );

    \I__898\ : InMux
    port map (
            O => \N__5374\,
            I => \N__5371\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5371\,
            I => \U712_CHIP_RAM.N_35\
        );

    \I__896\ : IoInMux
    port map (
            O => \N__5368\,
            I => \N__5365\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__5365\,
            I => \N__5362\
        );

    \I__894\ : Span4Mux_s3_h
    port map (
            O => \N__5362\,
            I => \N__5359\
        );

    \I__893\ : Sp12to4
    port map (
            O => \N__5359\,
            I => \N__5356\
        );

    \I__892\ : Span12Mux_s6_v
    port map (
            O => \N__5356\,
            I => \N__5353\
        );

    \I__891\ : Span12Mux_h
    port map (
            O => \N__5353\,
            I => \N__5350\
        );

    \I__890\ : Odrv12
    port map (
            O => \N__5350\,
            I => \CMA_c_3\
        );

    \I__889\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5344\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5344\,
            I => \N__5341\
        );

    \I__887\ : Span4Mux_v
    port map (
            O => \N__5341\,
            I => \N__5338\
        );

    \I__886\ : Sp12to4
    port map (
            O => \N__5338\,
            I => \N__5335\
        );

    \I__885\ : Span12Mux_h
    port map (
            O => \N__5335\,
            I => \N__5332\
        );

    \I__884\ : Odrv12
    port map (
            O => \N__5332\,
            I => \A_c_6\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__5329\,
            I => \N__5326\
        );

    \I__882\ : InMux
    port map (
            O => \N__5326\,
            I => \N__5323\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5323\,
            I => \N__5320\
        );

    \I__880\ : Span4Mux_v
    port map (
            O => \N__5320\,
            I => \N__5317\
        );

    \I__879\ : Span4Mux_v
    port map (
            O => \N__5317\,
            I => \N__5314\
        );

    \I__878\ : Sp12to4
    port map (
            O => \N__5314\,
            I => \N__5311\
        );

    \I__877\ : Span12Mux_h
    port map (
            O => \N__5311\,
            I => \N__5308\
        );

    \I__876\ : Odrv12
    port map (
            O => \N__5308\,
            I => \A_c_13\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__5305\,
            I => \U712_CHIP_RAM.N_36_cascade_\
        );

    \I__874\ : IoInMux
    port map (
            O => \N__5302\,
            I => \N__5299\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5299\,
            I => \N__5296\
        );

    \I__872\ : IoSpan4Mux
    port map (
            O => \N__5296\,
            I => \N__5293\
        );

    \I__871\ : Sp12to4
    port map (
            O => \N__5293\,
            I => \N__5290\
        );

    \I__870\ : Span12Mux_s9_v
    port map (
            O => \N__5290\,
            I => \N__5287\
        );

    \I__869\ : Span12Mux_h
    port map (
            O => \N__5287\,
            I => \N__5284\
        );

    \I__868\ : Odrv12
    port map (
            O => \N__5284\,
            I => \CMA_c_4\
        );

    \I__867\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5278\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5278\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_ns_1_2\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__5275\,
            I => \U712_CHIP_RAM.N_61_cascade_\
        );

    \I__864\ : CascadeMux
    port map (
            O => \N__5272\,
            I => \U712_CHIP_RAM.N_65_cascade_\
        );

    \I__863\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5266\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__5266\,
            I => \U712_CHIP_RAM.N_104_1\
        );

    \I__861\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5260\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__5260\,
            I => \N__5257\
        );

    \I__859\ : Span4Mux_v
    port map (
            O => \N__5257\,
            I => \N__5254\
        );

    \I__858\ : Sp12to4
    port map (
            O => \N__5254\,
            I => \N__5251\
        );

    \I__857\ : Span12Mux_h
    port map (
            O => \N__5251\,
            I => \N__5248\
        );

    \I__856\ : Odrv12
    port map (
            O => \N__5248\,
            I => \A_c_9\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__5245\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_\
        );

    \I__854\ : InMux
    port map (
            O => \N__5242\,
            I => \N__5239\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5239\,
            I => \N__5236\
        );

    \I__852\ : Span4Mux_v
    port map (
            O => \N__5236\,
            I => \N__5233\
        );

    \I__851\ : Sp12to4
    port map (
            O => \N__5233\,
            I => \N__5230\
        );

    \I__850\ : Span12Mux_h
    port map (
            O => \N__5230\,
            I => \N__5227\
        );

    \I__849\ : Span12Mux_v
    port map (
            O => \N__5227\,
            I => \N__5224\
        );

    \I__848\ : Odrv12
    port map (
            O => \N__5224\,
            I => \A_c_2\
        );

    \I__847\ : InMux
    port map (
            O => \N__5221\,
            I => \N__5218\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5218\,
            I => \U712_CHIP_RAM.N_32\
        );

    \I__845\ : InMux
    port map (
            O => \N__5215\,
            I => \N__5212\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5212\,
            I => \N__5209\
        );

    \I__843\ : Odrv4
    port map (
            O => \N__5209\,
            I => \U712_CHIP_RAM.N_37\
        );

    \I__842\ : IoInMux
    port map (
            O => \N__5206\,
            I => \N__5203\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5203\,
            I => \N__5200\
        );

    \I__840\ : Span4Mux_s3_h
    port map (
            O => \N__5200\,
            I => \N__5197\
        );

    \I__839\ : Span4Mux_v
    port map (
            O => \N__5197\,
            I => \N__5194\
        );

    \I__838\ : Sp12to4
    port map (
            O => \N__5194\,
            I => \N__5191\
        );

    \I__837\ : Span12Mux_h
    port map (
            O => \N__5191\,
            I => \N__5188\
        );

    \I__836\ : Odrv12
    port map (
            O => \N__5188\,
            I => \CMA_c_5\
        );

    \I__835\ : InMux
    port map (
            O => \N__5185\,
            I => \N__5181\
        );

    \I__834\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5178\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__5181\,
            I => \N__5173\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5178\,
            I => \N__5173\
        );

    \I__831\ : Span4Mux_v
    port map (
            O => \N__5173\,
            I => \N__5170\
        );

    \I__830\ : Span4Mux_v
    port map (
            O => \N__5170\,
            I => \N__5167\
        );

    \I__829\ : Sp12to4
    port map (
            O => \N__5167\,
            I => \N__5164\
        );

    \I__828\ : Span12Mux_h
    port map (
            O => \N__5164\,
            I => \N__5161\
        );

    \I__827\ : Odrv12
    port map (
            O => \N__5161\,
            I => \DRA_c_3\
        );

    \I__826\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5155\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5155\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__824\ : InMux
    port map (
            O => \N__5152\,
            I => \N__5149\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__5149\,
            I => \N__5145\
        );

    \I__822\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5142\
        );

    \I__821\ : Span4Mux_v
    port map (
            O => \N__5145\,
            I => \N__5139\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5142\,
            I => \N__5136\
        );

    \I__819\ : Sp12to4
    port map (
            O => \N__5139\,
            I => \N__5133\
        );

    \I__818\ : Sp12to4
    port map (
            O => \N__5136\,
            I => \N__5130\
        );

    \I__817\ : Span12Mux_h
    port map (
            O => \N__5133\,
            I => \N__5127\
        );

    \I__816\ : Span12Mux_v
    port map (
            O => \N__5130\,
            I => \N__5124\
        );

    \I__815\ : Span12Mux_v
    port map (
            O => \N__5127\,
            I => \N__5121\
        );

    \I__814\ : Span12Mux_h
    port map (
            O => \N__5124\,
            I => \N__5118\
        );

    \I__813\ : Odrv12
    port map (
            O => \N__5121\,
            I => \DRA_c_2\
        );

    \I__812\ : Odrv12
    port map (
            O => \N__5118\,
            I => \DRA_c_2\
        );

    \I__811\ : InMux
    port map (
            O => \N__5113\,
            I => \N__5110\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__5110\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__809\ : InMux
    port map (
            O => \N__5107\,
            I => \N__5104\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5104\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__807\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5098\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5098\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__805\ : InMux
    port map (
            O => \N__5095\,
            I => \N__5092\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5092\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_5\
        );

    \I__803\ : InMux
    port map (
            O => \N__5089\,
            I => \N__5085\
        );

    \I__802\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5082\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5085\,
            I => \N__5077\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__5082\,
            I => \N__5077\
        );

    \I__799\ : Span4Mux_v
    port map (
            O => \N__5077\,
            I => \N__5074\
        );

    \I__798\ : Span4Mux_v
    port map (
            O => \N__5074\,
            I => \N__5071\
        );

    \I__797\ : Sp12to4
    port map (
            O => \N__5071\,
            I => \N__5068\
        );

    \I__796\ : Span12Mux_h
    port map (
            O => \N__5068\,
            I => \N__5065\
        );

    \I__795\ : Odrv12
    port map (
            O => \N__5065\,
            I => \DRA_c_5\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__5062\,
            I => \N__5059\
        );

    \I__793\ : InMux
    port map (
            O => \N__5059\,
            I => \N__5056\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5056\,
            I => \N__5052\
        );

    \I__791\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5049\
        );

    \I__790\ : Odrv4
    port map (
            O => \N__5052\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5049\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__788\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5040\
        );

    \I__787\ : CascadeMux
    port map (
            O => \N__5043\,
            I => \N__5033\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5040\,
            I => \N__5030\
        );

    \I__785\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5027\
        );

    \I__784\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5024\
        );

    \I__783\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5017\
        );

    \I__782\ : InMux
    port map (
            O => \N__5036\,
            I => \N__5017\
        );

    \I__781\ : InMux
    port map (
            O => \N__5033\,
            I => \N__5017\
        );

    \I__780\ : Span4Mux_h
    port map (
            O => \N__5030\,
            I => \N__5014\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5027\,
            I => \N__5007\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5024\,
            I => \N__5007\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5017\,
            I => \N__5007\
        );

    \I__776\ : Odrv4
    port map (
            O => \N__5014\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__775\ : Odrv12
    port map (
            O => \N__5007\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__5002\,
            I => \N__4999\
        );

    \I__773\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4996\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__4996\,
            I => \N__4993\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__4993\,
            I => \U712_REG_SM.RnW_m\
        );

    \I__770\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4987\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4987\,
            I => \U712_REG_SM.un1_LDS_OUT_0_sqmuxa_1_0\
        );

    \I__768\ : InMux
    port map (
            O => \N__4984\,
            I => \N__4981\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4981\,
            I => \N__4978\
        );

    \I__766\ : Span12Mux_h
    port map (
            O => \N__4978\,
            I => \N__4975\
        );

    \I__765\ : Span12Mux_v
    port map (
            O => \N__4975\,
            I => \N__4972\
        );

    \I__764\ : Odrv12
    port map (
            O => \N__4972\,
            I => \DBRn_c\
        );

    \I__763\ : InMux
    port map (
            O => \N__4969\,
            I => \N__4965\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__4968\,
            I => \N__4962\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4965\,
            I => \N__4959\
        );

    \I__760\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4956\
        );

    \I__759\ : Span4Mux_v
    port map (
            O => \N__4959\,
            I => \N__4952\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4956\,
            I => \N__4949\
        );

    \I__757\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4945\
        );

    \I__756\ : Sp12to4
    port map (
            O => \N__4952\,
            I => \N__4940\
        );

    \I__755\ : Span12Mux_v
    port map (
            O => \N__4949\,
            I => \N__4940\
        );

    \I__754\ : InMux
    port map (
            O => \N__4948\,
            I => \N__4937\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4945\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__752\ : Odrv12
    port map (
            O => \N__4940\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4937\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__750\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4926\
        );

    \I__749\ : InMux
    port map (
            O => \N__4929\,
            I => \N__4923\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4926\,
            I => \N__4918\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__4923\,
            I => \N__4918\
        );

    \I__746\ : Span4Mux_h
    port map (
            O => \N__4918\,
            I => \N__4914\
        );

    \I__745\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4911\
        );

    \I__744\ : Odrv4
    port map (
            O => \N__4914\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__4911\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__742\ : InMux
    port map (
            O => \N__4906\,
            I => \N__4903\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4903\,
            I => \N__4899\
        );

    \I__740\ : InMux
    port map (
            O => \N__4902\,
            I => \N__4896\
        );

    \I__739\ : Span4Mux_v
    port map (
            O => \N__4899\,
            I => \N__4893\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4896\,
            I => \N__4890\
        );

    \I__737\ : Span4Mux_h
    port map (
            O => \N__4893\,
            I => \N__4887\
        );

    \I__736\ : Span4Mux_v
    port map (
            O => \N__4890\,
            I => \N__4884\
        );

    \I__735\ : Sp12to4
    port map (
            O => \N__4887\,
            I => \N__4879\
        );

    \I__734\ : Sp12to4
    port map (
            O => \N__4884\,
            I => \N__4879\
        );

    \I__733\ : Span12Mux_h
    port map (
            O => \N__4879\,
            I => \N__4876\
        );

    \I__732\ : Span12Mux_v
    port map (
            O => \N__4876\,
            I => \N__4873\
        );

    \I__731\ : Odrv12
    port map (
            O => \N__4873\,
            I => \SIZ_c_1\
        );

    \I__730\ : InMux
    port map (
            O => \N__4870\,
            I => \N__4866\
        );

    \I__729\ : CascadeMux
    port map (
            O => \N__4869\,
            I => \N__4863\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4866\,
            I => \N__4860\
        );

    \I__727\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4857\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__4860\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4857\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__724\ : IoInMux
    port map (
            O => \N__4852\,
            I => \N__4849\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__4849\,
            I => \N__4846\
        );

    \I__722\ : Span4Mux_s3_v
    port map (
            O => \N__4846\,
            I => \N__4843\
        );

    \I__721\ : Span4Mux_v
    port map (
            O => \N__4843\,
            I => \N__4840\
        );

    \I__720\ : Span4Mux_v
    port map (
            O => \N__4840\,
            I => \N__4837\
        );

    \I__719\ : Sp12to4
    port map (
            O => \N__4837\,
            I => \N__4834\
        );

    \I__718\ : Odrv12
    port map (
            O => \N__4834\,
            I => \U712_REG_SM_un1_UDSn_i\
        );

    \I__717\ : IoInMux
    port map (
            O => \N__4831\,
            I => \N__4828\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4828\,
            I => \N__4825\
        );

    \I__715\ : Odrv12
    port map (
            O => \N__4825\,
            I => \RESETn_c_i\
        );

    \I__714\ : InMux
    port map (
            O => \N__4822\,
            I => \N__4819\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__4819\,
            I => \N__4816\
        );

    \I__712\ : Span12Mux_v
    port map (
            O => \N__4816\,
            I => \N__4813\
        );

    \I__711\ : Span12Mux_h
    port map (
            O => \N__4813\,
            I => \N__4810\
        );

    \I__710\ : Odrv12
    port map (
            O => \N__4810\,
            I => \A_c_15\
        );

    \I__709\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4804\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4804\,
            I => \N__4801\
        );

    \I__707\ : Span4Mux_v
    port map (
            O => \N__4801\,
            I => \N__4798\
        );

    \I__706\ : Sp12to4
    port map (
            O => \N__4798\,
            I => \N__4795\
        );

    \I__705\ : Span12Mux_h
    port map (
            O => \N__4795\,
            I => \N__4792\
        );

    \I__704\ : Odrv12
    port map (
            O => \N__4792\,
            I => \A_c_8\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__4789\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_6_cascade_\
        );

    \I__702\ : InMux
    port map (
            O => \N__4786\,
            I => \N__4783\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__4783\,
            I => \N__4780\
        );

    \I__700\ : Span12Mux_v
    port map (
            O => \N__4780\,
            I => \N__4777\
        );

    \I__699\ : Span12Mux_h
    port map (
            O => \N__4777\,
            I => \N__4774\
        );

    \I__698\ : Odrv12
    port map (
            O => \N__4774\,
            I => \A_c_5\
        );

    \I__697\ : CascadeMux
    port map (
            O => \N__4771\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_\
        );

    \I__696\ : InMux
    port map (
            O => \N__4768\,
            I => \N__4765\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4765\,
            I => \N__4762\
        );

    \I__694\ : Span4Mux_v
    port map (
            O => \N__4762\,
            I => \N__4759\
        );

    \I__693\ : Sp12to4
    port map (
            O => \N__4759\,
            I => \N__4756\
        );

    \I__692\ : Span12Mux_h
    port map (
            O => \N__4756\,
            I => \N__4753\
        );

    \I__691\ : Odrv12
    port map (
            O => \N__4753\,
            I => \A_c_12\
        );

    \I__690\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4747\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__4747\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__688\ : InMux
    port map (
            O => \N__4744\,
            I => \N__4741\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__4741\,
            I => \N__4738\
        );

    \I__686\ : Odrv4
    port map (
            O => \N__4738\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__685\ : InMux
    port map (
            O => \N__4735\,
            I => \N__4730\
        );

    \I__684\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4727\
        );

    \I__683\ : InMux
    port map (
            O => \N__4733\,
            I => \N__4724\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__4730\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4727\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__4724\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__679\ : InMux
    port map (
            O => \N__4717\,
            I => \N__4714\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__4714\,
            I => \N__4709\
        );

    \I__677\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4706\
        );

    \I__676\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4703\
        );

    \I__675\ : Odrv4
    port map (
            O => \N__4709\,
            I => \U712_REG_SM.N_167_0\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__4706\,
            I => \U712_REG_SM.N_167_0\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4703\,
            I => \U712_REG_SM.N_167_0\
        );

    \I__672\ : InMux
    port map (
            O => \N__4696\,
            I => \N__4693\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4693\,
            I => \N__4690\
        );

    \I__670\ : Span4Mux_h
    port map (
            O => \N__4690\,
            I => \N__4687\
        );

    \I__669\ : Odrv4
    port map (
            O => \N__4687\,
            I => \U712_REG_SM.N_117\
        );

    \I__668\ : InMux
    port map (
            O => \N__4684\,
            I => \N__4681\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__4681\,
            I => \N__4677\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__4680\,
            I => \N__4673\
        );

    \I__665\ : Span4Mux_v
    port map (
            O => \N__4677\,
            I => \N__4670\
        );

    \I__664\ : InMux
    port map (
            O => \N__4676\,
            I => \N__4667\
        );

    \I__663\ : InMux
    port map (
            O => \N__4673\,
            I => \N__4664\
        );

    \I__662\ : Sp12to4
    port map (
            O => \N__4670\,
            I => \N__4659\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4667\,
            I => \N__4659\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4664\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__659\ : Odrv12
    port map (
            O => \N__4659\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__658\ : InMux
    port map (
            O => \N__4654\,
            I => \N__4647\
        );

    \I__657\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4647\
        );

    \I__656\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4644\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__4647\,
            I => \N__4639\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4644\,
            I => \N__4639\
        );

    \I__653\ : Sp12to4
    port map (
            O => \N__4639\,
            I => \N__4636\
        );

    \I__652\ : Span12Mux_v
    port map (
            O => \N__4636\,
            I => \N__4633\
        );

    \I__651\ : Span12Mux_h
    port map (
            O => \N__4633\,
            I => \N__4630\
        );

    \I__650\ : Odrv12
    port map (
            O => \N__4630\,
            I => \SIZ_c_0\
        );

    \I__649\ : InMux
    port map (
            O => \N__4627\,
            I => \N__4624\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4624\,
            I => \U712_REG_SM.LDS_OUT_2_0_0\
        );

    \I__647\ : InMux
    port map (
            O => \N__4621\,
            I => \N__4618\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__4618\,
            I => \U712_REG_SM.UDS_OUT_2_0_0\
        );

    \I__645\ : IoInMux
    port map (
            O => \N__4615\,
            I => \N__4612\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4612\,
            I => \N__4609\
        );

    \I__643\ : Span12Mux_s0_v
    port map (
            O => \N__4609\,
            I => \N__4606\
        );

    \I__642\ : Span12Mux_v
    port map (
            O => \N__4606\,
            I => \N__4603\
        );

    \I__641\ : Odrv12
    port map (
            O => \N__4603\,
            I => \CMA_c_0\
        );

    \I__640\ : InMux
    port map (
            O => \N__4600\,
            I => \N__4597\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4597\,
            I => \U712_CHIP_RAM.N_33\
        );

    \I__638\ : IoInMux
    port map (
            O => \N__4594\,
            I => \N__4591\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4591\,
            I => \N__4588\
        );

    \I__636\ : Span12Mux_s11_v
    port map (
            O => \N__4588\,
            I => \N__4585\
        );

    \I__635\ : Odrv12
    port map (
            O => \N__4585\,
            I => \CMA_c_1\
        );

    \I__634\ : IoInMux
    port map (
            O => \N__4582\,
            I => \N__4579\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4579\,
            I => \N__4576\
        );

    \I__632\ : IoSpan4Mux
    port map (
            O => \N__4576\,
            I => \N__4573\
        );

    \I__631\ : Sp12to4
    port map (
            O => \N__4573\,
            I => \N__4570\
        );

    \I__630\ : Span12Mux_s7_v
    port map (
            O => \N__4570\,
            I => \N__4567\
        );

    \I__629\ : Odrv12
    port map (
            O => \N__4567\,
            I => \CMA_c_2\
        );

    \I__628\ : InMux
    port map (
            O => \N__4564\,
            I => \N__4561\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__4561\,
            I => \N__4558\
        );

    \I__626\ : Span4Mux_v
    port map (
            O => \N__4558\,
            I => \N__4555\
        );

    \I__625\ : Span4Mux_v
    port map (
            O => \N__4555\,
            I => \N__4552\
        );

    \I__624\ : Sp12to4
    port map (
            O => \N__4552\,
            I => \N__4549\
        );

    \I__623\ : Span12Mux_h
    port map (
            O => \N__4549\,
            I => \N__4546\
        );

    \I__622\ : Odrv12
    port map (
            O => \N__4546\,
            I => \A_c_4\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__4543\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_\
        );

    \I__620\ : InMux
    port map (
            O => \N__4540\,
            I => \N__4537\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4537\,
            I => \N__4534\
        );

    \I__618\ : Span12Mux_v
    port map (
            O => \N__4534\,
            I => \N__4531\
        );

    \I__617\ : Span12Mux_h
    port map (
            O => \N__4531\,
            I => \N__4528\
        );

    \I__616\ : Odrv12
    port map (
            O => \N__4528\,
            I => \A_c_11\
        );

    \I__615\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4522\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__4522\,
            I => \U712_CHIP_RAM.N_34\
        );

    \I__613\ : InMux
    port map (
            O => \N__4519\,
            I => \N__4516\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4516\,
            I => \N__4513\
        );

    \I__611\ : Span4Mux_h
    port map (
            O => \N__4513\,
            I => \N__4510\
        );

    \I__610\ : Span4Mux_v
    port map (
            O => \N__4510\,
            I => \N__4507\
        );

    \I__609\ : Sp12to4
    port map (
            O => \N__4507\,
            I => \N__4504\
        );

    \I__608\ : Odrv12
    port map (
            O => \N__4504\,
            I => \A_c_7\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__4501\,
            I => \N__4498\
        );

    \I__606\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4495\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4495\,
            I => \N__4492\
        );

    \I__604\ : Span4Mux_v
    port map (
            O => \N__4492\,
            I => \N__4489\
        );

    \I__603\ : Span4Mux_v
    port map (
            O => \N__4489\,
            I => \N__4486\
        );

    \I__602\ : Sp12to4
    port map (
            O => \N__4486\,
            I => \N__4483\
        );

    \I__601\ : Span12Mux_h
    port map (
            O => \N__4483\,
            I => \N__4480\
        );

    \I__600\ : Odrv12
    port map (
            O => \N__4480\,
            I => \A_c_14\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__4477\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa_1_cascade_\
        );

    \I__598\ : InMux
    port map (
            O => \N__4474\,
            I => \N__4471\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4471\,
            I => \N__4467\
        );

    \I__596\ : InMux
    port map (
            O => \N__4470\,
            I => \N__4464\
        );

    \I__595\ : Odrv4
    port map (
            O => \N__4467\,
            I => \U712_REG_SM.N_68\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__4464\,
            I => \U712_REG_SM.N_68\
        );

    \I__593\ : CascadeMux
    port map (
            O => \N__4459\,
            I => \U712_REG_SM.N_188_cascade_\
        );

    \I__592\ : InMux
    port map (
            O => \N__4456\,
            I => \N__4451\
        );

    \I__591\ : InMux
    port map (
            O => \N__4455\,
            I => \N__4446\
        );

    \I__590\ : InMux
    port map (
            O => \N__4454\,
            I => \N__4446\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4451\,
            I => \U712_REG_SM.N_162_0\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4446\,
            I => \U712_REG_SM.N_162_0\
        );

    \I__587\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4437\
        );

    \I__586\ : InMux
    port map (
            O => \N__4440\,
            I => \N__4434\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__4437\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4434\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__583\ : IoInMux
    port map (
            O => \N__4429\,
            I => \N__4425\
        );

    \I__582\ : IoInMux
    port map (
            O => \N__4428\,
            I => \N__4422\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__4425\,
            I => \N__4419\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4422\,
            I => \N__4416\
        );

    \I__579\ : IoSpan4Mux
    port map (
            O => \N__4419\,
            I => \N__4413\
        );

    \I__578\ : IoSpan4Mux
    port map (
            O => \N__4416\,
            I => \N__4410\
        );

    \I__577\ : Span4Mux_s1_v
    port map (
            O => \N__4413\,
            I => \N__4407\
        );

    \I__576\ : Span4Mux_s1_v
    port map (
            O => \N__4410\,
            I => \N__4404\
        );

    \I__575\ : Sp12to4
    port map (
            O => \N__4407\,
            I => \N__4401\
        );

    \I__574\ : Sp12to4
    port map (
            O => \N__4404\,
            I => \N__4398\
        );

    \I__573\ : Span12Mux_v
    port map (
            O => \N__4401\,
            I => \N__4394\
        );

    \I__572\ : Span12Mux_v
    port map (
            O => \N__4398\,
            I => \N__4391\
        );

    \I__571\ : InMux
    port map (
            O => \N__4397\,
            I => \N__4388\
        );

    \I__570\ : Odrv12
    port map (
            O => \N__4394\,
            I => \ASn_c\
        );

    \I__569\ : Odrv12
    port map (
            O => \N__4391\,
            I => \ASn_c\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4388\,
            I => \ASn_c\
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__4381\,
            I => \N__4378\
        );

    \I__566\ : InMux
    port map (
            O => \N__4378\,
            I => \N__4372\
        );

    \I__565\ : InMux
    port map (
            O => \N__4377\,
            I => \N__4372\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4372\,
            I => \N__4369\
        );

    \I__563\ : Span4Mux_v
    port map (
            O => \N__4369\,
            I => \N__4366\
        );

    \I__562\ : Span4Mux_v
    port map (
            O => \N__4366\,
            I => \N__4363\
        );

    \I__561\ : Sp12to4
    port map (
            O => \N__4363\,
            I => \N__4360\
        );

    \I__560\ : Span12Mux_h
    port map (
            O => \N__4360\,
            I => \N__4357\
        );

    \I__559\ : Odrv12
    port map (
            O => \N__4357\,
            I => \REGSPACEn_c\
        );

    \I__558\ : InMux
    port map (
            O => \N__4354\,
            I => \N__4348\
        );

    \I__557\ : InMux
    port map (
            O => \N__4353\,
            I => \N__4348\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4348\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa_1\
        );

    \I__555\ : InMux
    port map (
            O => \N__4345\,
            I => \N__4336\
        );

    \I__554\ : InMux
    port map (
            O => \N__4344\,
            I => \N__4336\
        );

    \I__553\ : InMux
    port map (
            O => \N__4343\,
            I => \N__4336\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__4336\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__4333\,
            I => \N__4329\
        );

    \I__550\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4326\
        );

    \I__549\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4323\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4326\,
            I => \N__4320\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4323\,
            I => \N__4317\
        );

    \I__546\ : Span4Mux_v
    port map (
            O => \N__4320\,
            I => \N__4311\
        );

    \I__545\ : Span4Mux_v
    port map (
            O => \N__4317\,
            I => \N__4311\
        );

    \I__544\ : InMux
    port map (
            O => \N__4316\,
            I => \N__4308\
        );

    \I__543\ : Sp12to4
    port map (
            O => \N__4311\,
            I => \N__4303\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4308\,
            I => \N__4303\
        );

    \I__541\ : Span12Mux_h
    port map (
            O => \N__4303\,
            I => \N__4300\
        );

    \I__540\ : Span12Mux_v
    port map (
            O => \N__4300\,
            I => \N__4297\
        );

    \I__539\ : Odrv12
    port map (
            O => \N__4297\,
            I => \TSn_c\
        );

    \I__538\ : InMux
    port map (
            O => \N__4294\,
            I => \N__4291\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__4291\,
            I => \N__4287\
        );

    \I__536\ : IoInMux
    port map (
            O => \N__4290\,
            I => \N__4284\
        );

    \I__535\ : Span12Mux_h
    port map (
            O => \N__4287\,
            I => \N__4281\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__4284\,
            I => \N__4278\
        );

    \I__533\ : Span12Mux_v
    port map (
            O => \N__4281\,
            I => \N__4275\
        );

    \I__532\ : IoSpan4Mux
    port map (
            O => \N__4278\,
            I => \N__4272\
        );

    \I__531\ : Odrv12
    port map (
            O => \N__4275\,
            I => \RAMENn_c\
        );

    \I__530\ : Odrv4
    port map (
            O => \N__4272\,
            I => \RAMENn_c\
        );

    \I__529\ : InMux
    port map (
            O => \N__4267\,
            I => \N__4258\
        );

    \I__528\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4258\
        );

    \I__527\ : InMux
    port map (
            O => \N__4265\,
            I => \N__4253\
        );

    \I__526\ : InMux
    port map (
            O => \N__4264\,
            I => \N__4253\
        );

    \I__525\ : InMux
    port map (
            O => \N__4263\,
            I => \N__4250\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4258\,
            I => \U712_REG_SM.N_171_0\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4253\,
            I => \U712_REG_SM.N_171_0\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4250\,
            I => \U712_REG_SM.N_171_0\
        );

    \I__521\ : InMux
    port map (
            O => \N__4243\,
            I => \N__4236\
        );

    \I__520\ : InMux
    port map (
            O => \N__4242\,
            I => \N__4229\
        );

    \I__519\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4229\
        );

    \I__518\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4229\
        );

    \I__517\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4226\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4236\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4229\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__4226\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__4219\,
            I => \U712_REG_SM.N_165_0_cascade_\
        );

    \I__512\ : InMux
    port map (
            O => \N__4216\,
            I => \N__4210\
        );

    \I__511\ : InMux
    port map (
            O => \N__4215\,
            I => \N__4205\
        );

    \I__510\ : InMux
    port map (
            O => \N__4214\,
            I => \N__4205\
        );

    \I__509\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4202\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4210\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__4205\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4202\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__505\ : InMux
    port map (
            O => \N__4195\,
            I => \N__4192\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__4192\,
            I => \U712_CHIP_RAM.CPU_TACK_6\
        );

    \I__503\ : CascadeMux
    port map (
            O => \N__4189\,
            I => \N__4185\
        );

    \I__502\ : InMux
    port map (
            O => \N__4188\,
            I => \N__4179\
        );

    \I__501\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4179\
        );

    \I__500\ : InMux
    port map (
            O => \N__4184\,
            I => \N__4176\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4179\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4176\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__497\ : InMux
    port map (
            O => \N__4171\,
            I => \N__4167\
        );

    \I__496\ : InMux
    port map (
            O => \N__4170\,
            I => \N__4164\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4167\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4164\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__493\ : InMux
    port map (
            O => \N__4159\,
            I => \N__4156\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__4156\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\
        );

    \I__491\ : InMux
    port map (
            O => \N__4153\,
            I => \N__4150\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4150\,
            I => \N__4147\
        );

    \I__489\ : Span12Mux_h
    port map (
            O => \N__4147\,
            I => \N__4144\
        );

    \I__488\ : Span12Mux_v
    port map (
            O => \N__4144\,
            I => \N__4141\
        );

    \I__487\ : Odrv12
    port map (
            O => \N__4141\,
            I => \A_c_3\
        );

    \I__486\ : CascadeMux
    port map (
            O => \N__4138\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\
        );

    \I__485\ : InMux
    port map (
            O => \N__4135\,
            I => \N__4132\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4132\,
            I => \N__4129\
        );

    \I__483\ : Span4Mux_v
    port map (
            O => \N__4129\,
            I => \N__4126\
        );

    \I__482\ : Sp12to4
    port map (
            O => \N__4126\,
            I => \N__4123\
        );

    \I__481\ : Span12Mux_h
    port map (
            O => \N__4123\,
            I => \N__4120\
        );

    \I__480\ : Odrv12
    port map (
            O => \N__4120\,
            I => \A_c_10\
        );

    \I__479\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4114\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4114\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__477\ : InMux
    port map (
            O => \N__4111\,
            I => \N__4108\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4108\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_a3_0\
        );

    \I__475\ : CascadeMux
    port map (
            O => \N__4105\,
            I => \N__4102\
        );

    \I__474\ : InMux
    port map (
            O => \N__4102\,
            I => \N__4098\
        );

    \I__473\ : InMux
    port map (
            O => \N__4101\,
            I => \N__4095\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4098\,
            I => \CPU_TACKm\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4095\,
            I => \CPU_TACKm\
        );

    \I__470\ : CascadeMux
    port map (
            O => \N__4090\,
            I => \N__4087\
        );

    \I__469\ : InMux
    port map (
            O => \N__4087\,
            I => \N__4084\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4084\,
            I => \N__4079\
        );

    \I__467\ : InMux
    port map (
            O => \N__4083\,
            I => \N__4074\
        );

    \I__466\ : InMux
    port map (
            O => \N__4082\,
            I => \N__4074\
        );

    \I__465\ : Odrv12
    port map (
            O => \N__4079\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4074\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__463\ : CascadeMux
    port map (
            O => \N__4069\,
            I => \U712_REG_SM.N_173_0_cascade_\
        );

    \I__462\ : InMux
    port map (
            O => \N__4066\,
            I => \N__4061\
        );

    \I__461\ : InMux
    port map (
            O => \N__4065\,
            I => \N__4056\
        );

    \I__460\ : InMux
    port map (
            O => \N__4064\,
            I => \N__4056\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__4061\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4056\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__4051\,
            I => \U712_REG_SM.N_54_cascade_\
        );

    \I__456\ : InMux
    port map (
            O => \N__4048\,
            I => \N__4045\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4045\,
            I => \U712_REG_SM.un1_STATE_COUNT_5_0_1\
        );

    \I__454\ : InMux
    port map (
            O => \N__4042\,
            I => \N__4038\
        );

    \I__453\ : InMux
    port map (
            O => \N__4041\,
            I => \N__4035\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4038\,
            I => \REG_TACK\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__4035\,
            I => \REG_TACK\
        );

    \I__450\ : CascadeMux
    port map (
            O => \N__4030\,
            I => \U712_REG_SM.N_162_0_cascade_\
        );

    \I__449\ : InMux
    port map (
            O => \N__4027\,
            I => \N__4024\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4024\,
            I => \N__4014\
        );

    \I__447\ : InMux
    port map (
            O => \N__4023\,
            I => \N__4009\
        );

    \I__446\ : InMux
    port map (
            O => \N__4022\,
            I => \N__4009\
        );

    \I__445\ : InMux
    port map (
            O => \N__4021\,
            I => \N__4006\
        );

    \I__444\ : InMux
    port map (
            O => \N__4020\,
            I => \N__3999\
        );

    \I__443\ : InMux
    port map (
            O => \N__4019\,
            I => \N__3999\
        );

    \I__442\ : InMux
    port map (
            O => \N__4018\,
            I => \N__3999\
        );

    \I__441\ : InMux
    port map (
            O => \N__4017\,
            I => \N__3996\
        );

    \I__440\ : Span4Mux_v
    port map (
            O => \N__4014\,
            I => \N__3993\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4009\,
            I => \N__3986\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__4006\,
            I => \N__3986\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__3999\,
            I => \N__3986\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3996\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__435\ : Odrv4
    port map (
            O => \N__3993\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__434\ : Odrv4
    port map (
            O => \N__3986\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__433\ : InMux
    port map (
            O => \N__3979\,
            I => \N__3971\
        );

    \I__432\ : InMux
    port map (
            O => \N__3978\,
            I => \N__3971\
        );

    \I__431\ : InMux
    port map (
            O => \N__3977\,
            I => \N__3968\
        );

    \I__430\ : InMux
    port map (
            O => \N__3976\,
            I => \N__3965\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3971\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3968\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3965\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__3958\,
            I => \N__3953\
        );

    \I__425\ : InMux
    port map (
            O => \N__3957\,
            I => \N__3948\
        );

    \I__424\ : InMux
    port map (
            O => \N__3956\,
            I => \N__3943\
        );

    \I__423\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3943\
        );

    \I__422\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3940\
        );

    \I__421\ : InMux
    port map (
            O => \N__3951\,
            I => \N__3937\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3948\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3943\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3940\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3937\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__416\ : InMux
    port map (
            O => \N__3928\,
            I => \N__3925\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3925\,
            I => \N__3919\
        );

    \I__414\ : InMux
    port map (
            O => \N__3924\,
            I => \N__3912\
        );

    \I__413\ : InMux
    port map (
            O => \N__3923\,
            I => \N__3912\
        );

    \I__412\ : InMux
    port map (
            O => \N__3922\,
            I => \N__3912\
        );

    \I__411\ : Span4Mux_v
    port map (
            O => \N__3919\,
            I => \N__3909\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3912\,
            I => \N__3906\
        );

    \I__409\ : Span4Mux_v
    port map (
            O => \N__3909\,
            I => \N__3903\
        );

    \I__408\ : Span4Mux_h
    port map (
            O => \N__3906\,
            I => \N__3900\
        );

    \I__407\ : Sp12to4
    port map (
            O => \N__3903\,
            I => \N__3897\
        );

    \I__406\ : Sp12to4
    port map (
            O => \N__3900\,
            I => \N__3894\
        );

    \I__405\ : Span12Mux_h
    port map (
            O => \N__3897\,
            I => \N__3889\
        );

    \I__404\ : Span12Mux_v
    port map (
            O => \N__3894\,
            I => \N__3889\
        );

    \I__403\ : Odrv12
    port map (
            O => \N__3889\,
            I => \CLK40_OUT_i\
        );

    \I__402\ : InMux
    port map (
            O => \N__3886\,
            I => \N__3874\
        );

    \I__401\ : InMux
    port map (
            O => \N__3885\,
            I => \N__3874\
        );

    \I__400\ : InMux
    port map (
            O => \N__3884\,
            I => \N__3874\
        );

    \I__399\ : InMux
    port map (
            O => \N__3883\,
            I => \N__3874\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3874\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__397\ : InMux
    port map (
            O => \N__3871\,
            I => \N__3866\
        );

    \I__396\ : InMux
    port map (
            O => \N__3870\,
            I => \N__3863\
        );

    \I__395\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3860\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3866\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3863\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__3860\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__391\ : CascadeMux
    port map (
            O => \N__3853\,
            I => \N__3849\
        );

    \I__390\ : CascadeMux
    port map (
            O => \N__3852\,
            I => \N__3846\
        );

    \I__389\ : InMux
    port map (
            O => \N__3849\,
            I => \N__3843\
        );

    \I__388\ : InMux
    port map (
            O => \N__3846\,
            I => \N__3840\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__3843\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__3840\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__385\ : CascadeMux
    port map (
            O => \N__3835\,
            I => \N__3829\
        );

    \I__384\ : InMux
    port map (
            O => \N__3834\,
            I => \N__3826\
        );

    \I__383\ : InMux
    port map (
            O => \N__3833\,
            I => \N__3823\
        );

    \I__382\ : InMux
    port map (
            O => \N__3832\,
            I => \N__3818\
        );

    \I__381\ : InMux
    port map (
            O => \N__3829\,
            I => \N__3818\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__3826\,
            I => \N__3813\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__3823\,
            I => \N__3813\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3818\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__377\ : Odrv4
    port map (
            O => \N__3813\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__376\ : CascadeMux
    port map (
            O => \N__3808\,
            I => \U712_CYCLE_TERM.N_45_0_0_en_cascade_\
        );

    \I__375\ : CEMux
    port map (
            O => \N__3805\,
            I => \N__3802\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3802\,
            I => \U712_CYCLE_TERM.N_45_0_0_en_0\
        );

    \I__373\ : IoInMux
    port map (
            O => \N__3799\,
            I => \N__3796\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3796\,
            I => \N__3793\
        );

    \I__371\ : IoSpan4Mux
    port map (
            O => \N__3793\,
            I => \N__3790\
        );

    \I__370\ : Span4Mux_s3_v
    port map (
            O => \N__3790\,
            I => \N__3787\
        );

    \I__369\ : Sp12to4
    port map (
            O => \N__3787\,
            I => \N__3784\
        );

    \I__368\ : Odrv12
    port map (
            O => \N__3784\,
            I => \VBENn_c\
        );

    \I__367\ : CascadeMux
    port map (
            O => \N__3781\,
            I => \N__3777\
        );

    \I__366\ : CascadeMux
    port map (
            O => \N__3780\,
            I => \N__3774\
        );

    \I__365\ : InMux
    port map (
            O => \N__3777\,
            I => \N__3770\
        );

    \I__364\ : InMux
    port map (
            O => \N__3774\,
            I => \N__3767\
        );

    \I__363\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3764\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__3770\,
            I => \U712_REG_SM.N_73\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__3767\,
            I => \U712_REG_SM.N_73\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3764\,
            I => \U712_REG_SM.N_73\
        );

    \I__359\ : CascadeMux
    port map (
            O => \N__3757\,
            I => \U712_REG_SM.un1_STATE_COUNT_5_0_1_cascade_\
        );

    \I__358\ : InMux
    port map (
            O => \N__3754\,
            I => \N__3750\
        );

    \I__357\ : InMux
    port map (
            O => \N__3753\,
            I => \N__3747\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__3750\,
            I => \U712_REG_SM.N_86\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__3747\,
            I => \U712_REG_SM.N_86\
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__3742\,
            I => \U712_REG_SM.N_68_cascade_\
        );

    \I__353\ : CascadeMux
    port map (
            O => \N__3739\,
            I => \U712_REG_SM.N_73_cascade_\
        );

    \I__352\ : IoInMux
    port map (
            O => \N__3736\,
            I => \N__3733\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__3733\,
            I => \N__3730\
        );

    \I__350\ : IoSpan4Mux
    port map (
            O => \N__3730\,
            I => \N__3727\
        );

    \I__349\ : Sp12to4
    port map (
            O => \N__3727\,
            I => \N__3724\
        );

    \I__348\ : Span12Mux_h
    port map (
            O => \N__3724\,
            I => \N__3720\
        );

    \I__347\ : InMux
    port map (
            O => \N__3723\,
            I => \N__3717\
        );

    \I__346\ : Odrv12
    port map (
            O => \N__3720\,
            I => \TACK_OUTn\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__3717\,
            I => \TACK_OUTn\
        );

    \I__344\ : IoInMux
    port map (
            O => \N__3712\,
            I => \N__3708\
        );

    \I__343\ : InMux
    port map (
            O => \N__3711\,
            I => \N__3705\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3708\,
            I => \N__3702\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__3705\,
            I => \N__3699\
        );

    \I__340\ : Span4Mux_s3_h
    port map (
            O => \N__3702\,
            I => \N__3696\
        );

    \I__339\ : Span12Mux_h
    port map (
            O => \N__3699\,
            I => \N__3691\
        );

    \I__338\ : Sp12to4
    port map (
            O => \N__3696\,
            I => \N__3691\
        );

    \I__337\ : Span12Mux_v
    port map (
            O => \N__3691\,
            I => \N__3688\
        );

    \I__336\ : Odrv12
    port map (
            O => \N__3688\,
            I => \C1_c\
        );

    \I__335\ : IoInMux
    port map (
            O => \N__3685\,
            I => \N__3682\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__3682\,
            I => \N__3679\
        );

    \I__333\ : Span12Mux_s8_h
    port map (
            O => \N__3679\,
            I => \N__3676\
        );

    \I__332\ : Odrv12
    port map (
            O => \N__3676\,
            I => \CLK40_OUT_i_i\
        );

    \I__331\ : InMux
    port map (
            O => \N__3673\,
            I => \N__3670\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__3670\,
            I => \U712_REG_SM.N_120\
        );

    \I__329\ : InMux
    port map (
            O => \N__3667\,
            I => \N__3664\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__3664\,
            I => \N__3661\
        );

    \I__327\ : Span4Mux_v
    port map (
            O => \N__3661\,
            I => \N__3658\
        );

    \I__326\ : Sp12to4
    port map (
            O => \N__3658\,
            I => \N__3655\
        );

    \I__325\ : Span12Mux_h
    port map (
            O => \N__3655\,
            I => \N__3652\
        );

    \I__324\ : Odrv12
    port map (
            O => \N__3652\,
            I => \C3_c\
        );

    \I__323\ : IoInMux
    port map (
            O => \N__3649\,
            I => \N__3646\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__3646\,
            I => \N__3643\
        );

    \I__321\ : Span4Mux_s2_h
    port map (
            O => \N__3643\,
            I => \N__3640\
        );

    \I__320\ : Sp12to4
    port map (
            O => \N__3640\,
            I => \N__3637\
        );

    \I__319\ : Span12Mux_s11_v
    port map (
            O => \N__3637\,
            I => \N__3634\
        );

    \I__318\ : Odrv12
    port map (
            O => \N__3634\,
            I => \N_677_i\
        );

    \I__317\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3628\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__3628\,
            I => \TACK_EN_i_ess\
        );

    \I__315\ : IoInMux
    port map (
            O => \N__3625\,
            I => \N__3622\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__3622\,
            I => \N__3619\
        );

    \I__313\ : Span4Mux_s2_v
    port map (
            O => \N__3619\,
            I => \N__3616\
        );

    \I__312\ : Span4Mux_v
    port map (
            O => \N__3616\,
            I => \N__3613\
        );

    \I__311\ : Odrv4
    port map (
            O => \N__3613\,
            I => \CLK80_OUT_i_i\
        );

    \I__310\ : IoInMux
    port map (
            O => \N__3610\,
            I => \N__3607\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__3607\,
            I => \N__3604\
        );

    \I__308\ : Span4Mux_s0_v
    port map (
            O => \N__3604\,
            I => \N__3601\
        );

    \I__307\ : Span4Mux_v
    port map (
            O => \N__3601\,
            I => \N__3598\
        );

    \I__306\ : Sp12to4
    port map (
            O => \N__3598\,
            I => \N__3595\
        );

    \I__305\ : Span12Mux_h
    port map (
            O => \N__3595\,
            I => \N__3592\
        );

    \I__304\ : Span12Mux_v
    port map (
            O => \N__3592\,
            I => \N__3589\
        );

    \I__303\ : Odrv12
    port map (
            O => \N__3589\,
            I => \CLK40_IN_c\
        );

    \IN_MUX_bfv_14_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_4_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4831\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3712\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9577\,
            lcout => \CLK80_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK40C_obuf_RNO_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3928\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__4684\,
            in1 => \N__9158\,
            in2 => \N__4090\,
            in3 => \N__3673\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9569\,
            ce => 'H',
            sr => \N__9366\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4027\,
            in2 => \_gnd_net_\,
            in3 => \N__3753\,
            lcout => \U712_REG_SM.N_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3667\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9570\,
            ce => 'H',
            sr => \N__9353\
        );

    \TACKn_obuft_RNO_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3631\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_677_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIVAPS2_3_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__3773\,
            in1 => \N__4929\,
            in2 => \N__4968\,
            in3 => \N__4676\,
            lcout => \U712_REG_SM.N_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__3834\,
            in1 => \N__7816\,
            in2 => \_gnd_net_\,
            in3 => \N__3871\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9573\,
            ce => \N__3805\,
            sr => \N__9339\
        );

    \U712_REG_SM.C3_SYNC_2_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3957\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9555\,
            ce => 'H',
            sr => \N__9349\
        );

    \U712_REG_SM.C1_SYNC_2_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4243\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9555\,
            ce => 'H',
            sr => \N__9349\
        );

    \U712_REG_SM.C3_SYNC_1_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5044\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9555\,
            ce => 'H',
            sr => \N__9349\
        );

    \U712_REG_SM.C1_SYNC_1_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4023\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9555\,
            ce => 'H',
            sr => \N__9349\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110110000"
        )
    port map (
            in0 => \N__4066\,
            in1 => \N__3754\,
            in2 => \N__3781\,
            in3 => \N__4022\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9555\,
            ce => 'H',
            sr => \N__9349\
        );

    \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3976\,
            in2 => \_gnd_net_\,
            in3 => \N__3951\,
            lcout => \U712_REG_SM.N_68\,
            ltout => \U712_REG_SM.N_68_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI1FQR1_2_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__5038\,
            in1 => \N__4213\,
            in2 => \N__3742\,
            in3 => \N__4239\,
            lcout => \U712_REG_SM.N_73\,
            ltout => \U712_REG_SM.N_73_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4969\,
            in1 => \N__4930\,
            in2 => \N__3739\,
            in3 => \N__4017\,
            lcout => \U712_REG_SM.N_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4101\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4041\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4188\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => 'H',
            sr => \N__9340\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111100011111100"
        )
    port map (
            in0 => \N__3924\,
            in1 => \N__3723\,
            in2 => \N__4189\,
            in3 => \N__3885\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => 'H',
            sr => \N__9340\
        );

    \U712_REG_SM.C1_SYNC_0_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3711\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => 'H',
            sr => \N__9340\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000110000"
        )
    port map (
            in0 => \N__4159\,
            in1 => \N__3883\,
            in2 => \N__3853\,
            in3 => \N__3832\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => 'H',
            sr => \N__9340\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4171\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => 'H',
            sr => \N__9340\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__3923\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3884\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => 'H',
            sr => \N__9340\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110001000"
        )
    port map (
            in0 => \N__3886\,
            in1 => \N__3922\,
            in2 => \N__3835\,
            in3 => \N__3870\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9565\,
            ce => 'H',
            sr => \N__9340\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__7815\,
            in1 => \N__3869\,
            in2 => \N__3852\,
            in3 => \N__3833\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_45_0_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3808\,
            in3 => \N__9411\,
            lcout => \U712_CYCLE_TERM.N_45_0_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9173\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8116\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIFFKI2_4_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110001"
        )
    port map (
            in0 => \N__4065\,
            in1 => \N__4083\,
            in2 => \N__3780\,
            in3 => \N__4021\,
            lcout => \U712_REG_SM.un1_STATE_COUNT_5_0_1\,
            ltout => \U712_REG_SM.un1_STATE_COUNT_5_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__3979\,
            in1 => \N__3956\,
            in2 => \N__3757\,
            in3 => \N__4455\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9550\,
            ce => 'H',
            sr => \N__9344\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__4111\,
            in1 => \N__8267\,
            in2 => \N__4105\,
            in3 => \N__4195\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9550\,
            ce => 'H',
            sr => \N__9344\
        );

    \U712_REG_SM.STATE_COUNT_RNI1VLC2_5_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__4454\,
            in1 => \N__3978\,
            in2 => \N__3958\,
            in3 => \N__4082\,
            lcout => \U712_REG_SM.N_173_0\,
            ltout => \U712_REG_SM.N_173_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8189\,
            in2 => \N__4069\,
            in3 => \N__4064\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_54_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__6415\,
            in1 => \N__4042\,
            in2 => \N__4051\,
            in3 => \N__4048\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9550\,
            ce => 'H',
            sr => \N__9344\
        );

    \U712_REG_SM.C1_SYNC_RNIOEF21_2_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__5036\,
            in1 => \N__4215\,
            in2 => \_gnd_net_\,
            in3 => \N__4240\,
            lcout => \U712_REG_SM.N_183_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8179\,
            in2 => \_gnd_net_\,
            in3 => \N__4020\,
            lcout => \U712_REG_SM.RnW_m\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4018\,
            in1 => \N__4214\,
            in2 => \N__5043\,
            in3 => \N__4241\,
            lcout => \U712_REG_SM.N_162_0\,
            ltout => \U712_REG_SM.N_162_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4440\,
            in2 => \N__4030\,
            in3 => \N__4470\,
            lcout => \U712_REG_SM.N_171_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIQU741_2_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4019\,
            in1 => \N__3977\,
            in2 => \_gnd_net_\,
            in3 => \N__3952\,
            lcout => \U712_REG_SM.N_165_0\,
            ltout => \U712_REG_SM.N_165_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4242\,
            in1 => \N__5037\,
            in2 => \N__4219\,
            in3 => \N__4216\,
            lcout => \U712_REG_SM.N_167_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8096\,
            in2 => \_gnd_net_\,
            in3 => \N__6981\,
            lcout => \U712_CHIP_RAM.CPU_TACK_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4184\,
            in2 => \_gnd_net_\,
            in3 => \N__4170\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__4117\,
            in1 => \N__8104\,
            in2 => \N__8702\,
            in3 => \N__6001\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__8105\,
            in1 => \N__4153\,
            in2 => \N__4138\,
            in3 => \N__4135\,
            lcout => \U712_CHIP_RAM.N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5152\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9526\,
            ce => \N__8953\,
            sr => \N__9354\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIAEJU_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6387\,
            in2 => \_gnd_net_\,
            in3 => \N__6863\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__6864\,
            in1 => \N__6982\,
            in2 => \N__7894\,
            in3 => \N__8349\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6411\,
            in1 => \N__6450\,
            in2 => \_gnd_net_\,
            in3 => \N__6426\,
            lcout => \U712_REG_SM.DS_EN_0_sqmuxa_1\,
            ltout => \U712_REG_SM.DS_EN_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__4733\,
            in1 => \N__4712\,
            in2 => \N__4477\,
            in3 => \N__4263\,
            lcout => \U712_REG_SM.un1_LDS_OUT_0_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111011"
        )
    port map (
            in0 => \N__4332\,
            in1 => \N__4343\,
            in2 => \N__4381\,
            in3 => \N__4441\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_188_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__4345\,
            in1 => \N__4474\,
            in2 => \N__4459\,
            in3 => \N__4456\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9551\,
            ce => 'H',
            sr => \N__9329\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__4734\,
            in1 => \N__4713\,
            in2 => \_gnd_net_\,
            in3 => \N__4264\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9551\,
            ce => 'H',
            sr => \N__9329\
        );

    \U712_REG_SM.REGENn_1_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__4397\,
            in1 => \N__4353\,
            in2 => \_gnd_net_\,
            in3 => \N__4265\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9551\,
            ce => 'H',
            sr => \N__9329\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__4344\,
            in1 => \N__4377\,
            in2 => \N__4333\,
            in3 => \N__4354\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9551\,
            ce => 'H',
            sr => \N__9329\
        );

    \U712_REG_SM.UDS_OUT_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011111110000"
        )
    port map (
            in0 => \N__4654\,
            in1 => \N__4621\,
            in2 => \N__4869\,
            in3 => \N__4266\,
            lcout => \U712_REG_SM.UDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9556\,
            ce => 'H',
            sr => \N__9322\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110001"
        )
    port map (
            in0 => \N__4316\,
            in1 => \N__4294\,
            in2 => \N__5062\,
            in3 => \N__8075\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9556\,
            ce => 'H',
            sr => \N__9322\
        );

    \U712_REG_SM.LDS_OUT_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011111010"
        )
    port map (
            in0 => \N__4267\,
            in1 => \N__4627\,
            in2 => \N__6288\,
            in3 => \N__4653\,
            lcout => \U712_REG_SM.LDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9556\,
            ce => 'H',
            sr => \N__9322\
        );

    \U712_BYTE_ENABLE.LW_TRANS_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__4652\,
            in1 => \N__4902\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_BYTE_ENABLE.LW_TRANS_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDS_OUT_RNO_0_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5475\,
            in2 => \_gnd_net_\,
            in3 => \N__8163\,
            lcout => \U712_REG_SM.LDS_OUT_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_RNO_0_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__5476\,
            in1 => \_gnd_net_\,
            in2 => \N__8178\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.UDS_OUT_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__5221\,
            in1 => \_gnd_net_\,
            in2 => \N__8821\,
            in3 => \N__8530\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9522\,
            ce => \N__7395\,
            sr => \N__9352\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100011"
        )
    port map (
            in0 => \N__4600\,
            in1 => \N__8691\,
            in2 => \N__8539\,
            in3 => \N__8812\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9522\,
            ce => \N__7395\,
            sr => \N__9352\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8811\,
            in2 => \N__8540\,
            in3 => \N__4525\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9522\,
            ce => \N__7395\,
            sr => \N__9352\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__8695\,
            in1 => \N__4744\,
            in2 => \N__8121\,
            in3 => \N__5113\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__8092\,
            in1 => \N__4564\,
            in2 => \N__4543\,
            in3 => \N__4540\,
            lcout => \U712_CHIP_RAM.N_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010101"
        )
    port map (
            in0 => \N__5095\,
            in1 => \N__4519\,
            in2 => \N__4501\,
            in3 => \N__8090\,
            lcout => \U712_CHIP_RAM.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__8089\,
            in1 => \N__6565\,
            in2 => \N__8699\,
            in3 => \N__5107\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__4822\,
            in1 => \N__4807\,
            in2 => \N__4789\,
            in3 => \N__8091\,
            lcout => \U712_CHIP_RAM.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__4750\,
            in1 => \N__8065\,
            in2 => \N__8703\,
            in3 => \N__5158\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__8066\,
            in1 => \N__4786\,
            in2 => \N__4771\,
            in3 => \N__4768\,
            lcout => \U712_CHIP_RAM.N_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6549\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9530\,
            ce => \N__8935\,
            sr => \N__9338\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5184\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9530\,
            ce => \N__8935\,
            sr => \N__9338\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100000010"
        )
    port map (
            in0 => \N__5617\,
            in1 => \N__6388\,
            in2 => \N__6873\,
            in3 => \N__8024\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9534\,
            ce => 'H',
            sr => \N__9328\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__4735\,
            in1 => \N__4717\,
            in2 => \N__4680\,
            in3 => \N__4696\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9544\,
            ce => 'H',
            sr => \N__9321\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4917\,
            in1 => \N__4948\,
            in2 => \_gnd_net_\,
            in3 => \N__5055\,
            lcout => \U712_CHIP_RAM.un1_DBR_SYNC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111100"
        )
    port map (
            in0 => \N__6305\,
            in1 => \N__5039\,
            in2 => \N__5002\,
            in3 => \N__4990\,
            lcout => \U712_REG_SM.DS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9544\,
            ce => 'H',
            sr => \N__9321\
        );

    \U712_CHIP_RAM.DBR_SYNC_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4984\,
            lcout => \U712_REG_SM_DBR_SYNC_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9549\,
            ce => 'H',
            sr => \N__9320\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4955\,
            lcout => \U712_REG_SM_DBR_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9549\,
            ce => 'H',
            sr => \N__9320\
        );

    \U712_BYTE_ENABLE.LLBE_0_tz_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5477\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4906\,
            lcout => \U712_BYTE_ENABLE.LLBE_0_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_RNIUP9B_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4870\,
            in2 => \_gnd_net_\,
            in3 => \N__6312\,
            lcout => \U712_REG_SM_un1_UDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7780\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5643\,
            in2 => \_gnd_net_\,
            in3 => \N__5658\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__5694\,
            in1 => \N__5709\,
            in2 => \N__5677\,
            in3 => \N__5724\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__8680\,
            in1 => \N__5827\,
            in2 => \N__8122\,
            in3 => \N__5992\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8103\,
            in1 => \N__5263\,
            in2 => \N__5245\,
            in3 => \N__5242\,
            lcout => \U712_CHIP_RAM.N_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010101011"
        )
    port map (
            in0 => \N__5215\,
            in1 => \N__8816\,
            in2 => \N__8541\,
            in3 => \N__8690\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9524\,
            ce => \N__7394\,
            sr => \N__9363\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5185\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9527\,
            ce => \N__9064\,
            sr => \N__9355\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5148\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9527\,
            ce => \N__9064\,
            sr => \N__9355\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5818\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9527\,
            ce => \N__9064\,
            sr => \N__9355\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5089\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9527\,
            ce => \N__9064\,
            sr => \N__9355\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__8644\,
            in1 => \N__5794\,
            in2 => \N__8088\,
            in3 => \N__5101\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5088\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9531\,
            ce => \N__8945\,
            sr => \N__9350\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__5374\,
            in1 => \N__8769\,
            in2 => \_gnd_net_\,
            in3 => \N__8511\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9538\,
            ce => \N__7396\,
            sr => \N__9345\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__5347\,
            in1 => \N__6088\,
            in2 => \N__5329\,
            in3 => \N__8023\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8768\,
            in2 => \N__5305\,
            in3 => \N__8510\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9538\,
            ce => \N__7396\,
            sr => \N__9345\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__6069\,
            in1 => \N__5281\,
            in2 => \N__6055\,
            in3 => \N__7193\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9545\,
            ce => \N__6123\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__5404\,
            in1 => \N__7798\,
            in2 => \_gnd_net_\,
            in3 => \N__7236\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7014\,
            in1 => \N__7060\,
            in2 => \N__7089\,
            in3 => \N__7111\,
            lcout => \U712_CHIP_RAM.N_61\,
            ltout => \U712_CHIP_RAM.N_61_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5275\,
            in3 => \N__7855\,
            lcout => \U712_CHIP_RAM.N_65\,
            ltout => \U712_CHIP_RAM.N_65_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101011101"
        )
    port map (
            in0 => \N__7799\,
            in1 => \N__5269\,
            in2 => \N__5272\,
            in3 => \N__7701\,
            lcout => \U712_CHIP_RAM.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_1_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__6847\,
            in1 => \_gnd_net_\,
            in2 => \N__6976\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_104_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI399Q7_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000110011"
        )
    port map (
            in0 => \N__7251\,
            in1 => \N__7192\,
            in2 => \N__6019\,
            in3 => \N__7702\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER16_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIEBLDE_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__5403\,
            in1 => \N__8218\,
            in2 => \N__5392\,
            in3 => \N__6081\,
            lcout => \U712_CHIP_RAM.N_158_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8350\,
            in1 => \N__7576\,
            in2 => \N__6874\,
            in3 => \N__8251\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_0_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__6504\,
            in1 => \_gnd_net_\,
            in2 => \N__5389\,
            in3 => \N__7197\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5386\,
            in3 => \N__9410\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI3EN62_0_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__6380\,
            in1 => \N__7706\,
            in2 => \N__7630\,
            in3 => \N__6336\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_4_1_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6868\,
            in1 => \N__8250\,
            in2 => \N__6977\,
            in3 => \N__7853\,
            lcout => \U712_CHIP_RAM.N_67\,
            ltout => \U712_CHIP_RAM.N_67_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFQROA_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000110111"
        )
    port map (
            in0 => \N__7628\,
            in1 => \N__7707\,
            in2 => \N__5383\,
            in3 => \N__6103\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER18_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER18_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000010"
        )
    port map (
            in0 => \N__7198\,
            in1 => \N__6082\,
            in2 => \N__5380\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_m2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__7808\,
            in1 => \_gnd_net_\,
            in2 => \N__5377\,
            in3 => \N__6053\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9552\,
            ce => \N__6124\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011101110"
        )
    port map (
            in0 => \N__5768\,
            in1 => \N__5616\,
            in2 => \N__8968\,
            in3 => \N__5605\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9557\,
            ce => 'H',
            sr => \N__9323\
        );

    \U712_BYTE_ENABLE.un2_CUMBEn_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100000000"
        )
    port map (
            in0 => \N__5508\,
            in1 => \N__5566\,
            in2 => \N__5436\,
            in3 => \N__8119\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.un2_CUMBEnZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001101"
        )
    port map (
            in0 => \N__9125\,
            in1 => \N__6744\,
            in2 => \N__5593\,
            in3 => \N__5771\,
            lcout => \CUMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un2_CLLBEn_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000000"
        )
    port map (
            in0 => \N__5506\,
            in1 => \N__5565\,
            in2 => \N__5434\,
            in3 => \N__8117\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.un2_CLLBEnZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__9123\,
            in1 => \N__6743\,
            in2 => \N__5557\,
            in3 => \N__5769\,
            lcout => \CLLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un2_CLMBEn_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000000"
        )
    port map (
            in0 => \N__5507\,
            in1 => \N__5478\,
            in2 => \N__5435\,
            in3 => \N__8118\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.un2_CLMBEnZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__9124\,
            in1 => \N__6702\,
            in2 => \N__5533\,
            in3 => \N__5770\,
            lcout => \CLMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un2_CUUBEn_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100000000"
        )
    port map (
            in0 => \N__5509\,
            in1 => \N__5479\,
            in2 => \N__5437\,
            in3 => \N__8120\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.un2_CUUBEnZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001101"
        )
    port map (
            in0 => \N__9126\,
            in1 => \N__6703\,
            in2 => \N__5407\,
            in3 => \N__5772\,
            lcout => \CUUBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5725\,
            in2 => \_gnd_net_\,
            in3 => \N__5713\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_4_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__5626\,
            ce => 'H',
            sr => \N__6010\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5710\,
            in2 => \_gnd_net_\,
            in3 => \N__5698\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__5626\,
            ce => 'H',
            sr => \N__6010\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5695\,
            in2 => \_gnd_net_\,
            in3 => \N__5683\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__5626\,
            ce => 'H',
            sr => \N__6010\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6241\,
            in2 => \_gnd_net_\,
            in3 => \N__5680\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__5626\,
            ce => 'H',
            sr => \N__6010\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5676\,
            in2 => \_gnd_net_\,
            in3 => \N__5662\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__5626\,
            ce => 'H',
            sr => \N__6010\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5659\,
            in2 => \_gnd_net_\,
            in3 => \N__5647\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__5626\,
            ce => 'H',
            sr => \N__6010\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5644\,
            in2 => \_gnd_net_\,
            in3 => \N__5632\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__5626\,
            ce => 'H',
            sr => \N__6010\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6228\,
            in2 => \_gnd_net_\,
            in3 => \N__5629\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5626\,
            ce => 'H',
            sr => \N__6010\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8676\,
            in1 => \N__8515\,
            in2 => \N__8817\,
            in3 => \N__8879\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5860\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9528\,
            ce => \N__9063\,
            sr => \N__9367\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9007\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9528\,
            ce => \N__9063\,
            sr => \N__9367\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_2_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8800\,
            in1 => \N__8663\,
            in2 => \_gnd_net_\,
            in3 => \N__8516\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => \U712_CHIP_RAM.CMA_5_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__7264\,
            in1 => \N__5986\,
            in2 => \N__5965\,
            in3 => \N__8097\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9532\,
            ce => \N__7392\,
            sr => \N__9364\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8801\,
            in1 => \N__5941\,
            in2 => \_gnd_net_\,
            in3 => \N__8517\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9532\,
            ce => \N__7392\,
            sr => \N__9364\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__8407\,
            in1 => \N__5911\,
            in2 => \N__5905\,
            in3 => \N__8098\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9532\,
            ce => \N__7392\,
            sr => \N__9364\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5856\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9539\,
            ce => \N__8920\,
            sr => \N__9356\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5814\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9539\,
            ce => \N__8920\,
            sr => \N__9356\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100110001"
        )
    port map (
            in0 => \N__7795\,
            in1 => \N__6610\,
            in2 => \N__6054\,
            in3 => \N__8468\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9546\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000010011"
        )
    port map (
            in0 => \N__8615\,
            in1 => \N__8866\,
            in2 => \N__8781\,
            in3 => \N__8467\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__6517\,
            in1 => \N__8109\,
            in2 => \N__6097\,
            in3 => \N__8616\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__6807\,
            in1 => \_gnd_net_\,
            in2 => \N__6975\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITC5T1_1_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6846\,
            in1 => \N__6954\,
            in2 => \_gnd_net_\,
            in3 => \N__8348\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001101010101"
        )
    port map (
            in0 => \N__6025\,
            in1 => \N__6070\,
            in2 => \N__6058\,
            in3 => \N__6049\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9553\,
            ce => \N__6601\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__7753\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7235\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_1_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__6806\,
            in1 => \_gnd_net_\,
            in2 => \N__6974\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_2_1_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6804\,
            in2 => \_gnd_net_\,
            in3 => \N__6947\,
            lcout => \U712_CHIP_RAM.N_124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITDHQ2_0_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6805\,
            in1 => \N__7754\,
            in2 => \_gnd_net_\,
            in3 => \N__8249\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_0\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIO007I_0_0_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010101"
        )
    port map (
            in0 => \N__6625\,
            in1 => \N__8323\,
            in2 => \N__6127\,
            in3 => \N__8299\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6990\,
            in1 => \N__7041\,
            in2 => \N__6862\,
            in3 => \N__7523\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_5\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI971H6_2_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__7042\,
            in1 => \N__7033\,
            in2 => \N__6106\,
            in3 => \N__6991\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2VVR2_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7796\,
            in1 => \N__8248\,
            in2 => \N__7708\,
            in3 => \N__7609\,
            lcout => \U712_CHIP_RAM.N_108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__6586\,
            in1 => \N__9413\,
            in2 => \N__7026\,
            in3 => \N__7116\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__6837\,
            in1 => \N__6973\,
            in2 => \_gnd_net_\,
            in3 => \N__6885\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000010010"
        )
    port map (
            in0 => \N__6585\,
            in1 => \N__9412\,
            in2 => \N__7027\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__9415\,
            in1 => \N__6487\,
            in2 => \N__7066\,
            in3 => \N__7088\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__6486\,
            in1 => \N__9414\,
            in2 => \_gnd_net_\,
            in3 => \N__7065\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9558\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6378\,
            in2 => \_gnd_net_\,
            in3 => \N__6861\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9561\,
            ce => \N__6322\,
            sr => \N__9330\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__9409\,
            in1 => \N__6651\,
            in2 => \_gnd_net_\,
            in3 => \N__6665\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001010"
        )
    port map (
            in0 => \N__6652\,
            in1 => \N__9122\,
            in2 => \N__6670\,
            in3 => \N__6377\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9566\,
            ce => 'H',
            sr => \N__9324\
        );

    \U712_REG_SM.LDS_OUT_RNIL31J_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6316\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6292\,
            lcout => \U712_REG_SM_un1_LDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111111101"
        )
    port map (
            in0 => \N__6250\,
            in1 => \N__6240\,
            in2 => \N__6229\,
            in3 => \N__6214\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9523\,
            ce => 'H',
            sr => \N__9376\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__6139\,
            in1 => \N__8820\,
            in2 => \_gnd_net_\,
            in3 => \N__8534\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9525\,
            ce => \N__7379\,
            sr => \N__9374\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__6184\,
            in1 => \N__6133\,
            in2 => \N__6163\,
            in3 => \N__8123\,
            lcout => \U712_CHIP_RAM.N_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__6556\,
            in1 => \N__8099\,
            in2 => \N__8700\,
            in3 => \N__7303\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7330\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9540\,
            ce => \N__8952\,
            sr => \N__9368\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7297\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9540\,
            ce => \N__8952\,
            sr => \N__9368\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6550\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9547\,
            ce => \N__9059\,
            sr => \N__9365\
        );

    \U712_CHIP_RAM.DBDIR_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000001110100"
        )
    port map (
            in0 => \N__7933\,
            in1 => \N__6511\,
            in2 => \N__7460\,
            in3 => \N__7219\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9554\,
            ce => 'H',
            sr => \N__9357\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9417\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6493\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7117\,
            in1 => \N__7025\,
            in2 => \_gnd_net_\,
            in3 => \N__6584\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111100101010"
        )
    port map (
            in0 => \N__6475\,
            in1 => \N__6460\,
            in2 => \N__6439\,
            in3 => \N__6404\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9554\,
            ce => 'H',
            sr => \N__9357\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIG7JB2_1_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__7839\,
            in1 => \N__7752\,
            in2 => \N__6853\,
            in3 => \N__6957\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI3EN62_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__6379\,
            in1 => \N__7615\,
            in2 => \N__6343\,
            in3 => \N__7684\,
            lcout => \U712_CHIP_RAM.N_77\,
            ltout => \U712_CHIP_RAM.N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4B3NB_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__6643\,
            in1 => \N__6637\,
            in2 => \N__6628\,
            in3 => \N__7483\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIO007I_0_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__6619\,
            in1 => \N__8322\,
            in2 => \N__6613\,
            in3 => \N__8298\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6604\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6833\,
            in1 => \N__7570\,
            in2 => \_gnd_net_\,
            in3 => \N__7522\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100010010"
        )
    port map (
            in0 => \N__7217\,
            in1 => \N__6571\,
            in2 => \N__6854\,
            in3 => \N__7135\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9559\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVE5T1_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__6958\,
            in1 => \N__7840\,
            in2 => \N__7624\,
            in3 => \N__7683\,
            lcout => \U712_CHIP_RAM.N_121\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI7MV4_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8363\,
            in2 => \_gnd_net_\,
            in3 => \N__8376\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_2_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6956\,
            in1 => \N__7882\,
            in2 => \N__7525\,
            in3 => \N__7682\,
            lcout => \U712_CHIP_RAM.N_122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJ42D8_0_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__6856\,
            in1 => \N__9416\,
            in2 => \N__8272\,
            in3 => \N__8281\,
            lcout => \U712_CHIP_RAM.N_80\,
            ltout => \U712_CHIP_RAM.N_80_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQU7BE_0_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7134\,
            in2 => \N__7123\,
            in3 => \N__7207\,
            lcout => \U712_CHIP_RAM.N_50\,
            ltout => \U712_CHIP_RAM.N_50_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__6857\,
            in1 => \N__7521\,
            in2 => \N__7120\,
            in3 => \N__7575\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9562\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6955\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7881\,
            lcout => \U712_CHIP_RAM.N_127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7112\,
            in1 => \N__7090\,
            in2 => \_gnd_net_\,
            in3 => \N__7061\,
            lcout => \U712_CHIP_RAM.N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISDRT_2_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6855\,
            in2 => \_gnd_net_\,
            in3 => \N__7883\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER39_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_4_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7015\,
            in2 => \_gnd_net_\,
            in3 => \N__6959\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER39_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__6972\,
            in1 => \N__6886\,
            in2 => \N__6872\,
            in3 => \N__7887\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9567\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6745\,
            in2 => \_gnd_net_\,
            in3 => \N__6696\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9571\,
            ce => 'H',
            sr => \N__9331\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6669\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9571\,
            ce => 'H',
            sr => \N__9331\
        );

    \U712_BUFFERS.DRDDIR_0_i_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001010"
        )
    port map (
            in0 => \N__9139\,
            in1 => \N__8200\,
            in2 => \N__7467\,
            in3 => \N__9180\,
            lcout => \DRDDIR_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8819\,
            in1 => \N__8704\,
            in2 => \N__8886\,
            in3 => \N__8538\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9529\,
            ce => \N__7393\,
            sr => \N__9377\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7329\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9541\,
            ce => \N__9058\,
            sr => \N__9370\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7293\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9548\,
            ce => \N__9045\,
            sr => \N__9369\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7680\,
            in1 => \N__7255\,
            in2 => \N__7629\,
            in3 => \N__7240\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER49_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7218\,
            in2 => \N__7162\,
            in3 => \N__8365\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9563\,
            ce => 'H',
            sr => \N__9358\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7159\,
            in1 => \N__9141\,
            in2 => \_gnd_net_\,
            in3 => \N__8127\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9563\,
            ce => 'H',
            sr => \N__9358\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__7681\,
            in1 => \N__7147\,
            in2 => \_gnd_net_\,
            in3 => \N__8321\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9563\,
            ce => 'H',
            sr => \N__9358\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI20AV_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8377\,
            in1 => \N__8364\,
            in2 => \N__7524\,
            in3 => \N__7679\,
            lcout => \U712_CHIP_RAM.N_135\,
            ltout => \U712_CHIP_RAM.N_135_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMMGI5_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__7571\,
            in1 => \N__8320\,
            in2 => \N__8302\,
            in3 => \N__8297\,
            lcout => \U712_CHIP_RAM.N_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7543\,
            in1 => \N__7611\,
            in2 => \N__7854\,
            in3 => \N__7678\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__7900\,
            in1 => \N__8214\,
            in2 => \N__8275\,
            in3 => \N__8271\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9568\,
            ce => 'H',
            sr => \N__9351\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__8199\,
            in1 => \N__9140\,
            in2 => \N__8128\,
            in3 => \N__7929\,
            lcout => \U712_CHIP_RAM.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7513\,
            in2 => \_gnd_net_\,
            in3 => \N__7880\,
            lcout => \U712_CHIP_RAM.N_63\,
            ltout => \U712_CHIP_RAM.N_63_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN14U1_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7797\,
            in1 => \N__7677\,
            in2 => \N__7633\,
            in3 => \N__7610\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIFMO84_3_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__7569\,
            in1 => \N__7542\,
            in2 => \N__7528\,
            in3 => \N__7514\,
            lcout => \U712_CHIP_RAM.N_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9184\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9142\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__9418\,
            in1 => \N__8548\,
            in2 => \_gnd_net_\,
            in3 => \N__9592\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9003\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9572\,
            ce => \N__8934\,
            sr => \N__9359\
        );

    \U712_CHIP_RAM.CRCSn_LC_18_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8887\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9533\,
            ce => 'H',
            sr => \N__9380\
        );

    \U712_CHIP_RAM.RASn_LC_18_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8818\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9542\,
            ce => 'H',
            sr => \N__9379\
        );

    \U712_CHIP_RAM.CASn_LC_18_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8701\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9542\,
            ce => 'H',
            sr => \N__9379\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9591\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9560\,
            ce => 'H',
            sr => \N__9375\
        );

    \U712_CHIP_RAM.WEn_LC_19_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8542\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9543\,
            ce => 'H',
            sr => \N__9381\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_19_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8403\,
            in2 => \_gnd_net_\,
            in3 => \N__9601\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9564\,
            ce => 'H',
            sr => \N__9378\
        );

    \CONSTANT_ONE_LUT4_LC_20_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

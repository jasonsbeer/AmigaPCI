// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 15 2025 11:38:09

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    TM,
    TT,
    D,
    A,
    PIO_S0,
    PORTSIZE,
    TICK60,
    CIACS0n,
    CPUCONFn,
    CLK6,
    CLK_CIA,
    BUFENn,
    AUTOBOOT,
    RnW,
    PIO_P2,
    CIACS1n,
    BRIDGE_ENn,
    PIO_S1,
    PIO_P0,
    TICK50,
    TCIn,
    TBIn,
    RAMSPACEn,
    CLK40_IN,
    CLK28_IN,
    REGSPACEn,
    TSn,
    RTC_ENn,
    PIO_S2,
    ATA_ENn,
    RESETn,
    OVL,
    CONFIGENn,
    TACKn,
    ROMENn,
    PIO_P1);

    input [1:0] TM;
    input [1:0] TT;
    inout [7:4] D;
    input [31:1] A;
    output PIO_S0;
    output PORTSIZE;
    output TICK60;
    output CIACS0n;
    input CPUCONFn;
    input CLK6;
    output CLK_CIA;
    output BUFENn;
    input AUTOBOOT;
    input RnW;
    output PIO_P2;
    output CIACS1n;
    output BRIDGE_ENn;
    output PIO_S1;
    output PIO_P0;
    output TICK50;
    output TCIn;
    output TBIn;
    output RAMSPACEn;
    input CLK40_IN;
    input CLK28_IN;
    output REGSPACEn;
    input TSn;
    output RTC_ENn;
    output PIO_S2;
    output ATA_ENn;
    input RESETn;
    input OVL;
    output CONFIGENn;
    inout TACKn;
    output ROMENn;
    output PIO_P1;

    wire N__11575;
    wire N__11574;
    wire N__11573;
    wire N__11565;
    wire N__11564;
    wire N__11563;
    wire N__11555;
    wire N__11554;
    wire N__11553;
    wire N__11544;
    wire N__11543;
    wire N__11542;
    wire N__11535;
    wire N__11534;
    wire N__11533;
    wire N__11526;
    wire N__11525;
    wire N__11524;
    wire N__11517;
    wire N__11516;
    wire N__11515;
    wire N__11508;
    wire N__11507;
    wire N__11506;
    wire N__11499;
    wire N__11498;
    wire N__11497;
    wire N__11490;
    wire N__11489;
    wire N__11488;
    wire N__11481;
    wire N__11480;
    wire N__11479;
    wire N__11472;
    wire N__11471;
    wire N__11470;
    wire N__11463;
    wire N__11462;
    wire N__11461;
    wire N__11454;
    wire N__11453;
    wire N__11452;
    wire N__11445;
    wire N__11444;
    wire N__11443;
    wire N__11436;
    wire N__11435;
    wire N__11434;
    wire N__11427;
    wire N__11426;
    wire N__11425;
    wire N__11418;
    wire N__11417;
    wire N__11416;
    wire N__11409;
    wire N__11408;
    wire N__11407;
    wire N__11400;
    wire N__11399;
    wire N__11398;
    wire N__11391;
    wire N__11390;
    wire N__11389;
    wire N__11382;
    wire N__11381;
    wire N__11380;
    wire N__11373;
    wire N__11372;
    wire N__11371;
    wire N__11364;
    wire N__11363;
    wire N__11362;
    wire N__11355;
    wire N__11354;
    wire N__11353;
    wire N__11346;
    wire N__11345;
    wire N__11344;
    wire N__11337;
    wire N__11336;
    wire N__11335;
    wire N__11328;
    wire N__11327;
    wire N__11326;
    wire N__11319;
    wire N__11318;
    wire N__11317;
    wire N__11310;
    wire N__11309;
    wire N__11308;
    wire N__11301;
    wire N__11300;
    wire N__11299;
    wire N__11292;
    wire N__11291;
    wire N__11290;
    wire N__11283;
    wire N__11282;
    wire N__11281;
    wire N__11274;
    wire N__11273;
    wire N__11272;
    wire N__11265;
    wire N__11264;
    wire N__11263;
    wire N__11256;
    wire N__11255;
    wire N__11254;
    wire N__11247;
    wire N__11246;
    wire N__11245;
    wire N__11238;
    wire N__11237;
    wire N__11236;
    wire N__11229;
    wire N__11228;
    wire N__11227;
    wire N__11220;
    wire N__11219;
    wire N__11218;
    wire N__11211;
    wire N__11210;
    wire N__11209;
    wire N__11202;
    wire N__11201;
    wire N__11200;
    wire N__11193;
    wire N__11192;
    wire N__11191;
    wire N__11184;
    wire N__11183;
    wire N__11182;
    wire N__11175;
    wire N__11174;
    wire N__11173;
    wire N__11166;
    wire N__11165;
    wire N__11164;
    wire N__11157;
    wire N__11156;
    wire N__11155;
    wire N__11148;
    wire N__11147;
    wire N__11146;
    wire N__11139;
    wire N__11138;
    wire N__11137;
    wire N__11130;
    wire N__11129;
    wire N__11128;
    wire N__11121;
    wire N__11120;
    wire N__11119;
    wire N__11112;
    wire N__11111;
    wire N__11110;
    wire N__11103;
    wire N__11102;
    wire N__11101;
    wire N__11094;
    wire N__11093;
    wire N__11092;
    wire N__11085;
    wire N__11084;
    wire N__11083;
    wire N__11076;
    wire N__11075;
    wire N__11074;
    wire N__11067;
    wire N__11066;
    wire N__11065;
    wire N__11058;
    wire N__11057;
    wire N__11056;
    wire N__11049;
    wire N__11048;
    wire N__11047;
    wire N__11040;
    wire N__11039;
    wire N__11038;
    wire N__11031;
    wire N__11030;
    wire N__11029;
    wire N__11022;
    wire N__11021;
    wire N__11020;
    wire N__11013;
    wire N__11012;
    wire N__11011;
    wire N__11004;
    wire N__11003;
    wire N__11002;
    wire N__10995;
    wire N__10994;
    wire N__10993;
    wire N__10986;
    wire N__10985;
    wire N__10984;
    wire N__10967;
    wire N__10964;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10954;
    wire N__10951;
    wire N__10950;
    wire N__10947;
    wire N__10944;
    wire N__10941;
    wire N__10934;
    wire N__10933;
    wire N__10930;
    wire N__10929;
    wire N__10926;
    wire N__10923;
    wire N__10920;
    wire N__10919;
    wire N__10918;
    wire N__10917;
    wire N__10916;
    wire N__10915;
    wire N__10914;
    wire N__10913;
    wire N__10908;
    wire N__10905;
    wire N__10900;
    wire N__10897;
    wire N__10894;
    wire N__10893;
    wire N__10890;
    wire N__10889;
    wire N__10888;
    wire N__10885;
    wire N__10884;
    wire N__10881;
    wire N__10880;
    wire N__10879;
    wire N__10872;
    wire N__10871;
    wire N__10868;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10827;
    wire N__10826;
    wire N__10825;
    wire N__10818;
    wire N__10817;
    wire N__10816;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10794;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10782;
    wire N__10777;
    wire N__10774;
    wire N__10773;
    wire N__10770;
    wire N__10761;
    wire N__10758;
    wire N__10755;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10741;
    wire N__10736;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10714;
    wire N__10711;
    wire N__10708;
    wire N__10705;
    wire N__10702;
    wire N__10699;
    wire N__10696;
    wire N__10693;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10666;
    wire N__10663;
    wire N__10660;
    wire N__10655;
    wire N__10652;
    wire N__10651;
    wire N__10648;
    wire N__10645;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10609;
    wire N__10606;
    wire N__10603;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10586;
    wire N__10583;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10571;
    wire N__10570;
    wire N__10569;
    wire N__10568;
    wire N__10567;
    wire N__10566;
    wire N__10565;
    wire N__10564;
    wire N__10563;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10537;
    wire N__10536;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10514;
    wire N__10511;
    wire N__10510;
    wire N__10509;
    wire N__10506;
    wire N__10505;
    wire N__10504;
    wire N__10503;
    wire N__10498;
    wire N__10495;
    wire N__10492;
    wire N__10487;
    wire N__10478;
    wire N__10477;
    wire N__10474;
    wire N__10471;
    wire N__10466;
    wire N__10463;
    wire N__10462;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10450;
    wire N__10447;
    wire N__10444;
    wire N__10441;
    wire N__10438;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10426;
    wire N__10423;
    wire N__10420;
    wire N__10417;
    wire N__10414;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10363;
    wire N__10360;
    wire N__10357;
    wire N__10352;
    wire N__10349;
    wire N__10348;
    wire N__10345;
    wire N__10342;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10327;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10298;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10286;
    wire N__10283;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10238;
    wire N__10237;
    wire N__10234;
    wire N__10231;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10180;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10148;
    wire N__10147;
    wire N__10146;
    wire N__10145;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10127;
    wire N__10126;
    wire N__10125;
    wire N__10124;
    wire N__10123;
    wire N__10122;
    wire N__10119;
    wire N__10116;
    wire N__10109;
    wire N__10104;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10088;
    wire N__10087;
    wire N__10086;
    wire N__10083;
    wire N__10082;
    wire N__10079;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10061;
    wire N__10060;
    wire N__10059;
    wire N__10056;
    wire N__10051;
    wire N__10046;
    wire N__10045;
    wire N__10044;
    wire N__10041;
    wire N__10038;
    wire N__10035;
    wire N__10028;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__10000;
    wire N__9999;
    wire N__9998;
    wire N__9993;
    wire N__9990;
    wire N__9987;
    wire N__9980;
    wire N__9979;
    wire N__9978;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9964;
    wire N__9961;
    wire N__9960;
    wire N__9955;
    wire N__9952;
    wire N__9947;
    wire N__9946;
    wire N__9945;
    wire N__9944;
    wire N__9941;
    wire N__9936;
    wire N__9933;
    wire N__9930;
    wire N__9923;
    wire N__9922;
    wire N__9919;
    wire N__9916;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9883;
    wire N__9882;
    wire N__9879;
    wire N__9876;
    wire N__9873;
    wire N__9872;
    wire N__9871;
    wire N__9870;
    wire N__9869;
    wire N__9868;
    wire N__9865;
    wire N__9862;
    wire N__9859;
    wire N__9854;
    wire N__9847;
    wire N__9836;
    wire N__9833;
    wire N__9832;
    wire N__9831;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9819;
    wire N__9818;
    wire N__9817;
    wire N__9816;
    wire N__9815;
    wire N__9814;
    wire N__9811;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9793;
    wire N__9782;
    wire N__9781;
    wire N__9778;
    wire N__9777;
    wire N__9776;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9766;
    wire N__9765;
    wire N__9762;
    wire N__9761;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9743;
    wire N__9736;
    wire N__9733;
    wire N__9728;
    wire N__9719;
    wire N__9718;
    wire N__9715;
    wire N__9712;
    wire N__9707;
    wire N__9706;
    wire N__9703;
    wire N__9700;
    wire N__9697;
    wire N__9692;
    wire N__9689;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9653;
    wire N__9650;
    wire N__9649;
    wire N__9646;
    wire N__9643;
    wire N__9638;
    wire N__9637;
    wire N__9636;
    wire N__9633;
    wire N__9630;
    wire N__9629;
    wire N__9626;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9608;
    wire N__9607;
    wire N__9604;
    wire N__9601;
    wire N__9596;
    wire N__9593;
    wire N__9590;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9571;
    wire N__9568;
    wire N__9565;
    wire N__9560;
    wire N__9557;
    wire N__9556;
    wire N__9555;
    wire N__9554;
    wire N__9553;
    wire N__9552;
    wire N__9551;
    wire N__9548;
    wire N__9539;
    wire N__9534;
    wire N__9527;
    wire N__9526;
    wire N__9525;
    wire N__9524;
    wire N__9523;
    wire N__9522;
    wire N__9519;
    wire N__9518;
    wire N__9517;
    wire N__9508;
    wire N__9499;
    wire N__9494;
    wire N__9493;
    wire N__9492;
    wire N__9489;
    wire N__9486;
    wire N__9483;
    wire N__9482;
    wire N__9481;
    wire N__9480;
    wire N__9479;
    wire N__9470;
    wire N__9463;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9448;
    wire N__9445;
    wire N__9442;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9424;
    wire N__9421;
    wire N__9418;
    wire N__9413;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9401;
    wire N__9400;
    wire N__9397;
    wire N__9394;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9382;
    wire N__9379;
    wire N__9378;
    wire N__9373;
    wire N__9370;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9286;
    wire N__9283;
    wire N__9280;
    wire N__9275;
    wire N__9274;
    wire N__9271;
    wire N__9268;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9256;
    wire N__9253;
    wire N__9250;
    wire N__9245;
    wire N__9242;
    wire N__9241;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9224;
    wire N__9221;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9127;
    wire N__9126;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9108;
    wire N__9105;
    wire N__9100;
    wire N__9095;
    wire N__9092;
    wire N__9091;
    wire N__9088;
    wire N__9085;
    wire N__9084;
    wire N__9079;
    wire N__9076;
    wire N__9071;
    wire N__9070;
    wire N__9069;
    wire N__9066;
    wire N__9063;
    wire N__9060;
    wire N__9053;
    wire N__9052;
    wire N__9051;
    wire N__9048;
    wire N__9045;
    wire N__9042;
    wire N__9039;
    wire N__9032;
    wire N__9029;
    wire N__9028;
    wire N__9027;
    wire N__9024;
    wire N__9021;
    wire N__9018;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8980;
    wire N__8977;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8948;
    wire N__8947;
    wire N__8946;
    wire N__8943;
    wire N__8940;
    wire N__8937;
    wire N__8934;
    wire N__8931;
    wire N__8928;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8854;
    wire N__8851;
    wire N__8848;
    wire N__8843;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8835;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8825;
    wire N__8822;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8808;
    wire N__8805;
    wire N__8798;
    wire N__8795;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8782;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8767;
    wire N__8766;
    wire N__8765;
    wire N__8764;
    wire N__8763;
    wire N__8762;
    wire N__8753;
    wire N__8746;
    wire N__8741;
    wire N__8740;
    wire N__8739;
    wire N__8738;
    wire N__8737;
    wire N__8734;
    wire N__8731;
    wire N__8730;
    wire N__8727;
    wire N__8726;
    wire N__8715;
    wire N__8710;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8698;
    wire N__8697;
    wire N__8696;
    wire N__8695;
    wire N__8694;
    wire N__8689;
    wire N__8680;
    wire N__8675;
    wire N__8674;
    wire N__8673;
    wire N__8672;
    wire N__8671;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8663;
    wire N__8658;
    wire N__8655;
    wire N__8646;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8629;
    wire N__8628;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8616;
    wire N__8609;
    wire N__8608;
    wire N__8605;
    wire N__8602;
    wire N__8597;
    wire N__8596;
    wire N__8595;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8583;
    wire N__8576;
    wire N__8575;
    wire N__8574;
    wire N__8573;
    wire N__8572;
    wire N__8571;
    wire N__8570;
    wire N__8569;
    wire N__8568;
    wire N__8567;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8539;
    wire N__8536;
    wire N__8533;
    wire N__8530;
    wire N__8527;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8501;
    wire N__8500;
    wire N__8497;
    wire N__8494;
    wire N__8493;
    wire N__8492;
    wire N__8491;
    wire N__8488;
    wire N__8485;
    wire N__8480;
    wire N__8479;
    wire N__8476;
    wire N__8475;
    wire N__8474;
    wire N__8473;
    wire N__8472;
    wire N__8467;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8451;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8439;
    wire N__8434;
    wire N__8431;
    wire N__8428;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8406;
    wire N__8401;
    wire N__8398;
    wire N__8393;
    wire N__8390;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8382;
    wire N__8377;
    wire N__8374;
    wire N__8369;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8352;
    wire N__8351;
    wire N__8350;
    wire N__8347;
    wire N__8342;
    wire N__8337;
    wire N__8334;
    wire N__8333;
    wire N__8328;
    wire N__8327;
    wire N__8324;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8306;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8260;
    wire N__8259;
    wire N__8258;
    wire N__8257;
    wire N__8254;
    wire N__8253;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire N__8226;
    wire N__8221;
    wire N__8214;
    wire N__8211;
    wire N__8206;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8191;
    wire N__8190;
    wire N__8187;
    wire N__8184;
    wire N__8181;
    wire N__8178;
    wire N__8175;
    wire N__8172;
    wire N__8169;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8144;
    wire N__8143;
    wire N__8140;
    wire N__8137;
    wire N__8132;
    wire N__8131;
    wire N__8130;
    wire N__8125;
    wire N__8122;
    wire N__8117;
    wire N__8116;
    wire N__8115;
    wire N__8114;
    wire N__8113;
    wire N__8108;
    wire N__8107;
    wire N__8104;
    wire N__8101;
    wire N__8098;
    wire N__8097;
    wire N__8096;
    wire N__8095;
    wire N__8092;
    wire N__8081;
    wire N__8076;
    wire N__8071;
    wire N__8070;
    wire N__8067;
    wire N__8064;
    wire N__8061;
    wire N__8054;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8039;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8029;
    wire N__8026;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8014;
    wire N__8011;
    wire N__8008;
    wire N__8003;
    wire N__8002;
    wire N__8001;
    wire N__8000;
    wire N__7999;
    wire N__7998;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7971;
    wire N__7968;
    wire N__7965;
    wire N__7964;
    wire N__7963;
    wire N__7960;
    wire N__7957;
    wire N__7956;
    wire N__7955;
    wire N__7952;
    wire N__7951;
    wire N__7950;
    wire N__7949;
    wire N__7948;
    wire N__7947;
    wire N__7944;
    wire N__7943;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7891;
    wire N__7890;
    wire N__7889;
    wire N__7886;
    wire N__7879;
    wire N__7874;
    wire N__7873;
    wire N__7872;
    wire N__7869;
    wire N__7864;
    wire N__7859;
    wire N__7856;
    wire N__7853;
    wire N__7850;
    wire N__7847;
    wire N__7844;
    wire N__7843;
    wire N__7840;
    wire N__7837;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7811;
    wire N__7810;
    wire N__7807;
    wire N__7804;
    wire N__7801;
    wire N__7796;
    wire N__7793;
    wire N__7792;
    wire N__7789;
    wire N__7786;
    wire N__7783;
    wire N__7780;
    wire N__7775;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7756;
    wire N__7753;
    wire N__7750;
    wire N__7749;
    wire N__7744;
    wire N__7741;
    wire N__7738;
    wire N__7735;
    wire N__7730;
    wire N__7727;
    wire N__7724;
    wire N__7723;
    wire N__7722;
    wire N__7719;
    wire N__7714;
    wire N__7709;
    wire N__7708;
    wire N__7707;
    wire N__7706;
    wire N__7703;
    wire N__7702;
    wire N__7699;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7683;
    wire N__7676;
    wire N__7675;
    wire N__7674;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7662;
    wire N__7655;
    wire N__7654;
    wire N__7651;
    wire N__7648;
    wire N__7643;
    wire N__7640;
    wire N__7639;
    wire N__7636;
    wire N__7633;
    wire N__7632;
    wire N__7629;
    wire N__7624;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7601;
    wire N__7600;
    wire N__7599;
    wire N__7596;
    wire N__7591;
    wire N__7588;
    wire N__7585;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7570;
    wire N__7569;
    wire N__7566;
    wire N__7561;
    wire N__7556;
    wire N__7555;
    wire N__7550;
    wire N__7547;
    wire N__7546;
    wire N__7545;
    wire N__7544;
    wire N__7541;
    wire N__7540;
    wire N__7537;
    wire N__7528;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7516;
    wire N__7515;
    wire N__7512;
    wire N__7507;
    wire N__7504;
    wire N__7499;
    wire N__7496;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7486;
    wire N__7481;
    wire N__7480;
    wire N__7477;
    wire N__7476;
    wire N__7473;
    wire N__7470;
    wire N__7467;
    wire N__7464;
    wire N__7463;
    wire N__7462;
    wire N__7455;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7430;
    wire N__7427;
    wire N__7422;
    wire N__7417;
    wire N__7414;
    wire N__7411;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7399;
    wire N__7396;
    wire N__7393;
    wire N__7388;
    wire N__7387;
    wire N__7386;
    wire N__7381;
    wire N__7380;
    wire N__7377;
    wire N__7374;
    wire N__7371;
    wire N__7370;
    wire N__7367;
    wire N__7362;
    wire N__7359;
    wire N__7358;
    wire N__7355;
    wire N__7354;
    wire N__7351;
    wire N__7348;
    wire N__7345;
    wire N__7342;
    wire N__7339;
    wire N__7334;
    wire N__7331;
    wire N__7326;
    wire N__7321;
    wire N__7316;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7286;
    wire N__7285;
    wire N__7282;
    wire N__7279;
    wire N__7274;
    wire N__7271;
    wire N__7270;
    wire N__7267;
    wire N__7264;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7245;
    wire N__7240;
    wire N__7237;
    wire N__7236;
    wire N__7235;
    wire N__7234;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7181;
    wire N__7178;
    wire N__7175;
    wire N__7174;
    wire N__7169;
    wire N__7166;
    wire N__7165;
    wire N__7162;
    wire N__7159;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7136;
    wire N__7133;
    wire N__7130;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7118;
    wire N__7115;
    wire N__7114;
    wire N__7111;
    wire N__7108;
    wire N__7105;
    wire N__7100;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7081;
    wire N__7078;
    wire N__7075;
    wire N__7070;
    wire N__7069;
    wire N__7068;
    wire N__7067;
    wire N__7066;
    wire N__7065;
    wire N__7064;
    wire N__7063;
    wire N__7062;
    wire N__7061;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7046;
    wire N__7039;
    wire N__7036;
    wire N__7033;
    wire N__7032;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7024;
    wire N__7017;
    wire N__7016;
    wire N__7011;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6992;
    wire N__6989;
    wire N__6984;
    wire N__6981;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6963;
    wire N__6960;
    wire N__6955;
    wire N__6952;
    wire N__6947;
    wire N__6944;
    wire N__6943;
    wire N__6940;
    wire N__6937;
    wire N__6936;
    wire N__6933;
    wire N__6930;
    wire N__6927;
    wire N__6926;
    wire N__6919;
    wire N__6916;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6898;
    wire N__6895;
    wire N__6892;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6874;
    wire N__6871;
    wire N__6868;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6839;
    wire N__6838;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6824;
    wire N__6823;
    wire N__6822;
    wire N__6819;
    wire N__6818;
    wire N__6815;
    wire N__6812;
    wire N__6811;
    wire N__6806;
    wire N__6799;
    wire N__6794;
    wire N__6791;
    wire N__6790;
    wire N__6789;
    wire N__6788;
    wire N__6785;
    wire N__6780;
    wire N__6777;
    wire N__6770;
    wire N__6769;
    wire N__6768;
    wire N__6767;
    wire N__6766;
    wire N__6765;
    wire N__6762;
    wire N__6755;
    wire N__6752;
    wire N__6747;
    wire N__6740;
    wire N__6739;
    wire N__6738;
    wire N__6735;
    wire N__6730;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6718;
    wire N__6715;
    wire N__6714;
    wire N__6713;
    wire N__6710;
    wire N__6707;
    wire N__6702;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6682;
    wire N__6681;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6664;
    wire N__6661;
    wire N__6658;
    wire N__6653;
    wire N__6652;
    wire N__6651;
    wire N__6650;
    wire N__6647;
    wire N__6646;
    wire N__6643;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6631;
    wire N__6630;
    wire N__6625;
    wire N__6620;
    wire N__6617;
    wire N__6616;
    wire N__6613;
    wire N__6606;
    wire N__6603;
    wire N__6596;
    wire N__6593;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6581;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6548;
    wire N__6547;
    wire N__6546;
    wire N__6545;
    wire N__6544;
    wire N__6543;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6508;
    wire N__6505;
    wire N__6502;
    wire N__6497;
    wire N__6496;
    wire N__6493;
    wire N__6492;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6478;
    wire N__6477;
    wire N__6476;
    wire N__6475;
    wire N__6472;
    wire N__6467;
    wire N__6464;
    wire N__6459;
    wire N__6456;
    wire N__6453;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6437;
    wire N__6434;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6415;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6403;
    wire N__6402;
    wire N__6399;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6391;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6363;
    wire N__6362;
    wire N__6359;
    wire N__6354;
    wire N__6351;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6326;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6316;
    wire N__6315;
    wire N__6314;
    wire N__6313;
    wire N__6310;
    wire N__6303;
    wire N__6300;
    wire N__6293;
    wire N__6292;
    wire N__6291;
    wire N__6290;
    wire N__6287;
    wire N__6282;
    wire N__6279;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6241;
    wire N__6238;
    wire N__6235;
    wire N__6230;
    wire N__6227;
    wire N__6226;
    wire N__6225;
    wire N__6224;
    wire N__6223;
    wire N__6222;
    wire N__6221;
    wire N__6218;
    wire N__6213;
    wire N__6208;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6189;
    wire N__6184;
    wire N__6179;
    wire N__6176;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6166;
    wire N__6165;
    wire N__6162;
    wire N__6161;
    wire N__6160;
    wire N__6159;
    wire N__6158;
    wire N__6153;
    wire N__6150;
    wire N__6149;
    wire N__6148;
    wire N__6145;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6124;
    wire N__6121;
    wire N__6120;
    wire N__6115;
    wire N__6112;
    wire N__6107;
    wire N__6102;
    wire N__6099;
    wire N__6096;
    wire N__6083;
    wire N__6080;
    wire N__6079;
    wire N__6078;
    wire N__6077;
    wire N__6076;
    wire N__6075;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6063;
    wire N__6060;
    wire N__6057;
    wire N__6054;
    wire N__6041;
    wire N__6038;
    wire N__6037;
    wire N__6034;
    wire N__6033;
    wire N__6032;
    wire N__6031;
    wire N__6028;
    wire N__6027;
    wire N__6026;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6001;
    wire N__5990;
    wire N__5989;
    wire N__5986;
    wire N__5983;
    wire N__5982;
    wire N__5981;
    wire N__5980;
    wire N__5979;
    wire N__5976;
    wire N__5973;
    wire N__5972;
    wire N__5963;
    wire N__5960;
    wire N__5957;
    wire N__5954;
    wire N__5951;
    wire N__5942;
    wire N__5941;
    wire N__5940;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5927;
    wire N__5926;
    wire N__5925;
    wire N__5924;
    wire N__5921;
    wire N__5916;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5900;
    wire N__5895;
    wire N__5888;
    wire N__5887;
    wire N__5882;
    wire N__5879;
    wire N__5878;
    wire N__5877;
    wire N__5874;
    wire N__5869;
    wire N__5866;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5846;
    wire N__5845;
    wire N__5842;
    wire N__5839;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5825;
    wire N__5824;
    wire N__5819;
    wire N__5818;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5810;
    wire N__5809;
    wire N__5808;
    wire N__5805;
    wire N__5800;
    wire N__5797;
    wire N__5792;
    wire N__5791;
    wire N__5790;
    wire N__5787;
    wire N__5782;
    wire N__5779;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5765;
    wire N__5762;
    wire N__5759;
    wire N__5750;
    wire N__5747;
    wire N__5746;
    wire N__5741;
    wire N__5738;
    wire N__5737;
    wire N__5736;
    wire N__5735;
    wire N__5732;
    wire N__5725;
    wire N__5720;
    wire N__5719;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5705;
    wire N__5704;
    wire N__5703;
    wire N__5698;
    wire N__5695;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5671;
    wire N__5668;
    wire N__5665;
    wire N__5660;
    wire N__5657;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5634;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5618;
    wire N__5615;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5602;
    wire N__5601;
    wire N__5598;
    wire N__5595;
    wire N__5592;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5577;
    wire N__5574;
    wire N__5567;
    wire N__5564;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5554;
    wire N__5549;
    wire N__5546;
    wire N__5545;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5530;
    wire N__5525;
    wire N__5522;
    wire N__5519;
    wire N__5518;
    wire N__5515;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5505;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5450;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5437;
    wire N__5434;
    wire N__5431;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5384;
    wire N__5381;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5345;
    wire N__5342;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5272;
    wire N__5267;
    wire N__5264;
    wire N__5263;
    wire N__5262;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5180;
    wire N__5179;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5164;
    wire N__5161;
    wire N__5160;
    wire N__5157;
    wire N__5154;
    wire N__5151;
    wire N__5148;
    wire N__5145;
    wire N__5142;
    wire N__5139;
    wire N__5134;
    wire N__5129;
    wire N__5126;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5051;
    wire N__5048;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__5002;
    wire N__5001;
    wire N__5000;
    wire N__4999;
    wire N__4998;
    wire N__4997;
    wire N__4996;
    wire N__4991;
    wire N__4984;
    wire N__4983;
    wire N__4978;
    wire N__4977;
    wire N__4974;
    wire N__4973;
    wire N__4972;
    wire N__4971;
    wire N__4966;
    wire N__4963;
    wire N__4962;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4945;
    wire N__4940;
    wire N__4935;
    wire N__4930;
    wire N__4925;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4906;
    wire N__4903;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4885;
    wire N__4884;
    wire N__4883;
    wire N__4882;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4868;
    wire N__4863;
    wire N__4858;
    wire N__4857;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4845;
    wire N__4838;
    wire N__4835;
    wire N__4834;
    wire N__4831;
    wire N__4830;
    wire N__4827;
    wire N__4826;
    wire N__4825;
    wire N__4824;
    wire N__4823;
    wire N__4820;
    wire N__4815;
    wire N__4814;
    wire N__4809;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4784;
    wire N__4783;
    wire N__4778;
    wire N__4775;
    wire N__4770;
    wire N__4767;
    wire N__4762;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4741;
    wire N__4740;
    wire N__4737;
    wire N__4732;
    wire N__4731;
    wire N__4730;
    wire N__4727;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4702;
    wire N__4697;
    wire N__4694;
    wire N__4691;
    wire N__4690;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4669;
    wire N__4666;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4645;
    wire N__4640;
    wire N__4637;
    wire N__4636;
    wire N__4633;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4615;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4585;
    wire N__4584;
    wire N__4581;
    wire N__4576;
    wire N__4571;
    wire N__4570;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4562;
    wire N__4561;
    wire N__4560;
    wire N__4557;
    wire N__4556;
    wire N__4555;
    wire N__4554;
    wire N__4553;
    wire N__4548;
    wire N__4543;
    wire N__4540;
    wire N__4531;
    wire N__4530;
    wire N__4529;
    wire N__4526;
    wire N__4521;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4509;
    wire N__4506;
    wire N__4505;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4481;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4445;
    wire N__4442;
    wire N__4441;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4429;
    wire N__4426;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4378;
    wire N__4377;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4312;
    wire N__4309;
    wire N__4306;
    wire N__4305;
    wire N__4302;
    wire N__4299;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4278;
    wire N__4275;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4261;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4211;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4150;
    wire N__4149;
    wire N__4148;
    wire N__4147;
    wire N__4146;
    wire N__4145;
    wire N__4144;
    wire N__4143;
    wire N__4142;
    wire N__4141;
    wire N__4140;
    wire N__4115;
    wire CLK80_OUT;
    wire A_c_15;
    wire A_c_14;
    wire GNDG0;
    wire VCCG0;
    wire \U409_AUTOCONFIG.N_213_2_cascade_ ;
    wire \U409_AUTOCONFIG.N_249_cascade_ ;
    wire \U409_AUTOCONFIG.N_250_1 ;
    wire \U409_AUTOCONFIG.N_249 ;
    wire \U409_AUTOCONFIG.N_250_1_cascade_ ;
    wire \U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0 ;
    wire \U409_AUTOCONFIG.N_167_cascade_ ;
    wire \U409_AUTOCONFIG.N_233 ;
    wire \U409_AUTOCONFIG.N_231_cascade_ ;
    wire \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_a5_0_0 ;
    wire \U409_AUTOCONFIG.N_212 ;
    wire \U409_AUTOCONFIG.N_213_2 ;
    wire \U409_AUTOCONFIG.N_212_cascade_ ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_3_0_cascade_ ;
    wire \U409_AUTOCONFIG.N_165 ;
    wire \U409_AUTOCONFIG.un1_A_16Z0Z_2 ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_0 ;
    wire A_c_16;
    wire \U409_ADDRESS_DECODE.REG_SPACEZ0Z_0 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_0_0 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_1_0 ;
    wire \U409_AUTOCONFIG.N_168_cascade_ ;
    wire \U409_AUTOCONFIG.N_167 ;
    wire \U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0_cascade_ ;
    wire \U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0 ;
    wire \U409_AUTOCONFIG.N_166 ;
    wire \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ;
    wire \U409_AUTOCONFIG.N_173 ;
    wire \U409_AUTOCONFIG.N_249_1_cascade_ ;
    wire \U409_AUTOCONFIG.N_155_0 ;
    wire A_c_4;
    wire \U409_AUTOCONFIG.un1_A_19Z0Z_1_cascade_ ;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn_i;
    wire \U409_ADDRESS_DECODE.un2_REGSPACEn_0_0 ;
    wire \U409_ADDRESS_DECODE.REG_SPACEZ0 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_ ;
    wire A_c_2;
    wire \U409_AUTOCONFIG.un1_A_11Z0Z_0_cascade_ ;
    wire \U409_AUTOCONFIG.un1_AZ0Z_11 ;
    wire A_c_6;
    wire A_c_3;
    wire \U409_AUTOCONFIG.N_174 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ;
    wire \U409_ADDRESS_DECODE.REG_SPACE_3 ;
    wire A_c_25;
    wire \U409_ADDRESS_DECODE.REG_SPACE_3_cascade_ ;
    wire A_c_24;
    wire A_c_27;
    wire A_c_26;
    wire D_1_i;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ;
    wire U409_AUTOCONFIG_D_OUT_0_i_3;
    wire AUTOCONFIG_SPACE_cascade_;
    wire \U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0_a3_0 ;
    wire CPUCONFn_c;
    wire \U409_AUTOCONFIG.AC_STARTZ0 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ;
    wire U409_AUTOCONFIG_D_OUT_0_i_0;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNO_0Z0Z_1 ;
    wire \U409_AUTOCONFIG.N_265_0 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNO_0Z0Z_0 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ;
    wire \U409_AUTOCONFIG.un1_STATE_8_0_0 ;
    wire \U409_AUTOCONFIG.STATE4 ;
    wire \U409_AUTOCONFIG.un1_STATE_8Z0Z_0 ;
    wire \U409_AUTOCONFIG.N_248_0 ;
    wire \U409_AUTOCONFIG.un1_STATE_8Z0Z_0_cascade_ ;
    wire \INVU409_AUTOCONFIG.LIDE_OUT_1C_net ;
    wire \INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net ;
    wire U409_ADDRESS_DECODE_un1_RTC_ENn_i;
    wire TT_c_1;
    wire TT_c_0;
    wire \U409_ADDRESS_DECODE.CIA_SPACE_3 ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0 ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_4 ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_ ;
    wire \U409_ADDRESS_DECODE.CIA_SPACE_2_0 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6 ;
    wire \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7 ;
    wire U409_ADDRESS_DECODE_AUTOVECTOR_8;
    wire U409_ADDRESS_DECODE_AUTOVECTOR_10_cascade_;
    wire U409_ADDRESS_DECODE_AUTOVECTOR_9;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ;
    wire U409_AUTOCONFIG_D_OUT_0_i_1;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2 ;
    wire U409_AUTOCONFIG_D_OUT_0_i_2;
    wire \INVU409_AUTOCONFIG.STATE_1C_net ;
    wire \U409_AUTOCONFIG.STATE_d_2_cascade_ ;
    wire A_c_31;
    wire A_c_30;
    wire BRIDGE_BASE_3;
    wire A_c_29;
    wire A_c_28;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2Z0Z_0_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5 ;
    wire CONFIGENn_c;
    wire \INVU409_AUTOCONFIG.AC_TACKC_net ;
    wire A_c_7;
    wire \U409_AUTOCONFIG.ATA_BASE11Z0Z_1 ;
    wire A_c_5;
    wire \U409_AUTOCONFIG.STATEZ0Z_1 ;
    wire \U409_AUTOCONFIG.ATA_BASE11_cascade_ ;
    wire \U409_AUTOCONFIG.STATEZ0Z_0 ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_6 ;
    wire ATA_BASE_6;
    wire D_in_6;
    wire BRIDGE_BASE_2;
    wire A_c_20;
    wire ATA_BASE_4;
    wire \U409_AUTOCONFIG.LIDE_CONF_RNIDFPAZ0Z3 ;
    wire ATA_BASE_5;
    wire \INVU409_AUTOCONFIG.ATA_BASE_6C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_11_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_5_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_2 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ;
    wire \U409_AUTOCONFIG.STATE_d_2 ;
    wire \U409_AUTOCONFIG.un1_AZ0Z_16 ;
    wire \U409_AUTOCONFIG.LIDE_CONFZ0 ;
    wire D_in_4;
    wire BRIDGE_BASE_0;
    wire \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ;
    wire BRIDGE_BASE_1;
    wire \INVU409_AUTOCONFIG.LIDE_CONFC_net ;
    wire A_c_19;
    wire A_c_18;
    wire ATA_BASE_2;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2_cascade_ ;
    wire ATA_BASE_7;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_0 ;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_5_cascade_ ;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_ ;
    wire \U409_AUTOCONFIG.un1_STATE_6_0 ;
    wire A_c_1;
    wire A_c_17;
    wire \U409_ADDRESS_DECODE.un2_ATA_SPACEZ0Z_0 ;
    wire U409_ADDRESS_DECODE_un1_RTC_ENn;
    wire U409_ADDRESS_DECODE_PORTSIZE_0_cascade_;
    wire PORTSIZE_0_i;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.un1_AUTOVECTOR_0 ;
    wire TSn_c;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ;
    wire \U409_TRANSFER_ACK.N_17_mux_cascade_ ;
    wire \U409_TRANSFER_ACK.N_3_0_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0 ;
    wire \U409_TRANSFER_ACK.N_3_0 ;
    wire \U409_TRANSFER_ACK.N_6_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_17_mux ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_0C_net ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1Z0Z_0 ;
    wire A_c_22;
    wire A_c_23;
    wire \U409_TRANSFER_ACK.N_43 ;
    wire ROMENn_c;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0 ;
    wire \INVU409_TRANSFER_ACK.ROMENnC_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire AC_TACK;
    wire \U409_TRANSFER_ACK.TACK_COUNTER5_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ;
    wire \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ;
    wire TACK_OUTn;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_1_out ;
    wire \INVU409_TRANSFER_ACK.TACK_OUTnC_net ;
    wire \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ;
    wire TM_c_0;
    wire TM_c_1;
    wire CONFIGURED;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1 ;
    wire \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_1 ;
    wire \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_2 ;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_ ;
    wire U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i;
    wire RnW_c;
    wire D_in_5;
    wire un1_AUTOCONFIG_SPACE_cascade_;
    wire ATA_BASE_1;
    wire \U409_AUTOCONFIG.STATE_RNIS3FU2Z0Z_0 ;
    wire un1_AUTOCONFIG_SPACE;
    wire D_in_7;
    wire ATA_BASE_3;
    wire \INVU409_AUTOCONFIG.ATA_BASE_1C_net ;
    wire CLK40_IN_c_g;
    wire GB_BUFFER_CLK40_IN_c_g_THRU_CO;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ;
    wire TICK50_c;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn_i;
    wire \U409_TRANSFER_ACK.N_28 ;
    wire \U409_TRANSFER_ACK.N_22 ;
    wire U409_ADDRESS_DECODE_ROMEN_1;
    wire \U409_TRANSFER_ACK.N_33_1 ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0_cascade_ ;
    wire \U409_TRANSFER_ACK.N_33 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_34 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.N_45 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.TACK_ENC_net ;
    wire RESETn_c_i_g;
    wire \U409_ADDRESS_DECODE.un1_REGSPACEnZ0 ;
    wire \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0 ;
    wire A_c_21;
    wire OVL_c;
    wire AGNUS_SPACE_0_cascade_;
    wire TACKn_in;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5 ;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4 ;
    wire BUFENn_c;
    wire U409_ADDRESS_DECODE_PORTSIZE_0;
    wire AGNUS_SPACE_0;
    wire TACK_EN;
    wire TCIn_1_i;
    wire RESETn_c_i;
    wire bfn_13_6_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire bfn_13_7_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_ADDRESS_DECODE.ATA_ENZ0 ;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0 ;
    wire U409_ADDRESS_DECODE_un1_ATA_ENn_i;
    wire \U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_ ;
    wire CIA_SPACE;
    wire \U409_CIA.VMA_RNOZ0Z_0_cascade_ ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.TICK503_8 ;
    wire \U409_TICK.TICK503_11_cascade_ ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire TICK60_c;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.TICK603_11 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.TICK603_8_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire bfn_15_4_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_5 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_6 ;
    wire \U409_CIA.CLK_CIA_r_1_0 ;
    wire \U409_CIA.CLK_CIA6_3_cascade_ ;
    wire CLK_CIA_c;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_7 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_6 ;
    wire \U409_CIA.CLK_CIA6_4 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_0 ;
    wire \U409_CIA.CLK_CIA6_4_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire CLK28_IN_c_g;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire bfn_15_6_0_;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire bfn_15_7_0_;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire CLK6_c_g;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2 ;
    wire CONSTANT_ONE_NET;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_CIACS1n_i;
    wire \U409_CIA.VMAZ0 ;
    wire RESETn_c;
    wire CIA_ENABLE;
    wire A_c_12;
    wire CIA_ENABLE_cascade_;
    wire U409_ADDRESS_DECODE_un1_CIACS0n_i;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__7904),
            .RESETB(N__10466),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11573),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__11575),
            .DIN(N__11574),
            .DOUT(N__11573),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__11575),
            .PADOUT(N__11574),
            .PADIN(N__11573),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11563),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__11565),
            .DIN(N__11564),
            .DOUT(N__11563),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__11565),
            .PADOUT(N__11564),
            .PADIN(N__11563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK40_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11553),
            .GLOBALBUFFEROUTPUT(CLK40_IN_c_g));
    IO_PAD CLK40_IN_ibuf_gb_io_iopad (
            .OE(N__11555),
            .DIN(N__11554),
            .DOUT(N__11553),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_gb_io_preio (
            .PADOEN(N__11555),
            .PADOUT(N__11554),
            .PADIN(N__11553),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11544),
            .DIN(N__11543),
            .DOUT(N__11542),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11544),
            .PADOUT(N__11543),
            .PADIN(N__11542),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__11535),
            .DIN(N__11534),
            .DOUT(N__11533),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__11535),
            .PADOUT(N__11534),
            .PADIN(N__11533),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_P1_obuf_iopad (
            .OE(N__11526),
            .DIN(N__11525),
            .DOUT(N__11524),
            .PACKAGEPIN(PIO_P1));
    defparam PIO_P1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_P1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_P1_obuf_preio (
            .PADOEN(N__11526),
            .PADOUT(N__11525),
            .PADIN(N__11524),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10433),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_7_iopad (
            .OE(N__11517),
            .DIN(N__11516),
            .DOUT(N__11515),
            .PACKAGEPIN(D[7]));
    defparam D_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_7_preio (
            .PADOEN(N__11517),
            .PADOUT(N__11516),
            .PADIN(N__11515),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5178),
            .DIN0(D_in_7),
            .DOUT0(N__5114),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11508),
            .DIN(N__11507),
            .DOUT(N__11506),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11508),
            .PADOUT(N__11507),
            .PADIN(N__11506),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CPUCONFn_ibuf_iopad (
            .OE(N__11499),
            .DIN(N__11498),
            .DOUT(N__11497),
            .PACKAGEPIN(CPUCONFn));
    defparam CPUCONFn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUCONFn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CPUCONFn_ibuf_preio (
            .PADOEN(N__11499),
            .PADOUT(N__11498),
            .PADIN(N__11497),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CPUCONFn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RTC_ENn_obuf_iopad (
            .OE(N__11490),
            .DIN(N__11489),
            .DOUT(N__11488),
            .PACKAGEPIN(RTC_ENn));
    defparam RTC_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RTC_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RTC_ENn_obuf_preio (
            .PADOEN(N__11490),
            .PADOUT(N__11489),
            .PADIN(N__11488),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5237),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__11481),
            .DIN(N__11480),
            .DOUT(N__11479),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__11481),
            .PADOUT(N__11480),
            .PADIN(N__11479),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_4_iopad (
            .OE(N__11472),
            .DIN(N__11471),
            .DOUT(N__11470),
            .PACKAGEPIN(D[4]));
    defparam D_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_4_preio (
            .PADOEN(N__11472),
            .PADOUT(N__11471),
            .PADIN(N__11470),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5160),
            .DIN0(D_in_4),
            .DOUT0(N__5036),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11463),
            .DIN(N__11462),
            .DOUT(N__11461),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11463),
            .PADOUT(N__11462),
            .PADIN(N__11461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_1_iopad (
            .OE(N__11454),
            .DIN(N__11453),
            .DOUT(N__11452),
            .PACKAGEPIN(TM[1]));
    defparam TM_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_1_preio (
            .PADOEN(N__11454),
            .PADOUT(N__11453),
            .PADIN(N__11452),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__11445),
            .DIN(N__11444),
            .DOUT(N__11443),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__11445),
            .PADOUT(N__11444),
            .PADIN(N__11443),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_obuf_iopad (
            .OE(N__11436),
            .DIN(N__11435),
            .DOUT(N__11434),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMSPACEn_obuf_preio (
            .PADOEN(N__11436),
            .PADOUT(N__11435),
            .PADIN(N__11434),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8879),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11427),
            .DIN(N__11426),
            .DOUT(N__11425),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11427),
            .PADOUT(N__11426),
            .PADIN(N__11425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ROMENn_obuf_iopad (
            .OE(N__11418),
            .DIN(N__11417),
            .DOUT(N__11416),
            .PACKAGEPIN(ROMENn));
    defparam ROMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ROMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ROMENn_obuf_preio (
            .PADOEN(N__11418),
            .PADOUT(N__11417),
            .PADIN(N__11416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7304),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__11409),
            .DIN(N__11408),
            .DOUT(N__11407),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__11409),
            .PADOUT(N__11408),
            .PADIN(N__11407),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8969),
            .DIN0(),
            .DOUT0(N__7756),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11400),
            .DIN(N__11399),
            .DOUT(N__11398),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11400),
            .PADOUT(N__11399),
            .PADIN(N__11398),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__11391),
            .DIN(N__11390),
            .DOUT(N__11389),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__11391),
            .PADOUT(N__11390),
            .PADIN(N__11389),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6860),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_P2_obuf_iopad (
            .OE(N__11382),
            .DIN(N__11381),
            .DOUT(N__11380),
            .PACKAGEPIN(PIO_P2));
    defparam PIO_P2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_P2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_P2_obuf_preio (
            .PADOEN(N__11382),
            .PADOUT(N__11381),
            .PADIN(N__11380),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4175),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11373),
            .DIN(N__11372),
            .DOUT(N__11371),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11373),
            .PADOUT(N__11372),
            .PADIN(N__11371),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BRIDGE_ENn_obuf_iopad (
            .OE(N__11364),
            .DIN(N__11363),
            .DOUT(N__11362),
            .PACKAGEPIN(BRIDGE_ENn));
    defparam BRIDGE_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BRIDGE_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BRIDGE_ENn_obuf_preio (
            .PADOEN(N__11364),
            .PADOUT(N__11363),
            .PADIN(N__11362),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8276),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__11355),
            .DIN(N__11354),
            .DOUT(N__11353),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__11355),
            .PADOUT(N__11354),
            .PADIN(N__11353),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11346),
            .DIN(N__11345),
            .DOUT(N__11344),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11346),
            .PADOUT(N__11345),
            .PADIN(N__11344),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11337),
            .DIN(N__11336),
            .DOUT(N__11335),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11337),
            .PADOUT(N__11336),
            .PADIN(N__11335),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11328),
            .DIN(N__11327),
            .DOUT(N__11326),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11328),
            .PADOUT(N__11327),
            .PADIN(N__11326),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__11319),
            .DIN(N__11318),
            .DOUT(N__11317),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__11319),
            .PADOUT(N__11318),
            .PADIN(N__11317),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS0n_obuf_iopad (
            .OE(N__11310),
            .DIN(N__11309),
            .DOUT(N__11308),
            .PACKAGEPIN(CIACS0n));
    defparam CIACS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS0n_obuf_preio (
            .PADOEN(N__11310),
            .PADOUT(N__11309),
            .PADIN(N__11308),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10685),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__11301),
            .DIN(N__11300),
            .DOUT(N__11299),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__11301),
            .PADOUT(N__11300),
            .PADIN(N__11299),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7859),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11292),
            .DIN(N__11291),
            .DOUT(N__11290),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11292),
            .PADOUT(N__11291),
            .PADIN(N__11290),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__11283),
            .DIN(N__11282),
            .DOUT(N__11281),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__11283),
            .PADOUT(N__11282),
            .PADIN(N__11281),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__11274),
            .DIN(N__11273),
            .DOUT(N__11272),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__11274),
            .PADOUT(N__11273),
            .PADIN(N__11272),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__11265),
            .DIN(N__11264),
            .DOUT(N__11263),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__11265),
            .PADOUT(N__11264),
            .PADIN(N__11263),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__11256),
            .DIN(N__11255),
            .DOUT(N__11254),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__11256),
            .PADOUT(N__11255),
            .PADIN(N__11254),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8921),
            .DIN0(),
            .DOUT0(N__7757),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_5_iopad (
            .OE(N__11247),
            .DIN(N__11246),
            .DOUT(N__11245),
            .PACKAGEPIN(D[5]));
    defparam D_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_5_preio (
            .PADOEN(N__11247),
            .PADOUT(N__11246),
            .PADIN(N__11245),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5179),
            .DIN0(D_in_5),
            .DOUT0(N__5369),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__11238),
            .DIN(N__11237),
            .DOUT(N__11236),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__11238),
            .PADOUT(N__11237),
            .PADIN(N__11236),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11229),
            .DIN(N__11228),
            .DOUT(N__11227),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11229),
            .PADOUT(N__11228),
            .PADIN(N__11227),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11220),
            .DIN(N__11219),
            .DOUT(N__11218),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11220),
            .PADOUT(N__11219),
            .PADIN(N__11218),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CONFIGENn_obuf_iopad (
            .OE(N__11211),
            .DIN(N__11210),
            .DOUT(N__11209),
            .PACKAGEPIN(CONFIGENn));
    defparam CONFIGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CONFIGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CONFIGENn_obuf_preio (
            .PADOEN(N__11211),
            .PADOUT(N__11210),
            .PADIN(N__11209),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5681),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__11202),
            .DIN(N__11201),
            .DOUT(N__11200),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__11202),
            .PADOUT(N__11201),
            .PADIN(N__11200),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9365),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__11193),
            .DIN(N__11192),
            .DOUT(N__11191),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__11193),
            .PADOUT(N__11192),
            .PADIN(N__11191),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_P0_obuf_iopad (
            .OE(N__11184),
            .DIN(N__11183),
            .DOUT(N__11182),
            .PACKAGEPIN(PIO_P0));
    defparam PIO_P0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_P0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_P0_obuf_preio (
            .PADOEN(N__11184),
            .PADOUT(N__11183),
            .PADIN(N__11182),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10730),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__11175),
            .DIN(N__11174),
            .DOUT(N__11173),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__11175),
            .PADOUT(N__11174),
            .PADIN(N__11173),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__11166),
            .DIN(N__11165),
            .DOUT(N__11164),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__11166),
            .PADOUT(N__11165),
            .PADIN(N__11164),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ATA_ENn_obuf_iopad (
            .OE(N__11157),
            .DIN(N__11156),
            .DOUT(N__11155),
            .PACKAGEPIN(ATA_ENn));
    defparam ATA_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ATA_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ATA_ENn_obuf_preio (
            .PADOEN(N__11157),
            .PADOUT(N__11156),
            .PADIN(N__11155),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9197),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__11148),
            .DIN(N__11147),
            .DOUT(N__11146),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__11148),
            .PADOUT(N__11147),
            .PADIN(N__11146),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS1n_obuf_iopad (
            .OE(N__11139),
            .DIN(N__11138),
            .DOUT(N__11137),
            .PACKAGEPIN(CIACS1n));
    defparam CIACS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS1n_obuf_preio (
            .PADOEN(N__11139),
            .PADOUT(N__11138),
            .PADIN(N__11137),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10397),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_obuf_iopad (
            .OE(N__11130),
            .DIN(N__11129),
            .DOUT(N__11128),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGSPACEn_obuf_preio (
            .PADOEN(N__11130),
            .PADOUT(N__11129),
            .PADIN(N__11128),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4460),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__11121),
            .DIN(N__11120),
            .DOUT(N__11119),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__11121),
            .PADOUT(N__11120),
            .PADIN(N__11119),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_CIA_obuf_iopad (
            .OE(N__11112),
            .DIN(N__11111),
            .DOUT(N__11110),
            .PACKAGEPIN(CLK_CIA));
    defparam CLK_CIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_CIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_CIA_obuf_preio (
            .PADOEN(N__11112),
            .PADOUT(N__11111),
            .PADIN(N__11110),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10193),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__11103),
            .DIN(N__11102),
            .DOUT(N__11101),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__11103),
            .PADOUT(N__11102),
            .PADIN(N__11101),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__11094),
            .DIN(N__11093),
            .DOUT(N__11092),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__11094),
            .PADOUT(N__11093),
            .PADIN(N__11092),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8959),
            .DIN0(TACKn_in),
            .DOUT0(N__7749),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__11085),
            .DIN(N__11084),
            .DOUT(N__11083),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__11085),
            .PADOUT(N__11084),
            .PADIN(N__11083),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__11076),
            .DIN(N__11075),
            .DOUT(N__11074),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__11076),
            .PADOUT(N__11075),
            .PADIN(N__11074),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9011),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_S0_obuf_iopad (
            .OE(N__11067),
            .DIN(N__11066),
            .DOUT(N__11065),
            .PACKAGEPIN(PIO_S0));
    defparam PIO_S0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_S0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_S0_obuf_preio (
            .PADOEN(N__11067),
            .PADOUT(N__11066),
            .PADIN(N__11065),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4199),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__11058),
            .DIN(N__11057),
            .DOUT(N__11056),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__11058),
            .PADOUT(N__11057),
            .PADIN(N__11056),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_S2_obuf_iopad (
            .OE(N__11049),
            .DIN(N__11048),
            .DOUT(N__11047),
            .PACKAGEPIN(PIO_S2));
    defparam PIO_S2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_S2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_S2_obuf_preio (
            .PADOEN(N__11049),
            .PADOUT(N__11048),
            .PADIN(N__11047),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10462),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_6_iopad (
            .OE(N__11040),
            .DIN(N__11039),
            .DOUT(N__11038),
            .PACKAGEPIN(D[6]));
    defparam D_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_6_preio (
            .PADOEN(N__11040),
            .PADOUT(N__11039),
            .PADIN(N__11038),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5180),
            .DIN0(D_in_6),
            .DOUT0(N__5330),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11031),
            .DIN(N__11030),
            .DOUT(N__11029),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11031),
            .PADOUT(N__11030),
            .PADIN(N__11029),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__11022),
            .DIN(N__11021),
            .DOUT(N__11020),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__11022),
            .PADOUT(N__11021),
            .PADIN(N__11020),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PIO_S1_obuf_iopad (
            .OE(N__11013),
            .DIN(N__11012),
            .DOUT(N__11011),
            .PACKAGEPIN(PIO_S1));
    defparam PIO_S1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PIO_S1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PIO_S1_obuf_preio (
            .PADOEN(N__11013),
            .PADOUT(N__11012),
            .PADIN(N__11011),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4316),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_0_iopad (
            .OE(N__11004),
            .DIN(N__11003),
            .DOUT(N__11002),
            .PACKAGEPIN(TM[0]));
    defparam TM_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_0_preio (
            .PADOEN(N__11004),
            .PADOUT(N__11003),
            .PADIN(N__11002),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__10995),
            .DIN(N__10994),
            .DOUT(N__10993),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__10995),
            .PADOUT(N__10994),
            .PADIN(N__10993),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__10986),
            .DIN(N__10985),
            .DOUT(N__10984),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__10986),
            .PADOUT(N__10985),
            .PADIN(N__10984),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2644 (
            .O(N__10967),
            .I(N__10964));
    LocalMux I__2643 (
            .O(N__10964),
            .I(N__10960));
    InMux I__2642 (
            .O(N__10963),
            .I(N__10957));
    Span4Mux_v I__2641 (
            .O(N__10960),
            .I(N__10954));
    LocalMux I__2640 (
            .O(N__10957),
            .I(N__10951));
    Sp12to4 I__2639 (
            .O(N__10954),
            .I(N__10947));
    Span4Mux_v I__2638 (
            .O(N__10951),
            .I(N__10944));
    InMux I__2637 (
            .O(N__10950),
            .I(N__10941));
    Odrv12 I__2636 (
            .O(N__10947),
            .I(\U409_CIA.VMAZ0 ));
    Odrv4 I__2635 (
            .O(N__10944),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__2634 (
            .O(N__10941),
            .I(\U409_CIA.VMAZ0 ));
    CascadeMux I__2633 (
            .O(N__10934),
            .I(N__10930));
    InMux I__2632 (
            .O(N__10933),
            .I(N__10926));
    InMux I__2631 (
            .O(N__10930),
            .I(N__10923));
    CascadeMux I__2630 (
            .O(N__10929),
            .I(N__10920));
    LocalMux I__2629 (
            .O(N__10926),
            .I(N__10908));
    LocalMux I__2628 (
            .O(N__10923),
            .I(N__10908));
    InMux I__2627 (
            .O(N__10920),
            .I(N__10905));
    InMux I__2626 (
            .O(N__10919),
            .I(N__10900));
    InMux I__2625 (
            .O(N__10918),
            .I(N__10900));
    InMux I__2624 (
            .O(N__10917),
            .I(N__10897));
    CascadeMux I__2623 (
            .O(N__10916),
            .I(N__10894));
    CascadeMux I__2622 (
            .O(N__10915),
            .I(N__10890));
    CascadeMux I__2621 (
            .O(N__10914),
            .I(N__10885));
    CascadeMux I__2620 (
            .O(N__10913),
            .I(N__10881));
    Span4Mux_v I__2619 (
            .O(N__10908),
            .I(N__10872));
    LocalMux I__2618 (
            .O(N__10905),
            .I(N__10872));
    LocalMux I__2617 (
            .O(N__10900),
            .I(N__10872));
    LocalMux I__2616 (
            .O(N__10897),
            .I(N__10868));
    InMux I__2615 (
            .O(N__10894),
            .I(N__10859));
    InMux I__2614 (
            .O(N__10893),
            .I(N__10859));
    InMux I__2613 (
            .O(N__10890),
            .I(N__10859));
    InMux I__2612 (
            .O(N__10889),
            .I(N__10859));
    InMux I__2611 (
            .O(N__10888),
            .I(N__10856));
    InMux I__2610 (
            .O(N__10885),
            .I(N__10853));
    InMux I__2609 (
            .O(N__10884),
            .I(N__10850));
    InMux I__2608 (
            .O(N__10881),
            .I(N__10847));
    InMux I__2607 (
            .O(N__10880),
            .I(N__10842));
    InMux I__2606 (
            .O(N__10879),
            .I(N__10842));
    Span4Mux_v I__2605 (
            .O(N__10872),
            .I(N__10839));
    InMux I__2604 (
            .O(N__10871),
            .I(N__10836));
    Span4Mux_h I__2603 (
            .O(N__10868),
            .I(N__10827));
    LocalMux I__2602 (
            .O(N__10859),
            .I(N__10827));
    LocalMux I__2601 (
            .O(N__10856),
            .I(N__10827));
    LocalMux I__2600 (
            .O(N__10853),
            .I(N__10827));
    LocalMux I__2599 (
            .O(N__10850),
            .I(N__10818));
    LocalMux I__2598 (
            .O(N__10847),
            .I(N__10818));
    LocalMux I__2597 (
            .O(N__10842),
            .I(N__10818));
    Span4Mux_h I__2596 (
            .O(N__10839),
            .I(N__10811));
    LocalMux I__2595 (
            .O(N__10836),
            .I(N__10811));
    Span4Mux_v I__2594 (
            .O(N__10827),
            .I(N__10808));
    InMux I__2593 (
            .O(N__10826),
            .I(N__10805));
    InMux I__2592 (
            .O(N__10825),
            .I(N__10802));
    Span4Mux_v I__2591 (
            .O(N__10818),
            .I(N__10799));
    InMux I__2590 (
            .O(N__10817),
            .I(N__10794));
    InMux I__2589 (
            .O(N__10816),
            .I(N__10794));
    Span4Mux_v I__2588 (
            .O(N__10811),
            .I(N__10790));
    Span4Mux_h I__2587 (
            .O(N__10808),
            .I(N__10787));
    LocalMux I__2586 (
            .O(N__10805),
            .I(N__10782));
    LocalMux I__2585 (
            .O(N__10802),
            .I(N__10782));
    Span4Mux_v I__2584 (
            .O(N__10799),
            .I(N__10777));
    LocalMux I__2583 (
            .O(N__10794),
            .I(N__10777));
    InMux I__2582 (
            .O(N__10793),
            .I(N__10774));
    Sp12to4 I__2581 (
            .O(N__10790),
            .I(N__10770));
    Sp12to4 I__2580 (
            .O(N__10787),
            .I(N__10761));
    Span12Mux_v I__2579 (
            .O(N__10782),
            .I(N__10761));
    Sp12to4 I__2578 (
            .O(N__10777),
            .I(N__10761));
    LocalMux I__2577 (
            .O(N__10774),
            .I(N__10761));
    InMux I__2576 (
            .O(N__10773),
            .I(N__10758));
    Span12Mux_h I__2575 (
            .O(N__10770),
            .I(N__10755));
    Span12Mux_v I__2574 (
            .O(N__10761),
            .I(N__10752));
    LocalMux I__2573 (
            .O(N__10758),
            .I(N__10749));
    Span12Mux_v I__2572 (
            .O(N__10755),
            .I(N__10746));
    Span12Mux_h I__2571 (
            .O(N__10752),
            .I(N__10741));
    Span12Mux_v I__2570 (
            .O(N__10749),
            .I(N__10741));
    Odrv12 I__2569 (
            .O(N__10746),
            .I(RESETn_c));
    Odrv12 I__2568 (
            .O(N__10741),
            .I(RESETn_c));
    InMux I__2567 (
            .O(N__10736),
            .I(N__10733));
    LocalMux I__2566 (
            .O(N__10733),
            .I(CIA_ENABLE));
    IoInMux I__2565 (
            .O(N__10730),
            .I(N__10727));
    LocalMux I__2564 (
            .O(N__10727),
            .I(N__10724));
    Span4Mux_s0_h I__2563 (
            .O(N__10724),
            .I(N__10720));
    InMux I__2562 (
            .O(N__10723),
            .I(N__10717));
    Sp12to4 I__2561 (
            .O(N__10720),
            .I(N__10714));
    LocalMux I__2560 (
            .O(N__10717),
            .I(N__10711));
    Span12Mux_s10_v I__2559 (
            .O(N__10714),
            .I(N__10708));
    Span12Mux_s10_v I__2558 (
            .O(N__10711),
            .I(N__10705));
    Span12Mux_h I__2557 (
            .O(N__10708),
            .I(N__10702));
    Span12Mux_h I__2556 (
            .O(N__10705),
            .I(N__10699));
    Span12Mux_h I__2555 (
            .O(N__10702),
            .I(N__10696));
    Span12Mux_h I__2554 (
            .O(N__10699),
            .I(N__10693));
    Odrv12 I__2553 (
            .O(N__10696),
            .I(A_c_12));
    Odrv12 I__2552 (
            .O(N__10693),
            .I(A_c_12));
    CascadeMux I__2551 (
            .O(N__10688),
            .I(CIA_ENABLE_cascade_));
    IoInMux I__2550 (
            .O(N__10685),
            .I(N__10682));
    LocalMux I__2549 (
            .O(N__10682),
            .I(N__10679));
    Span4Mux_s3_h I__2548 (
            .O(N__10679),
            .I(N__10676));
    Span4Mux_v I__2547 (
            .O(N__10676),
            .I(N__10673));
    Odrv4 I__2546 (
            .O(N__10673),
            .I(U409_ADDRESS_DECODE_un1_CIACS0n_i));
    InMux I__2545 (
            .O(N__10670),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__2544 (
            .O(N__10667),
            .I(N__10663));
    InMux I__2543 (
            .O(N__10666),
            .I(N__10660));
    LocalMux I__2542 (
            .O(N__10663),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__2541 (
            .O(N__10660),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    InMux I__2540 (
            .O(N__10655),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__2539 (
            .O(N__10652),
            .I(N__10648));
    InMux I__2538 (
            .O(N__10651),
            .I(N__10645));
    LocalMux I__2537 (
            .O(N__10648),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__2536 (
            .O(N__10645),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__2535 (
            .O(N__10640),
            .I(N__10637));
    LocalMux I__2534 (
            .O(N__10637),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__2533 (
            .O(N__10634),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__2532 (
            .O(N__10631),
            .I(N__10627));
    InMux I__2531 (
            .O(N__10630),
            .I(N__10624));
    LocalMux I__2530 (
            .O(N__10627),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__2529 (
            .O(N__10624),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    InMux I__2528 (
            .O(N__10619),
            .I(N__10616));
    LocalMux I__2527 (
            .O(N__10616),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__2526 (
            .O(N__10613),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__2525 (
            .O(N__10610),
            .I(N__10606));
    InMux I__2524 (
            .O(N__10609),
            .I(N__10603));
    LocalMux I__2523 (
            .O(N__10606),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__2522 (
            .O(N__10603),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    CascadeMux I__2521 (
            .O(N__10598),
            .I(N__10595));
    InMux I__2520 (
            .O(N__10595),
            .I(N__10592));
    LocalMux I__2519 (
            .O(N__10592),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__2518 (
            .O(N__10589),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__2517 (
            .O(N__10586),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__2516 (
            .O(N__10583),
            .I(N__10579));
    InMux I__2515 (
            .O(N__10582),
            .I(N__10576));
    LocalMux I__2514 (
            .O(N__10579),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__2513 (
            .O(N__10576),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    ClkMux I__2512 (
            .O(N__10571),
            .I(N__10544));
    ClkMux I__2511 (
            .O(N__10570),
            .I(N__10544));
    ClkMux I__2510 (
            .O(N__10569),
            .I(N__10544));
    ClkMux I__2509 (
            .O(N__10568),
            .I(N__10544));
    ClkMux I__2508 (
            .O(N__10567),
            .I(N__10544));
    ClkMux I__2507 (
            .O(N__10566),
            .I(N__10544));
    ClkMux I__2506 (
            .O(N__10565),
            .I(N__10544));
    ClkMux I__2505 (
            .O(N__10564),
            .I(N__10544));
    ClkMux I__2504 (
            .O(N__10563),
            .I(N__10544));
    GlobalMux I__2503 (
            .O(N__10544),
            .I(N__10541));
    gio2CtrlBuf I__2502 (
            .O(N__10541),
            .I(CLK6_c_g));
    InMux I__2501 (
            .O(N__10538),
            .I(N__10532));
    InMux I__2500 (
            .O(N__10537),
            .I(N__10529));
    InMux I__2499 (
            .O(N__10536),
            .I(N__10526));
    InMux I__2498 (
            .O(N__10535),
            .I(N__10523));
    LocalMux I__2497 (
            .O(N__10532),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__2496 (
            .O(N__10529),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__2495 (
            .O(N__10526),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__2494 (
            .O(N__10523),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    CascadeMux I__2493 (
            .O(N__10514),
            .I(N__10511));
    InMux I__2492 (
            .O(N__10511),
            .I(N__10506));
    InMux I__2491 (
            .O(N__10510),
            .I(N__10498));
    InMux I__2490 (
            .O(N__10509),
            .I(N__10498));
    LocalMux I__2489 (
            .O(N__10506),
            .I(N__10495));
    InMux I__2488 (
            .O(N__10505),
            .I(N__10492));
    InMux I__2487 (
            .O(N__10504),
            .I(N__10487));
    InMux I__2486 (
            .O(N__10503),
            .I(N__10487));
    LocalMux I__2485 (
            .O(N__10498),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    Odrv4 I__2484 (
            .O(N__10495),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__2483 (
            .O(N__10492),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__2482 (
            .O(N__10487),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    InMux I__2481 (
            .O(N__10478),
            .I(N__10474));
    InMux I__2480 (
            .O(N__10477),
            .I(N__10471));
    LocalMux I__2479 (
            .O(N__10474),
            .I(\U409_CIA.CIA_CLK_COUNT11_2 ));
    LocalMux I__2478 (
            .O(N__10471),
            .I(\U409_CIA.CIA_CLK_COUNT11_2 ));
    IoInMux I__2477 (
            .O(N__10466),
            .I(N__10463));
    LocalMux I__2476 (
            .O(N__10463),
            .I(N__10459));
    IoInMux I__2475 (
            .O(N__10462),
            .I(N__10456));
    Span4Mux_s0_v I__2474 (
            .O(N__10459),
            .I(N__10453));
    LocalMux I__2473 (
            .O(N__10456),
            .I(N__10450));
    Sp12to4 I__2472 (
            .O(N__10453),
            .I(N__10447));
    Span4Mux_s3_h I__2471 (
            .O(N__10450),
            .I(N__10444));
    Span12Mux_h I__2470 (
            .O(N__10447),
            .I(N__10441));
    Span4Mux_v I__2469 (
            .O(N__10444),
            .I(N__10438));
    Odrv12 I__2468 (
            .O(N__10441),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2467 (
            .O(N__10438),
            .I(CONSTANT_ONE_NET));
    IoInMux I__2466 (
            .O(N__10433),
            .I(N__10430));
    LocalMux I__2465 (
            .O(N__10430),
            .I(N__10427));
    IoSpan4Mux I__2464 (
            .O(N__10427),
            .I(N__10423));
    InMux I__2463 (
            .O(N__10426),
            .I(N__10420));
    IoSpan4Mux I__2462 (
            .O(N__10423),
            .I(N__10417));
    LocalMux I__2461 (
            .O(N__10420),
            .I(N__10414));
    Span4Mux_s3_h I__2460 (
            .O(N__10417),
            .I(N__10409));
    Span4Mux_v I__2459 (
            .O(N__10414),
            .I(N__10409));
    Sp12to4 I__2458 (
            .O(N__10409),
            .I(N__10406));
    Span12Mux_h I__2457 (
            .O(N__10406),
            .I(N__10403));
    Span12Mux_h I__2456 (
            .O(N__10403),
            .I(N__10400));
    Odrv12 I__2455 (
            .O(N__10400),
            .I(A_c_13));
    IoInMux I__2454 (
            .O(N__10397),
            .I(N__10394));
    LocalMux I__2453 (
            .O(N__10394),
            .I(N__10391));
    Span4Mux_s3_h I__2452 (
            .O(N__10391),
            .I(N__10388));
    Span4Mux_v I__2451 (
            .O(N__10388),
            .I(N__10385));
    Odrv4 I__2450 (
            .O(N__10385),
            .I(U409_ADDRESS_DECODE_un1_CIACS1n_i));
    InMux I__2449 (
            .O(N__10382),
            .I(N__10378));
    InMux I__2448 (
            .O(N__10381),
            .I(N__10375));
    LocalMux I__2447 (
            .O(N__10378),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__2446 (
            .O(N__10375),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__2445 (
            .O(N__10370),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    CascadeMux I__2444 (
            .O(N__10367),
            .I(N__10364));
    InMux I__2443 (
            .O(N__10364),
            .I(N__10360));
    InMux I__2442 (
            .O(N__10363),
            .I(N__10357));
    LocalMux I__2441 (
            .O(N__10360),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__2440 (
            .O(N__10357),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    InMux I__2439 (
            .O(N__10352),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__2438 (
            .O(N__10349),
            .I(N__10345));
    InMux I__2437 (
            .O(N__10348),
            .I(N__10342));
    LocalMux I__2436 (
            .O(N__10345),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__2435 (
            .O(N__10342),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__2434 (
            .O(N__10337),
            .I(N__10334));
    LocalMux I__2433 (
            .O(N__10334),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__2432 (
            .O(N__10331),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    InMux I__2431 (
            .O(N__10328),
            .I(N__10324));
    InMux I__2430 (
            .O(N__10327),
            .I(N__10321));
    LocalMux I__2429 (
            .O(N__10324),
            .I(N__10318));
    LocalMux I__2428 (
            .O(N__10321),
            .I(N__10315));
    Odrv4 I__2427 (
            .O(N__10318),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    Odrv4 I__2426 (
            .O(N__10315),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    InMux I__2425 (
            .O(N__10310),
            .I(N__10307));
    LocalMux I__2424 (
            .O(N__10307),
            .I(N__10304));
    Odrv4 I__2423 (
            .O(N__10304),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__2422 (
            .O(N__10301),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__2421 (
            .O(N__10298),
            .I(N__10294));
    InMux I__2420 (
            .O(N__10297),
            .I(N__10291));
    LocalMux I__2419 (
            .O(N__10294),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__2418 (
            .O(N__10291),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    InMux I__2417 (
            .O(N__10286),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__2416 (
            .O(N__10283),
            .I(N__10279));
    InMux I__2415 (
            .O(N__10282),
            .I(N__10276));
    LocalMux I__2414 (
            .O(N__10279),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__2413 (
            .O(N__10276),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__2412 (
            .O(N__10271),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    CascadeMux I__2411 (
            .O(N__10268),
            .I(N__10265));
    InMux I__2410 (
            .O(N__10265),
            .I(N__10261));
    InMux I__2409 (
            .O(N__10264),
            .I(N__10258));
    LocalMux I__2408 (
            .O(N__10261),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__2407 (
            .O(N__10258),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    CascadeMux I__2406 (
            .O(N__10253),
            .I(N__10250));
    InMux I__2405 (
            .O(N__10250),
            .I(N__10247));
    LocalMux I__2404 (
            .O(N__10247),
            .I(N__10244));
    Odrv12 I__2403 (
            .O(N__10244),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__2402 (
            .O(N__10241),
            .I(bfn_15_7_0_));
    InMux I__2401 (
            .O(N__10238),
            .I(N__10234));
    InMux I__2400 (
            .O(N__10237),
            .I(N__10231));
    LocalMux I__2399 (
            .O(N__10234),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__2398 (
            .O(N__10231),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    InMux I__2397 (
            .O(N__10226),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__2396 (
            .O(N__10223),
            .I(N__10220));
    LocalMux I__2395 (
            .O(N__10220),
            .I(N__10216));
    InMux I__2394 (
            .O(N__10219),
            .I(N__10213));
    Odrv4 I__2393 (
            .O(N__10216),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__2392 (
            .O(N__10213),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__2391 (
            .O(N__10208),
            .I(N__10205));
    LocalMux I__2390 (
            .O(N__10205),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__2389 (
            .O(N__10202),
            .I(N__10199));
    LocalMux I__2388 (
            .O(N__10199),
            .I(\U409_CIA.CLK_CIA_r_1_0 ));
    CascadeMux I__2387 (
            .O(N__10196),
            .I(\U409_CIA.CLK_CIA6_3_cascade_ ));
    IoInMux I__2386 (
            .O(N__10193),
            .I(N__10190));
    LocalMux I__2385 (
            .O(N__10190),
            .I(N__10187));
    IoSpan4Mux I__2384 (
            .O(N__10187),
            .I(N__10184));
    Span4Mux_s3_v I__2383 (
            .O(N__10184),
            .I(N__10181));
    Sp12to4 I__2382 (
            .O(N__10181),
            .I(N__10176));
    InMux I__2381 (
            .O(N__10180),
            .I(N__10173));
    CascadeMux I__2380 (
            .O(N__10179),
            .I(N__10169));
    Span12Mux_s10_v I__2379 (
            .O(N__10176),
            .I(N__10166));
    LocalMux I__2378 (
            .O(N__10173),
            .I(N__10163));
    InMux I__2377 (
            .O(N__10172),
            .I(N__10160));
    InMux I__2376 (
            .O(N__10169),
            .I(N__10157));
    Odrv12 I__2375 (
            .O(N__10166),
            .I(CLK_CIA_c));
    Odrv12 I__2374 (
            .O(N__10163),
            .I(CLK_CIA_c));
    LocalMux I__2373 (
            .O(N__10160),
            .I(CLK_CIA_c));
    LocalMux I__2372 (
            .O(N__10157),
            .I(CLK_CIA_c));
    InMux I__2371 (
            .O(N__10148),
            .I(N__10140));
    InMux I__2370 (
            .O(N__10147),
            .I(N__10140));
    InMux I__2369 (
            .O(N__10146),
            .I(N__10137));
    InMux I__2368 (
            .O(N__10145),
            .I(N__10134));
    LocalMux I__2367 (
            .O(N__10140),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__2366 (
            .O(N__10137),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__2365 (
            .O(N__10134),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    CascadeMux I__2364 (
            .O(N__10127),
            .I(N__10119));
    InMux I__2363 (
            .O(N__10126),
            .I(N__10116));
    InMux I__2362 (
            .O(N__10125),
            .I(N__10109));
    InMux I__2361 (
            .O(N__10124),
            .I(N__10109));
    InMux I__2360 (
            .O(N__10123),
            .I(N__10109));
    InMux I__2359 (
            .O(N__10122),
            .I(N__10104));
    InMux I__2358 (
            .O(N__10119),
            .I(N__10104));
    LocalMux I__2357 (
            .O(N__10116),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__2356 (
            .O(N__10109),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__2355 (
            .O(N__10104),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    CascadeMux I__2354 (
            .O(N__10097),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ));
    InMux I__2353 (
            .O(N__10094),
            .I(N__10091));
    LocalMux I__2352 (
            .O(N__10091),
            .I(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5 ));
    CascadeMux I__2351 (
            .O(N__10088),
            .I(N__10083));
    CascadeMux I__2350 (
            .O(N__10087),
            .I(N__10079));
    InMux I__2349 (
            .O(N__10086),
            .I(N__10074));
    InMux I__2348 (
            .O(N__10083),
            .I(N__10074));
    InMux I__2347 (
            .O(N__10082),
            .I(N__10071));
    InMux I__2346 (
            .O(N__10079),
            .I(N__10068));
    LocalMux I__2345 (
            .O(N__10074),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__2344 (
            .O(N__10071),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__2343 (
            .O(N__10068),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    InMux I__2342 (
            .O(N__10061),
            .I(N__10056));
    InMux I__2341 (
            .O(N__10060),
            .I(N__10051));
    InMux I__2340 (
            .O(N__10059),
            .I(N__10051));
    LocalMux I__2339 (
            .O(N__10056),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__2338 (
            .O(N__10051),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    InMux I__2337 (
            .O(N__10046),
            .I(N__10041));
    InMux I__2336 (
            .O(N__10045),
            .I(N__10038));
    InMux I__2335 (
            .O(N__10044),
            .I(N__10035));
    LocalMux I__2334 (
            .O(N__10041),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__2333 (
            .O(N__10038),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__2332 (
            .O(N__10035),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    InMux I__2331 (
            .O(N__10028),
            .I(N__10024));
    InMux I__2330 (
            .O(N__10027),
            .I(N__10021));
    LocalMux I__2329 (
            .O(N__10024),
            .I(\U409_CIA.CLK_CIA6_4 ));
    LocalMux I__2328 (
            .O(N__10021),
            .I(\U409_CIA.CLK_CIA6_4 ));
    InMux I__2327 (
            .O(N__10016),
            .I(N__10013));
    LocalMux I__2326 (
            .O(N__10013),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0 ));
    CascadeMux I__2325 (
            .O(N__10010),
            .I(\U409_CIA.CLK_CIA6_4_cascade_ ));
    InMux I__2324 (
            .O(N__10007),
            .I(N__10004));
    LocalMux I__2323 (
            .O(N__10004),
            .I(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3 ));
    InMux I__2322 (
            .O(N__10001),
            .I(N__9993));
    InMux I__2321 (
            .O(N__10000),
            .I(N__9993));
    InMux I__2320 (
            .O(N__9999),
            .I(N__9990));
    InMux I__2319 (
            .O(N__9998),
            .I(N__9987));
    LocalMux I__2318 (
            .O(N__9993),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__2317 (
            .O(N__9990),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__2316 (
            .O(N__9987),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    ClkMux I__2315 (
            .O(N__9980),
            .I(N__9971));
    ClkMux I__2314 (
            .O(N__9979),
            .I(N__9971));
    ClkMux I__2313 (
            .O(N__9978),
            .I(N__9971));
    GlobalMux I__2312 (
            .O(N__9971),
            .I(N__9968));
    gio2CtrlBuf I__2311 (
            .O(N__9968),
            .I(CLK28_IN_c_g));
    CascadeMux I__2310 (
            .O(N__9965),
            .I(N__9961));
    InMux I__2309 (
            .O(N__9964),
            .I(N__9955));
    InMux I__2308 (
            .O(N__9961),
            .I(N__9955));
    InMux I__2307 (
            .O(N__9960),
            .I(N__9952));
    LocalMux I__2306 (
            .O(N__9955),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__2305 (
            .O(N__9952),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    CascadeMux I__2304 (
            .O(N__9947),
            .I(N__9941));
    InMux I__2303 (
            .O(N__9946),
            .I(N__9936));
    InMux I__2302 (
            .O(N__9945),
            .I(N__9936));
    InMux I__2301 (
            .O(N__9944),
            .I(N__9933));
    InMux I__2300 (
            .O(N__9941),
            .I(N__9930));
    LocalMux I__2299 (
            .O(N__9936),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2298 (
            .O(N__9933),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2297 (
            .O(N__9930),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__2296 (
            .O(N__9923),
            .I(N__9919));
    InMux I__2295 (
            .O(N__9922),
            .I(N__9916));
    LocalMux I__2294 (
            .O(N__9919),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__2293 (
            .O(N__9916),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__2292 (
            .O(N__9911),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__2291 (
            .O(N__9908),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__2290 (
            .O(N__9905),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__2289 (
            .O(N__9902),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__2288 (
            .O(N__9899),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    InMux I__2287 (
            .O(N__9896),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ));
    InMux I__2286 (
            .O(N__9893),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ));
    InMux I__2285 (
            .O(N__9890),
            .I(N__9887));
    LocalMux I__2284 (
            .O(N__9887),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__2283 (
            .O(N__9884),
            .I(N__9879));
    InMux I__2282 (
            .O(N__9883),
            .I(N__9876));
    InMux I__2281 (
            .O(N__9882),
            .I(N__9873));
    LocalMux I__2280 (
            .O(N__9879),
            .I(N__9865));
    LocalMux I__2279 (
            .O(N__9876),
            .I(N__9862));
    LocalMux I__2278 (
            .O(N__9873),
            .I(N__9859));
    InMux I__2277 (
            .O(N__9872),
            .I(N__9854));
    InMux I__2276 (
            .O(N__9871),
            .I(N__9854));
    InMux I__2275 (
            .O(N__9870),
            .I(N__9847));
    InMux I__2274 (
            .O(N__9869),
            .I(N__9847));
    InMux I__2273 (
            .O(N__9868),
            .I(N__9847));
    Odrv4 I__2272 (
            .O(N__9865),
            .I(\U409_TICK.TICK503_14 ));
    Odrv4 I__2271 (
            .O(N__9862),
            .I(\U409_TICK.TICK503_14 ));
    Odrv4 I__2270 (
            .O(N__9859),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__2269 (
            .O(N__9854),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__2268 (
            .O(N__9847),
            .I(\U409_TICK.TICK503_14 ));
    InMux I__2267 (
            .O(N__9836),
            .I(N__9833));
    LocalMux I__2266 (
            .O(N__9833),
            .I(N__9827));
    InMux I__2265 (
            .O(N__9832),
            .I(N__9824));
    InMux I__2264 (
            .O(N__9831),
            .I(N__9819));
    InMux I__2263 (
            .O(N__9830),
            .I(N__9819));
    Span4Mux_h I__2262 (
            .O(N__9827),
            .I(N__9811));
    LocalMux I__2261 (
            .O(N__9824),
            .I(N__9806));
    LocalMux I__2260 (
            .O(N__9819),
            .I(N__9806));
    InMux I__2259 (
            .O(N__9818),
            .I(N__9803));
    InMux I__2258 (
            .O(N__9817),
            .I(N__9800));
    InMux I__2257 (
            .O(N__9816),
            .I(N__9793));
    InMux I__2256 (
            .O(N__9815),
            .I(N__9793));
    InMux I__2255 (
            .O(N__9814),
            .I(N__9793));
    Odrv4 I__2254 (
            .O(N__9811),
            .I(\U409_TICK.TICK503_10 ));
    Odrv12 I__2253 (
            .O(N__9806),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__2252 (
            .O(N__9803),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__2251 (
            .O(N__9800),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__2250 (
            .O(N__9793),
            .I(\U409_TICK.TICK503_10 ));
    CascadeMux I__2249 (
            .O(N__9782),
            .I(N__9778));
    CascadeMux I__2248 (
            .O(N__9781),
            .I(N__9772));
    InMux I__2247 (
            .O(N__9778),
            .I(N__9769));
    CascadeMux I__2246 (
            .O(N__9777),
            .I(N__9766));
    CascadeMux I__2245 (
            .O(N__9776),
            .I(N__9762));
    CascadeMux I__2244 (
            .O(N__9775),
            .I(N__9757));
    InMux I__2243 (
            .O(N__9772),
            .I(N__9754));
    LocalMux I__2242 (
            .O(N__9769),
            .I(N__9751));
    InMux I__2241 (
            .O(N__9766),
            .I(N__9748));
    InMux I__2240 (
            .O(N__9765),
            .I(N__9743));
    InMux I__2239 (
            .O(N__9762),
            .I(N__9743));
    InMux I__2238 (
            .O(N__9761),
            .I(N__9736));
    InMux I__2237 (
            .O(N__9760),
            .I(N__9736));
    InMux I__2236 (
            .O(N__9757),
            .I(N__9736));
    LocalMux I__2235 (
            .O(N__9754),
            .I(N__9733));
    Span4Mux_v I__2234 (
            .O(N__9751),
            .I(N__9728));
    LocalMux I__2233 (
            .O(N__9748),
            .I(N__9728));
    LocalMux I__2232 (
            .O(N__9743),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__2231 (
            .O(N__9736),
            .I(\U409_TICK.TICK503_9 ));
    Odrv4 I__2230 (
            .O(N__9733),
            .I(\U409_TICK.TICK503_9 ));
    Odrv4 I__2229 (
            .O(N__9728),
            .I(\U409_TICK.TICK503_9 ));
    InMux I__2228 (
            .O(N__9719),
            .I(N__9715));
    InMux I__2227 (
            .O(N__9718),
            .I(N__9712));
    LocalMux I__2226 (
            .O(N__9715),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__2225 (
            .O(N__9712),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    CascadeMux I__2224 (
            .O(N__9707),
            .I(N__9703));
    InMux I__2223 (
            .O(N__9706),
            .I(N__9700));
    InMux I__2222 (
            .O(N__9703),
            .I(N__9697));
    LocalMux I__2221 (
            .O(N__9700),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__2220 (
            .O(N__9697),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    CascadeMux I__2219 (
            .O(N__9692),
            .I(N__9689));
    InMux I__2218 (
            .O(N__9689),
            .I(N__9685));
    InMux I__2217 (
            .O(N__9688),
            .I(N__9682));
    LocalMux I__2216 (
            .O(N__9685),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__2215 (
            .O(N__9682),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    InMux I__2214 (
            .O(N__9677),
            .I(N__9674));
    LocalMux I__2213 (
            .O(N__9674),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    CascadeMux I__2212 (
            .O(N__9671),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    CascadeMux I__2211 (
            .O(N__9668),
            .I(N__9664));
    InMux I__2210 (
            .O(N__9667),
            .I(N__9661));
    InMux I__2209 (
            .O(N__9664),
            .I(N__9658));
    LocalMux I__2208 (
            .O(N__9661),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__2207 (
            .O(N__9658),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__2206 (
            .O(N__9653),
            .I(N__9650));
    LocalMux I__2205 (
            .O(N__9650),
            .I(N__9646));
    InMux I__2204 (
            .O(N__9649),
            .I(N__9643));
    Odrv4 I__2203 (
            .O(N__9646),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__2202 (
            .O(N__9643),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    CascadeMux I__2201 (
            .O(N__9638),
            .I(N__9633));
    CascadeMux I__2200 (
            .O(N__9637),
            .I(N__9630));
    CascadeMux I__2199 (
            .O(N__9636),
            .I(N__9626));
    InMux I__2198 (
            .O(N__9633),
            .I(N__9621));
    InMux I__2197 (
            .O(N__9630),
            .I(N__9621));
    InMux I__2196 (
            .O(N__9629),
            .I(N__9618));
    InMux I__2195 (
            .O(N__9626),
            .I(N__9615));
    LocalMux I__2194 (
            .O(N__9621),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__2193 (
            .O(N__9618),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__2192 (
            .O(N__9615),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__2191 (
            .O(N__9608),
            .I(N__9604));
    InMux I__2190 (
            .O(N__9607),
            .I(N__9601));
    LocalMux I__2189 (
            .O(N__9604),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__2188 (
            .O(N__9601),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__2187 (
            .O(N__9596),
            .I(N__9593));
    LocalMux I__2186 (
            .O(N__9593),
            .I(\U409_TICK.TICK603_11 ));
    InMux I__2185 (
            .O(N__9590),
            .I(N__9586));
    InMux I__2184 (
            .O(N__9589),
            .I(N__9583));
    LocalMux I__2183 (
            .O(N__9586),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__2182 (
            .O(N__9583),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    CascadeMux I__2181 (
            .O(N__9578),
            .I(\U409_TICK.TICK603_8_cascade_ ));
    InMux I__2180 (
            .O(N__9575),
            .I(N__9572));
    LocalMux I__2179 (
            .O(N__9572),
            .I(N__9568));
    InMux I__2178 (
            .O(N__9571),
            .I(N__9565));
    Odrv4 I__2177 (
            .O(N__9568),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__2176 (
            .O(N__9565),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    CascadeMux I__2175 (
            .O(N__9560),
            .I(N__9557));
    InMux I__2174 (
            .O(N__9557),
            .I(N__9548));
    InMux I__2173 (
            .O(N__9556),
            .I(N__9539));
    InMux I__2172 (
            .O(N__9555),
            .I(N__9539));
    InMux I__2171 (
            .O(N__9554),
            .I(N__9539));
    InMux I__2170 (
            .O(N__9553),
            .I(N__9539));
    InMux I__2169 (
            .O(N__9552),
            .I(N__9534));
    InMux I__2168 (
            .O(N__9551),
            .I(N__9534));
    LocalMux I__2167 (
            .O(N__9548),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__2166 (
            .O(N__9539),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__2165 (
            .O(N__9534),
            .I(\U409_TICK.TICK603_14 ));
    CascadeMux I__2164 (
            .O(N__9527),
            .I(N__9519));
    InMux I__2163 (
            .O(N__9526),
            .I(N__9508));
    InMux I__2162 (
            .O(N__9525),
            .I(N__9508));
    InMux I__2161 (
            .O(N__9524),
            .I(N__9508));
    InMux I__2160 (
            .O(N__9523),
            .I(N__9508));
    InMux I__2159 (
            .O(N__9522),
            .I(N__9499));
    InMux I__2158 (
            .O(N__9519),
            .I(N__9499));
    InMux I__2157 (
            .O(N__9518),
            .I(N__9499));
    InMux I__2156 (
            .O(N__9517),
            .I(N__9499));
    LocalMux I__2155 (
            .O(N__9508),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__2154 (
            .O(N__9499),
            .I(\U409_TICK.TICK603_10 ));
    CascadeMux I__2153 (
            .O(N__9494),
            .I(N__9489));
    CascadeMux I__2152 (
            .O(N__9493),
            .I(N__9486));
    CascadeMux I__2151 (
            .O(N__9492),
            .I(N__9483));
    InMux I__2150 (
            .O(N__9489),
            .I(N__9470));
    InMux I__2149 (
            .O(N__9486),
            .I(N__9470));
    InMux I__2148 (
            .O(N__9483),
            .I(N__9470));
    InMux I__2147 (
            .O(N__9482),
            .I(N__9470));
    InMux I__2146 (
            .O(N__9481),
            .I(N__9463));
    InMux I__2145 (
            .O(N__9480),
            .I(N__9463));
    InMux I__2144 (
            .O(N__9479),
            .I(N__9463));
    LocalMux I__2143 (
            .O(N__9470),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__2142 (
            .O(N__9463),
            .I(\U409_TICK.TICK603_9 ));
    CascadeMux I__2141 (
            .O(N__9458),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    InMux I__2140 (
            .O(N__9455),
            .I(N__9452));
    LocalMux I__2139 (
            .O(N__9452),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__2138 (
            .O(N__9449),
            .I(N__9445));
    InMux I__2137 (
            .O(N__9448),
            .I(N__9442));
    LocalMux I__2136 (
            .O(N__9445),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__2135 (
            .O(N__9442),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    InMux I__2134 (
            .O(N__9437),
            .I(N__9434));
    LocalMux I__2133 (
            .O(N__9434),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__2132 (
            .O(N__9431),
            .I(N__9428));
    LocalMux I__2131 (
            .O(N__9428),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__2130 (
            .O(N__9425),
            .I(N__9421));
    InMux I__2129 (
            .O(N__9424),
            .I(N__9418));
    LocalMux I__2128 (
            .O(N__9421),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__2127 (
            .O(N__9418),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__2126 (
            .O(N__9413),
            .I(N__9409));
    InMux I__2125 (
            .O(N__9412),
            .I(N__9406));
    LocalMux I__2124 (
            .O(N__9409),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__2123 (
            .O(N__9406),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    InMux I__2122 (
            .O(N__9401),
            .I(N__9397));
    InMux I__2121 (
            .O(N__9400),
            .I(N__9394));
    LocalMux I__2120 (
            .O(N__9397),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__2119 (
            .O(N__9394),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    InMux I__2118 (
            .O(N__9389),
            .I(N__9386));
    LocalMux I__2117 (
            .O(N__9386),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    CascadeMux I__2116 (
            .O(N__9383),
            .I(N__9379));
    InMux I__2115 (
            .O(N__9382),
            .I(N__9373));
    InMux I__2114 (
            .O(N__9379),
            .I(N__9373));
    InMux I__2113 (
            .O(N__9378),
            .I(N__9370));
    LocalMux I__2112 (
            .O(N__9373),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__2111 (
            .O(N__9370),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    IoInMux I__2110 (
            .O(N__9365),
            .I(N__9362));
    LocalMux I__2109 (
            .O(N__9362),
            .I(N__9359));
    Span4Mux_s3_v I__2108 (
            .O(N__9359),
            .I(N__9356));
    Span4Mux_h I__2107 (
            .O(N__9356),
            .I(N__9353));
    Sp12to4 I__2106 (
            .O(N__9353),
            .I(N__9349));
    InMux I__2105 (
            .O(N__9352),
            .I(N__9346));
    Odrv12 I__2104 (
            .O(N__9349),
            .I(TICK60_c));
    LocalMux I__2103 (
            .O(N__9346),
            .I(TICK60_c));
    InMux I__2102 (
            .O(N__9341),
            .I(N__9338));
    LocalMux I__2101 (
            .O(N__9338),
            .I(N__9335));
    Span4Mux_h I__2100 (
            .O(N__9335),
            .I(N__9332));
    Span4Mux_v I__2099 (
            .O(N__9332),
            .I(N__9329));
    Span4Mux_v I__2098 (
            .O(N__9329),
            .I(N__9325));
    InMux I__2097 (
            .O(N__9328),
            .I(N__9322));
    Sp12to4 I__2096 (
            .O(N__9325),
            .I(N__9317));
    LocalMux I__2095 (
            .O(N__9322),
            .I(N__9317));
    Odrv12 I__2094 (
            .O(N__9317),
            .I(CIA_SPACE));
    CascadeMux I__2093 (
            .O(N__9314),
            .I(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ));
    CascadeMux I__2092 (
            .O(N__9311),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    InMux I__2091 (
            .O(N__9308),
            .I(N__9305));
    LocalMux I__2090 (
            .O(N__9305),
            .I(\U409_TICK.TICK503_8 ));
    CascadeMux I__2089 (
            .O(N__9302),
            .I(\U409_TICK.TICK503_11_cascade_ ));
    CascadeMux I__2088 (
            .O(N__9299),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    InMux I__2087 (
            .O(N__9296),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__2086 (
            .O(N__9293),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__2085 (
            .O(N__9290),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__2084 (
            .O(N__9287),
            .I(N__9283));
    InMux I__2083 (
            .O(N__9286),
            .I(N__9280));
    LocalMux I__2082 (
            .O(N__9283),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__2081 (
            .O(N__9280),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__2080 (
            .O(N__9275),
            .I(N__9271));
    InMux I__2079 (
            .O(N__9274),
            .I(N__9268));
    LocalMux I__2078 (
            .O(N__9271),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__2077 (
            .O(N__9268),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    CascadeMux I__2076 (
            .O(N__9263),
            .I(N__9260));
    InMux I__2075 (
            .O(N__9260),
            .I(N__9257));
    LocalMux I__2074 (
            .O(N__9257),
            .I(N__9253));
    InMux I__2073 (
            .O(N__9256),
            .I(N__9250));
    Odrv4 I__2072 (
            .O(N__9253),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__2071 (
            .O(N__9250),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__2070 (
            .O(N__9245),
            .I(N__9242));
    LocalMux I__2069 (
            .O(N__9242),
            .I(N__9237));
    InMux I__2068 (
            .O(N__9241),
            .I(N__9234));
    InMux I__2067 (
            .O(N__9240),
            .I(N__9231));
    Odrv12 I__2066 (
            .O(N__9237),
            .I(\U409_ADDRESS_DECODE.ATA_ENZ0 ));
    LocalMux I__2065 (
            .O(N__9234),
            .I(\U409_ADDRESS_DECODE.ATA_ENZ0 ));
    LocalMux I__2064 (
            .O(N__9231),
            .I(\U409_ADDRESS_DECODE.ATA_ENZ0 ));
    InMux I__2063 (
            .O(N__9224),
            .I(N__9221));
    LocalMux I__2062 (
            .O(N__9221),
            .I(N__9217));
    InMux I__2061 (
            .O(N__9220),
            .I(N__9214));
    Span4Mux_v I__2060 (
            .O(N__9217),
            .I(N__9210));
    LocalMux I__2059 (
            .O(N__9214),
            .I(N__9207));
    InMux I__2058 (
            .O(N__9213),
            .I(N__9204));
    Odrv4 I__2057 (
            .O(N__9210),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0 ));
    Odrv4 I__2056 (
            .O(N__9207),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0 ));
    LocalMux I__2055 (
            .O(N__9204),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0 ));
    IoInMux I__2054 (
            .O(N__9197),
            .I(N__9194));
    LocalMux I__2053 (
            .O(N__9194),
            .I(N__9191));
    IoSpan4Mux I__2052 (
            .O(N__9191),
            .I(N__9188));
    Sp12to4 I__2051 (
            .O(N__9188),
            .I(N__9185));
    Span12Mux_s7_h I__2050 (
            .O(N__9185),
            .I(N__9182));
    Odrv12 I__2049 (
            .O(N__9182),
            .I(U409_ADDRESS_DECODE_un1_ATA_ENn_i));
    CascadeMux I__2048 (
            .O(N__9179),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_ ));
    InMux I__2047 (
            .O(N__9176),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    InMux I__2046 (
            .O(N__9173),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__2045 (
            .O(N__9170),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__2044 (
            .O(N__9167),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__2043 (
            .O(N__9164),
            .I(bfn_13_7_0_));
    InMux I__2042 (
            .O(N__9161),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__2041 (
            .O(N__9158),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__2040 (
            .O(N__9155),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__2039 (
            .O(N__9152),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    CascadeMux I__2038 (
            .O(N__9149),
            .I(AGNUS_SPACE_0_cascade_));
    InMux I__2037 (
            .O(N__9146),
            .I(N__9143));
    LocalMux I__2036 (
            .O(N__9143),
            .I(N__9140));
    Span12Mux_v I__2035 (
            .O(N__9140),
            .I(N__9137));
    Span12Mux_h I__2034 (
            .O(N__9137),
            .I(N__9134));
    Odrv12 I__2033 (
            .O(N__9134),
            .I(TACKn_in));
    SRMux I__2032 (
            .O(N__9131),
            .I(N__9128));
    LocalMux I__2031 (
            .O(N__9128),
            .I(N__9122));
    SRMux I__2030 (
            .O(N__9127),
            .I(N__9119));
    SRMux I__2029 (
            .O(N__9126),
            .I(N__9116));
    SRMux I__2028 (
            .O(N__9125),
            .I(N__9113));
    Span4Mux_v I__2027 (
            .O(N__9122),
            .I(N__9108));
    LocalMux I__2026 (
            .O(N__9119),
            .I(N__9108));
    LocalMux I__2025 (
            .O(N__9116),
            .I(N__9105));
    LocalMux I__2024 (
            .O(N__9113),
            .I(N__9100));
    Span4Mux_v I__2023 (
            .O(N__9108),
            .I(N__9100));
    Span4Mux_v I__2022 (
            .O(N__9105),
            .I(N__9095));
    Span4Mux_v I__2021 (
            .O(N__9100),
            .I(N__9095));
    Odrv4 I__2020 (
            .O(N__9095),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__2019 (
            .O(N__9092),
            .I(N__9088));
    InMux I__2018 (
            .O(N__9091),
            .I(N__9085));
    LocalMux I__2017 (
            .O(N__9088),
            .I(N__9079));
    LocalMux I__2016 (
            .O(N__9085),
            .I(N__9079));
    InMux I__2015 (
            .O(N__9084),
            .I(N__9076));
    Span4Mux_h I__2014 (
            .O(N__9079),
            .I(N__9071));
    LocalMux I__2013 (
            .O(N__9076),
            .I(N__9071));
    Span4Mux_v I__2012 (
            .O(N__9071),
            .I(N__9066));
    InMux I__2011 (
            .O(N__9070),
            .I(N__9063));
    InMux I__2010 (
            .O(N__9069),
            .I(N__9060));
    Odrv4 I__2009 (
            .O(N__9066),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5 ));
    LocalMux I__2008 (
            .O(N__9063),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5 ));
    LocalMux I__2007 (
            .O(N__9060),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5 ));
    CascadeMux I__2006 (
            .O(N__9053),
            .I(N__9048));
    InMux I__2005 (
            .O(N__9052),
            .I(N__9045));
    InMux I__2004 (
            .O(N__9051),
            .I(N__9042));
    InMux I__2003 (
            .O(N__9048),
            .I(N__9039));
    LocalMux I__2002 (
            .O(N__9045),
            .I(N__9032));
    LocalMux I__2001 (
            .O(N__9042),
            .I(N__9032));
    LocalMux I__2000 (
            .O(N__9039),
            .I(N__9032));
    Span4Mux_h I__1999 (
            .O(N__9032),
            .I(N__9029));
    Span4Mux_v I__1998 (
            .O(N__9029),
            .I(N__9024));
    InMux I__1997 (
            .O(N__9028),
            .I(N__9021));
    InMux I__1996 (
            .O(N__9027),
            .I(N__9018));
    Odrv4 I__1995 (
            .O(N__9024),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4 ));
    LocalMux I__1994 (
            .O(N__9021),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4 ));
    LocalMux I__1993 (
            .O(N__9018),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4 ));
    IoInMux I__1992 (
            .O(N__9011),
            .I(N__9008));
    LocalMux I__1991 (
            .O(N__9008),
            .I(N__9005));
    IoSpan4Mux I__1990 (
            .O(N__9005),
            .I(N__9002));
    Span4Mux_s3_v I__1989 (
            .O(N__9002),
            .I(N__8999));
    Sp12to4 I__1988 (
            .O(N__8999),
            .I(N__8996));
    Span12Mux_h I__1987 (
            .O(N__8996),
            .I(N__8993));
    Odrv12 I__1986 (
            .O(N__8993),
            .I(BUFENn_c));
    InMux I__1985 (
            .O(N__8990),
            .I(N__8987));
    LocalMux I__1984 (
            .O(N__8987),
            .I(N__8984));
    Odrv12 I__1983 (
            .O(N__8984),
            .I(U409_ADDRESS_DECODE_PORTSIZE_0));
    CascadeMux I__1982 (
            .O(N__8981),
            .I(N__8977));
    InMux I__1981 (
            .O(N__8980),
            .I(N__8972));
    InMux I__1980 (
            .O(N__8977),
            .I(N__8972));
    LocalMux I__1979 (
            .O(N__8972),
            .I(AGNUS_SPACE_0));
    IoInMux I__1978 (
            .O(N__8969),
            .I(N__8966));
    LocalMux I__1977 (
            .O(N__8966),
            .I(N__8963));
    IoSpan4Mux I__1976 (
            .O(N__8963),
            .I(N__8960));
    Span4Mux_s0_v I__1975 (
            .O(N__8960),
            .I(N__8956));
    IoInMux I__1974 (
            .O(N__8959),
            .I(N__8953));
    Sp12to4 I__1973 (
            .O(N__8956),
            .I(N__8948));
    LocalMux I__1972 (
            .O(N__8953),
            .I(N__8948));
    Span12Mux_s11_v I__1971 (
            .O(N__8948),
            .I(N__8943));
    InMux I__1970 (
            .O(N__8947),
            .I(N__8940));
    CascadeMux I__1969 (
            .O(N__8946),
            .I(N__8937));
    Span12Mux_h I__1968 (
            .O(N__8943),
            .I(N__8934));
    LocalMux I__1967 (
            .O(N__8940),
            .I(N__8931));
    InMux I__1966 (
            .O(N__8937),
            .I(N__8928));
    Odrv12 I__1965 (
            .O(N__8934),
            .I(TACK_EN));
    Odrv4 I__1964 (
            .O(N__8931),
            .I(TACK_EN));
    LocalMux I__1963 (
            .O(N__8928),
            .I(TACK_EN));
    IoInMux I__1962 (
            .O(N__8921),
            .I(N__8918));
    LocalMux I__1961 (
            .O(N__8918),
            .I(N__8915));
    IoSpan4Mux I__1960 (
            .O(N__8915),
            .I(N__8912));
    Span4Mux_s2_v I__1959 (
            .O(N__8912),
            .I(N__8909));
    Sp12to4 I__1958 (
            .O(N__8909),
            .I(N__8906));
    Span12Mux_h I__1957 (
            .O(N__8906),
            .I(N__8903));
    Odrv12 I__1956 (
            .O(N__8903),
            .I(TCIn_1_i));
    IoInMux I__1955 (
            .O(N__8900),
            .I(N__8897));
    LocalMux I__1954 (
            .O(N__8897),
            .I(N__8894));
    Span12Mux_s2_v I__1953 (
            .O(N__8894),
            .I(N__8891));
    Odrv12 I__1952 (
            .O(N__8891),
            .I(RESETn_c_i));
    InMux I__1951 (
            .O(N__8888),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__1950 (
            .O(N__8885),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__1949 (
            .O(N__8882),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    IoInMux I__1948 (
            .O(N__8879),
            .I(N__8876));
    LocalMux I__1947 (
            .O(N__8876),
            .I(N__8873));
    Span12Mux_s7_v I__1946 (
            .O(N__8873),
            .I(N__8870));
    Odrv12 I__1945 (
            .O(N__8870),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn_i));
    InMux I__1944 (
            .O(N__8867),
            .I(N__8864));
    LocalMux I__1943 (
            .O(N__8864),
            .I(\U409_TRANSFER_ACK.N_28 ));
    InMux I__1942 (
            .O(N__8861),
            .I(N__8858));
    LocalMux I__1941 (
            .O(N__8858),
            .I(N__8855));
    Span4Mux_v I__1940 (
            .O(N__8855),
            .I(N__8851));
    InMux I__1939 (
            .O(N__8854),
            .I(N__8848));
    Odrv4 I__1938 (
            .O(N__8851),
            .I(\U409_TRANSFER_ACK.N_22 ));
    LocalMux I__1937 (
            .O(N__8848),
            .I(\U409_TRANSFER_ACK.N_22 ));
    CascadeMux I__1936 (
            .O(N__8843),
            .I(N__8839));
    InMux I__1935 (
            .O(N__8842),
            .I(N__8836));
    InMux I__1934 (
            .O(N__8839),
            .I(N__8832));
    LocalMux I__1933 (
            .O(N__8836),
            .I(N__8829));
    InMux I__1932 (
            .O(N__8835),
            .I(N__8826));
    LocalMux I__1931 (
            .O(N__8832),
            .I(N__8822));
    Span4Mux_h I__1930 (
            .O(N__8829),
            .I(N__8817));
    LocalMux I__1929 (
            .O(N__8826),
            .I(N__8817));
    InMux I__1928 (
            .O(N__8825),
            .I(N__8814));
    Span12Mux_v I__1927 (
            .O(N__8822),
            .I(N__8811));
    Span4Mux_h I__1926 (
            .O(N__8817),
            .I(N__8808));
    LocalMux I__1925 (
            .O(N__8814),
            .I(N__8805));
    Odrv12 I__1924 (
            .O(N__8811),
            .I(U409_ADDRESS_DECODE_ROMEN_1));
    Odrv4 I__1923 (
            .O(N__8808),
            .I(U409_ADDRESS_DECODE_ROMEN_1));
    Odrv4 I__1922 (
            .O(N__8805),
            .I(U409_ADDRESS_DECODE_ROMEN_1));
    InMux I__1921 (
            .O(N__8798),
            .I(N__8795));
    LocalMux I__1920 (
            .O(N__8795),
            .I(N__8791));
    CascadeMux I__1919 (
            .O(N__8794),
            .I(N__8788));
    Span4Mux_h I__1918 (
            .O(N__8791),
            .I(N__8785));
    InMux I__1917 (
            .O(N__8788),
            .I(N__8782));
    Odrv4 I__1916 (
            .O(N__8785),
            .I(\U409_TRANSFER_ACK.N_33_1 ));
    LocalMux I__1915 (
            .O(N__8782),
            .I(\U409_TRANSFER_ACK.N_33_1 ));
    CascadeMux I__1914 (
            .O(N__8777),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0_cascade_ ));
    InMux I__1913 (
            .O(N__8774),
            .I(N__8771));
    LocalMux I__1912 (
            .O(N__8771),
            .I(\U409_TRANSFER_ACK.N_33 ));
    InMux I__1911 (
            .O(N__8768),
            .I(N__8753));
    InMux I__1910 (
            .O(N__8767),
            .I(N__8753));
    InMux I__1909 (
            .O(N__8766),
            .I(N__8753));
    InMux I__1908 (
            .O(N__8765),
            .I(N__8753));
    InMux I__1907 (
            .O(N__8764),
            .I(N__8746));
    InMux I__1906 (
            .O(N__8763),
            .I(N__8746));
    InMux I__1905 (
            .O(N__8762),
            .I(N__8746));
    LocalMux I__1904 (
            .O(N__8753),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1903 (
            .O(N__8746),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    CascadeMux I__1902 (
            .O(N__8741),
            .I(N__8734));
    CascadeMux I__1901 (
            .O(N__8740),
            .I(N__8731));
    CascadeMux I__1900 (
            .O(N__8739),
            .I(N__8727));
    InMux I__1899 (
            .O(N__8738),
            .I(N__8715));
    InMux I__1898 (
            .O(N__8737),
            .I(N__8715));
    InMux I__1897 (
            .O(N__8734),
            .I(N__8715));
    InMux I__1896 (
            .O(N__8731),
            .I(N__8715));
    InMux I__1895 (
            .O(N__8730),
            .I(N__8715));
    InMux I__1894 (
            .O(N__8727),
            .I(N__8710));
    InMux I__1893 (
            .O(N__8726),
            .I(N__8710));
    LocalMux I__1892 (
            .O(N__8715),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1891 (
            .O(N__8710),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    InMux I__1890 (
            .O(N__8705),
            .I(N__8702));
    LocalMux I__1889 (
            .O(N__8702),
            .I(\U409_TRANSFER_ACK.N_34 ));
    InMux I__1888 (
            .O(N__8699),
            .I(N__8689));
    InMux I__1887 (
            .O(N__8698),
            .I(N__8689));
    InMux I__1886 (
            .O(N__8697),
            .I(N__8680));
    InMux I__1885 (
            .O(N__8696),
            .I(N__8680));
    InMux I__1884 (
            .O(N__8695),
            .I(N__8680));
    InMux I__1883 (
            .O(N__8694),
            .I(N__8680));
    LocalMux I__1882 (
            .O(N__8689),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1881 (
            .O(N__8680),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    CascadeMux I__1880 (
            .O(N__8675),
            .I(N__8667));
    CascadeMux I__1879 (
            .O(N__8674),
            .I(N__8664));
    InMux I__1878 (
            .O(N__8673),
            .I(N__8658));
    InMux I__1877 (
            .O(N__8672),
            .I(N__8658));
    InMux I__1876 (
            .O(N__8671),
            .I(N__8655));
    InMux I__1875 (
            .O(N__8670),
            .I(N__8646));
    InMux I__1874 (
            .O(N__8667),
            .I(N__8646));
    InMux I__1873 (
            .O(N__8664),
            .I(N__8646));
    InMux I__1872 (
            .O(N__8663),
            .I(N__8646));
    LocalMux I__1871 (
            .O(N__8658),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1870 (
            .O(N__8655),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1869 (
            .O(N__8646),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    InMux I__1868 (
            .O(N__8639),
            .I(N__8636));
    LocalMux I__1867 (
            .O(N__8636),
            .I(N__8633));
    Odrv4 I__1866 (
            .O(N__8633),
            .I(\U409_TRANSFER_ACK.N_45 ));
    InMux I__1865 (
            .O(N__8630),
            .I(N__8624));
    InMux I__1864 (
            .O(N__8629),
            .I(N__8621));
    InMux I__1863 (
            .O(N__8628),
            .I(N__8616));
    InMux I__1862 (
            .O(N__8627),
            .I(N__8616));
    LocalMux I__1861 (
            .O(N__8624),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__1860 (
            .O(N__8621),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__1859 (
            .O(N__8616),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    InMux I__1858 (
            .O(N__8609),
            .I(N__8605));
    InMux I__1857 (
            .O(N__8608),
            .I(N__8602));
    LocalMux I__1856 (
            .O(N__8605),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    LocalMux I__1855 (
            .O(N__8602),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    InMux I__1854 (
            .O(N__8597),
            .I(N__8591));
    InMux I__1853 (
            .O(N__8596),
            .I(N__8588));
    InMux I__1852 (
            .O(N__8595),
            .I(N__8583));
    InMux I__1851 (
            .O(N__8594),
            .I(N__8583));
    LocalMux I__1850 (
            .O(N__8591),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__1849 (
            .O(N__8588),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__1848 (
            .O(N__8583),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    SRMux I__1847 (
            .O(N__8576),
            .I(N__8546));
    SRMux I__1846 (
            .O(N__8575),
            .I(N__8546));
    SRMux I__1845 (
            .O(N__8574),
            .I(N__8546));
    SRMux I__1844 (
            .O(N__8573),
            .I(N__8546));
    SRMux I__1843 (
            .O(N__8572),
            .I(N__8546));
    SRMux I__1842 (
            .O(N__8571),
            .I(N__8546));
    SRMux I__1841 (
            .O(N__8570),
            .I(N__8546));
    SRMux I__1840 (
            .O(N__8569),
            .I(N__8546));
    SRMux I__1839 (
            .O(N__8568),
            .I(N__8546));
    SRMux I__1838 (
            .O(N__8567),
            .I(N__8546));
    GlobalMux I__1837 (
            .O(N__8546),
            .I(N__8543));
    gio2CtrlBuf I__1836 (
            .O(N__8543),
            .I(RESETn_c_i_g));
    InMux I__1835 (
            .O(N__8540),
            .I(N__8536));
    InMux I__1834 (
            .O(N__8539),
            .I(N__8533));
    LocalMux I__1833 (
            .O(N__8536),
            .I(N__8530));
    LocalMux I__1832 (
            .O(N__8533),
            .I(N__8527));
    Span4Mux_h I__1831 (
            .O(N__8530),
            .I(N__8522));
    Span4Mux_v I__1830 (
            .O(N__8527),
            .I(N__8522));
    Odrv4 I__1829 (
            .O(N__8522),
            .I(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0 ));
    InMux I__1828 (
            .O(N__8519),
            .I(N__8516));
    LocalMux I__1827 (
            .O(N__8516),
            .I(N__8513));
    Span4Mux_v I__1826 (
            .O(N__8513),
            .I(N__8509));
    InMux I__1825 (
            .O(N__8512),
            .I(N__8506));
    Odrv4 I__1824 (
            .O(N__8509),
            .I(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0 ));
    LocalMux I__1823 (
            .O(N__8506),
            .I(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0 ));
    InMux I__1822 (
            .O(N__8501),
            .I(N__8497));
    CascadeMux I__1821 (
            .O(N__8500),
            .I(N__8494));
    LocalMux I__1820 (
            .O(N__8497),
            .I(N__8488));
    InMux I__1819 (
            .O(N__8494),
            .I(N__8485));
    InMux I__1818 (
            .O(N__8493),
            .I(N__8480));
    InMux I__1817 (
            .O(N__8492),
            .I(N__8480));
    InMux I__1816 (
            .O(N__8491),
            .I(N__8476));
    Span4Mux_v I__1815 (
            .O(N__8488),
            .I(N__8467));
    LocalMux I__1814 (
            .O(N__8485),
            .I(N__8467));
    LocalMux I__1813 (
            .O(N__8480),
            .I(N__8464));
    InMux I__1812 (
            .O(N__8479),
            .I(N__8461));
    LocalMux I__1811 (
            .O(N__8476),
            .I(N__8458));
    InMux I__1810 (
            .O(N__8475),
            .I(N__8451));
    InMux I__1809 (
            .O(N__8474),
            .I(N__8451));
    InMux I__1808 (
            .O(N__8473),
            .I(N__8451));
    CascadeMux I__1807 (
            .O(N__8472),
            .I(N__8447));
    Span4Mux_v I__1806 (
            .O(N__8467),
            .I(N__8444));
    Span4Mux_v I__1805 (
            .O(N__8464),
            .I(N__8439));
    LocalMux I__1804 (
            .O(N__8461),
            .I(N__8439));
    Span4Mux_v I__1803 (
            .O(N__8458),
            .I(N__8434));
    LocalMux I__1802 (
            .O(N__8451),
            .I(N__8434));
    InMux I__1801 (
            .O(N__8450),
            .I(N__8431));
    InMux I__1800 (
            .O(N__8447),
            .I(N__8428));
    Span4Mux_h I__1799 (
            .O(N__8444),
            .I(N__8423));
    Span4Mux_v I__1798 (
            .O(N__8439),
            .I(N__8423));
    Span4Mux_v I__1797 (
            .O(N__8434),
            .I(N__8420));
    LocalMux I__1796 (
            .O(N__8431),
            .I(N__8417));
    LocalMux I__1795 (
            .O(N__8428),
            .I(N__8414));
    Span4Mux_h I__1794 (
            .O(N__8423),
            .I(N__8411));
    Span4Mux_h I__1793 (
            .O(N__8420),
            .I(N__8406));
    Span4Mux_v I__1792 (
            .O(N__8417),
            .I(N__8406));
    Span12Mux_v I__1791 (
            .O(N__8414),
            .I(N__8401));
    Sp12to4 I__1790 (
            .O(N__8411),
            .I(N__8401));
    Span4Mux_h I__1789 (
            .O(N__8406),
            .I(N__8398));
    Odrv12 I__1788 (
            .O(N__8401),
            .I(A_c_21));
    Odrv4 I__1787 (
            .O(N__8398),
            .I(A_c_21));
    InMux I__1786 (
            .O(N__8393),
            .I(N__8390));
    LocalMux I__1785 (
            .O(N__8390),
            .I(N__8386));
    InMux I__1784 (
            .O(N__8389),
            .I(N__8383));
    Span4Mux_v I__1783 (
            .O(N__8386),
            .I(N__8377));
    LocalMux I__1782 (
            .O(N__8383),
            .I(N__8377));
    InMux I__1781 (
            .O(N__8382),
            .I(N__8374));
    Sp12to4 I__1780 (
            .O(N__8377),
            .I(N__8369));
    LocalMux I__1779 (
            .O(N__8374),
            .I(N__8369));
    Span12Mux_v I__1778 (
            .O(N__8369),
            .I(N__8366));
    Span12Mux_h I__1777 (
            .O(N__8366),
            .I(N__8363));
    Odrv12 I__1776 (
            .O(N__8363),
            .I(OVL_c));
    CascadeMux I__1775 (
            .O(N__8360),
            .I(N__8356));
    CascadeMux I__1774 (
            .O(N__8359),
            .I(N__8353));
    InMux I__1773 (
            .O(N__8356),
            .I(N__8347));
    InMux I__1772 (
            .O(N__8353),
            .I(N__8342));
    InMux I__1771 (
            .O(N__8352),
            .I(N__8342));
    InMux I__1770 (
            .O(N__8351),
            .I(N__8337));
    InMux I__1769 (
            .O(N__8350),
            .I(N__8337));
    LocalMux I__1768 (
            .O(N__8347),
            .I(N__8334));
    LocalMux I__1767 (
            .O(N__8342),
            .I(N__8328));
    LocalMux I__1766 (
            .O(N__8337),
            .I(N__8328));
    Span4Mux_v I__1765 (
            .O(N__8334),
            .I(N__8324));
    InMux I__1764 (
            .O(N__8333),
            .I(N__8321));
    Span4Mux_h I__1763 (
            .O(N__8328),
            .I(N__8318));
    InMux I__1762 (
            .O(N__8327),
            .I(N__8315));
    Odrv4 I__1761 (
            .O(N__8324),
            .I(CONFIGURED));
    LocalMux I__1760 (
            .O(N__8321),
            .I(CONFIGURED));
    Odrv4 I__1759 (
            .O(N__8318),
            .I(CONFIGURED));
    LocalMux I__1758 (
            .O(N__8315),
            .I(CONFIGURED));
    InMux I__1757 (
            .O(N__8306),
            .I(N__8303));
    LocalMux I__1756 (
            .O(N__8303),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1 ));
    InMux I__1755 (
            .O(N__8300),
            .I(N__8297));
    LocalMux I__1754 (
            .O(N__8297),
            .I(N__8294));
    Span4Mux_v I__1753 (
            .O(N__8294),
            .I(N__8291));
    Odrv4 I__1752 (
            .O(N__8291),
            .I(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_1 ));
    InMux I__1751 (
            .O(N__8288),
            .I(N__8285));
    LocalMux I__1750 (
            .O(N__8285),
            .I(N__8282));
    Odrv4 I__1749 (
            .O(N__8282),
            .I(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_2 ));
    CascadeMux I__1748 (
            .O(N__8279),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_ ));
    IoInMux I__1747 (
            .O(N__8276),
            .I(N__8273));
    LocalMux I__1746 (
            .O(N__8273),
            .I(N__8270));
    Span12Mux_s5_h I__1745 (
            .O(N__8270),
            .I(N__8267));
    Span12Mux_h I__1744 (
            .O(N__8267),
            .I(N__8264));
    Odrv12 I__1743 (
            .O(N__8264),
            .I(U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i));
    InMux I__1742 (
            .O(N__8261),
            .I(N__8254));
    InMux I__1741 (
            .O(N__8260),
            .I(N__8249));
    InMux I__1740 (
            .O(N__8259),
            .I(N__8246));
    InMux I__1739 (
            .O(N__8258),
            .I(N__8243));
    InMux I__1738 (
            .O(N__8257),
            .I(N__8240));
    LocalMux I__1737 (
            .O(N__8254),
            .I(N__8237));
    InMux I__1736 (
            .O(N__8253),
            .I(N__8234));
    InMux I__1735 (
            .O(N__8252),
            .I(N__8231));
    LocalMux I__1734 (
            .O(N__8249),
            .I(N__8226));
    LocalMux I__1733 (
            .O(N__8246),
            .I(N__8226));
    LocalMux I__1732 (
            .O(N__8243),
            .I(N__8221));
    LocalMux I__1731 (
            .O(N__8240),
            .I(N__8221));
    Span4Mux_v I__1730 (
            .O(N__8237),
            .I(N__8214));
    LocalMux I__1729 (
            .O(N__8234),
            .I(N__8214));
    LocalMux I__1728 (
            .O(N__8231),
            .I(N__8214));
    Span4Mux_v I__1727 (
            .O(N__8226),
            .I(N__8211));
    Span4Mux_v I__1726 (
            .O(N__8221),
            .I(N__8206));
    Span4Mux_v I__1725 (
            .O(N__8214),
            .I(N__8206));
    Sp12to4 I__1724 (
            .O(N__8211),
            .I(N__8201));
    Sp12to4 I__1723 (
            .O(N__8206),
            .I(N__8201));
    Span12Mux_h I__1722 (
            .O(N__8201),
            .I(N__8198));
    Span12Mux_v I__1721 (
            .O(N__8198),
            .I(N__8195));
    Odrv12 I__1720 (
            .O(N__8195),
            .I(RnW_c));
    InMux I__1719 (
            .O(N__8192),
            .I(N__8187));
    CascadeMux I__1718 (
            .O(N__8191),
            .I(N__8184));
    InMux I__1717 (
            .O(N__8190),
            .I(N__8181));
    LocalMux I__1716 (
            .O(N__8187),
            .I(N__8178));
    InMux I__1715 (
            .O(N__8184),
            .I(N__8175));
    LocalMux I__1714 (
            .O(N__8181),
            .I(N__8172));
    Span4Mux_h I__1713 (
            .O(N__8178),
            .I(N__8169));
    LocalMux I__1712 (
            .O(N__8175),
            .I(N__8164));
    Span4Mux_v I__1711 (
            .O(N__8172),
            .I(N__8164));
    Span4Mux_v I__1710 (
            .O(N__8169),
            .I(N__8161));
    Sp12to4 I__1709 (
            .O(N__8164),
            .I(N__8158));
    Sp12to4 I__1708 (
            .O(N__8161),
            .I(N__8153));
    Span12Mux_h I__1707 (
            .O(N__8158),
            .I(N__8153));
    Span12Mux_v I__1706 (
            .O(N__8153),
            .I(N__8150));
    Odrv12 I__1705 (
            .O(N__8150),
            .I(D_in_5));
    CascadeMux I__1704 (
            .O(N__8147),
            .I(un1_AUTOCONFIG_SPACE_cascade_));
    InMux I__1703 (
            .O(N__8144),
            .I(N__8140));
    InMux I__1702 (
            .O(N__8143),
            .I(N__8137));
    LocalMux I__1701 (
            .O(N__8140),
            .I(ATA_BASE_1));
    LocalMux I__1700 (
            .O(N__8137),
            .I(ATA_BASE_1));
    InMux I__1699 (
            .O(N__8132),
            .I(N__8125));
    InMux I__1698 (
            .O(N__8131),
            .I(N__8125));
    InMux I__1697 (
            .O(N__8130),
            .I(N__8122));
    LocalMux I__1696 (
            .O(N__8125),
            .I(\U409_AUTOCONFIG.STATE_RNIS3FU2Z0Z_0 ));
    LocalMux I__1695 (
            .O(N__8122),
            .I(\U409_AUTOCONFIG.STATE_RNIS3FU2Z0Z_0 ));
    InMux I__1694 (
            .O(N__8117),
            .I(N__8108));
    InMux I__1693 (
            .O(N__8116),
            .I(N__8108));
    CascadeMux I__1692 (
            .O(N__8115),
            .I(N__8104));
    CascadeMux I__1691 (
            .O(N__8114),
            .I(N__8101));
    CascadeMux I__1690 (
            .O(N__8113),
            .I(N__8098));
    LocalMux I__1689 (
            .O(N__8108),
            .I(N__8092));
    InMux I__1688 (
            .O(N__8107),
            .I(N__8081));
    InMux I__1687 (
            .O(N__8104),
            .I(N__8081));
    InMux I__1686 (
            .O(N__8101),
            .I(N__8081));
    InMux I__1685 (
            .O(N__8098),
            .I(N__8081));
    InMux I__1684 (
            .O(N__8097),
            .I(N__8081));
    InMux I__1683 (
            .O(N__8096),
            .I(N__8076));
    InMux I__1682 (
            .O(N__8095),
            .I(N__8076));
    Span4Mux_h I__1681 (
            .O(N__8092),
            .I(N__8071));
    LocalMux I__1680 (
            .O(N__8081),
            .I(N__8071));
    LocalMux I__1679 (
            .O(N__8076),
            .I(N__8067));
    Span4Mux_h I__1678 (
            .O(N__8071),
            .I(N__8064));
    InMux I__1677 (
            .O(N__8070),
            .I(N__8061));
    Odrv4 I__1676 (
            .O(N__8067),
            .I(un1_AUTOCONFIG_SPACE));
    Odrv4 I__1675 (
            .O(N__8064),
            .I(un1_AUTOCONFIG_SPACE));
    LocalMux I__1674 (
            .O(N__8061),
            .I(un1_AUTOCONFIG_SPACE));
    CascadeMux I__1673 (
            .O(N__8054),
            .I(N__8050));
    InMux I__1672 (
            .O(N__8053),
            .I(N__8047));
    InMux I__1671 (
            .O(N__8050),
            .I(N__8044));
    LocalMux I__1670 (
            .O(N__8047),
            .I(N__8039));
    LocalMux I__1669 (
            .O(N__8044),
            .I(N__8039));
    Span4Mux_v I__1668 (
            .O(N__8039),
            .I(N__8035));
    CascadeMux I__1667 (
            .O(N__8038),
            .I(N__8032));
    Span4Mux_h I__1666 (
            .O(N__8035),
            .I(N__8029));
    InMux I__1665 (
            .O(N__8032),
            .I(N__8026));
    Sp12to4 I__1664 (
            .O(N__8029),
            .I(N__8021));
    LocalMux I__1663 (
            .O(N__8026),
            .I(N__8021));
    Span12Mux_v I__1662 (
            .O(N__8021),
            .I(N__8018));
    Odrv12 I__1661 (
            .O(N__8018),
            .I(D_in_7));
    InMux I__1660 (
            .O(N__8015),
            .I(N__8011));
    InMux I__1659 (
            .O(N__8014),
            .I(N__8008));
    LocalMux I__1658 (
            .O(N__8011),
            .I(ATA_BASE_3));
    LocalMux I__1657 (
            .O(N__8008),
            .I(ATA_BASE_3));
    CascadeMux I__1656 (
            .O(N__8003),
            .I(N__7994));
    CascadeMux I__1655 (
            .O(N__8002),
            .I(N__7991));
    InMux I__1654 (
            .O(N__8001),
            .I(N__7988));
    InMux I__1653 (
            .O(N__8000),
            .I(N__7985));
    InMux I__1652 (
            .O(N__7999),
            .I(N__7982));
    InMux I__1651 (
            .O(N__7998),
            .I(N__7979));
    InMux I__1650 (
            .O(N__7997),
            .I(N__7976));
    InMux I__1649 (
            .O(N__7994),
            .I(N__7971));
    InMux I__1648 (
            .O(N__7991),
            .I(N__7971));
    LocalMux I__1647 (
            .O(N__7988),
            .I(N__7968));
    LocalMux I__1646 (
            .O(N__7985),
            .I(N__7965));
    LocalMux I__1645 (
            .O(N__7982),
            .I(N__7960));
    LocalMux I__1644 (
            .O(N__7979),
            .I(N__7957));
    LocalMux I__1643 (
            .O(N__7976),
            .I(N__7952));
    LocalMux I__1642 (
            .O(N__7971),
            .I(N__7944));
    Glb2LocalMux I__1641 (
            .O(N__7968),
            .I(N__7910));
    Glb2LocalMux I__1640 (
            .O(N__7965),
            .I(N__7910));
    ClkMux I__1639 (
            .O(N__7964),
            .I(N__7910));
    ClkMux I__1638 (
            .O(N__7963),
            .I(N__7910));
    Glb2LocalMux I__1637 (
            .O(N__7960),
            .I(N__7910));
    Glb2LocalMux I__1636 (
            .O(N__7957),
            .I(N__7910));
    ClkMux I__1635 (
            .O(N__7956),
            .I(N__7910));
    ClkMux I__1634 (
            .O(N__7955),
            .I(N__7910));
    Glb2LocalMux I__1633 (
            .O(N__7952),
            .I(N__7910));
    ClkMux I__1632 (
            .O(N__7951),
            .I(N__7910));
    ClkMux I__1631 (
            .O(N__7950),
            .I(N__7910));
    ClkMux I__1630 (
            .O(N__7949),
            .I(N__7910));
    ClkMux I__1629 (
            .O(N__7948),
            .I(N__7910));
    ClkMux I__1628 (
            .O(N__7947),
            .I(N__7910));
    Glb2LocalMux I__1627 (
            .O(N__7944),
            .I(N__7910));
    ClkMux I__1626 (
            .O(N__7943),
            .I(N__7910));
    GlobalMux I__1625 (
            .O(N__7910),
            .I(N__7907));
    gio2CtrlBuf I__1624 (
            .O(N__7907),
            .I(CLK40_IN_c_g));
    IoInMux I__1623 (
            .O(N__7904),
            .I(N__7901));
    LocalMux I__1622 (
            .O(N__7901),
            .I(N__7898));
    Span12Mux_s6_v I__1621 (
            .O(N__7898),
            .I(N__7895));
    Odrv12 I__1620 (
            .O(N__7895),
            .I(GB_BUFFER_CLK40_IN_c_g_THRU_CO));
    InMux I__1619 (
            .O(N__7892),
            .I(N__7886));
    InMux I__1618 (
            .O(N__7891),
            .I(N__7879));
    InMux I__1617 (
            .O(N__7890),
            .I(N__7879));
    InMux I__1616 (
            .O(N__7889),
            .I(N__7879));
    LocalMux I__1615 (
            .O(N__7886),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__1614 (
            .O(N__7879),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    InMux I__1613 (
            .O(N__7874),
            .I(N__7869));
    InMux I__1612 (
            .O(N__7873),
            .I(N__7864));
    InMux I__1611 (
            .O(N__7872),
            .I(N__7864));
    LocalMux I__1610 (
            .O(N__7869),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    LocalMux I__1609 (
            .O(N__7864),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    IoInMux I__1608 (
            .O(N__7859),
            .I(N__7856));
    LocalMux I__1607 (
            .O(N__7856),
            .I(N__7853));
    Span4Mux_s3_v I__1606 (
            .O(N__7853),
            .I(N__7850));
    Span4Mux_v I__1605 (
            .O(N__7850),
            .I(N__7847));
    Span4Mux_v I__1604 (
            .O(N__7847),
            .I(N__7844));
    Span4Mux_h I__1603 (
            .O(N__7844),
            .I(N__7840));
    InMux I__1602 (
            .O(N__7843),
            .I(N__7837));
    Odrv4 I__1601 (
            .O(N__7840),
            .I(TICK50_c));
    LocalMux I__1600 (
            .O(N__7837),
            .I(TICK50_c));
    InMux I__1599 (
            .O(N__7832),
            .I(N__7829));
    LocalMux I__1598 (
            .O(N__7829),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0 ));
    CascadeMux I__1597 (
            .O(N__7826),
            .I(N__7823));
    InMux I__1596 (
            .O(N__7823),
            .I(N__7819));
    InMux I__1595 (
            .O(N__7822),
            .I(N__7816));
    LocalMux I__1594 (
            .O(N__7819),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__1593 (
            .O(N__7816),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__1592 (
            .O(N__7811),
            .I(N__7807));
    InMux I__1591 (
            .O(N__7810),
            .I(N__7804));
    LocalMux I__1590 (
            .O(N__7807),
            .I(N__7801));
    LocalMux I__1589 (
            .O(N__7804),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    Odrv12 I__1588 (
            .O(N__7801),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    CascadeMux I__1587 (
            .O(N__7796),
            .I(N__7793));
    InMux I__1586 (
            .O(N__7793),
            .I(N__7789));
    CascadeMux I__1585 (
            .O(N__7792),
            .I(N__7786));
    LocalMux I__1584 (
            .O(N__7789),
            .I(N__7783));
    InMux I__1583 (
            .O(N__7786),
            .I(N__7780));
    Odrv4 I__1582 (
            .O(N__7783),
            .I(AC_TACK));
    LocalMux I__1581 (
            .O(N__7780),
            .I(AC_TACK));
    InMux I__1580 (
            .O(N__7775),
            .I(N__7772));
    LocalMux I__1579 (
            .O(N__7772),
            .I(N__7769));
    Span4Mux_h I__1578 (
            .O(N__7769),
            .I(N__7766));
    Odrv4 I__1577 (
            .O(N__7766),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER5_1 ));
    CascadeMux I__1576 (
            .O(N__7763),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ));
    CascadeMux I__1575 (
            .O(N__7760),
            .I(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ));
    IoInMux I__1574 (
            .O(N__7757),
            .I(N__7753));
    IoInMux I__1573 (
            .O(N__7756),
            .I(N__7750));
    LocalMux I__1572 (
            .O(N__7753),
            .I(N__7744));
    LocalMux I__1571 (
            .O(N__7750),
            .I(N__7744));
    IoInMux I__1570 (
            .O(N__7749),
            .I(N__7741));
    IoSpan4Mux I__1569 (
            .O(N__7744),
            .I(N__7738));
    LocalMux I__1568 (
            .O(N__7741),
            .I(N__7735));
    Span4Mux_s2_v I__1567 (
            .O(N__7738),
            .I(N__7730));
    Span4Mux_s2_v I__1566 (
            .O(N__7735),
            .I(N__7730));
    Span4Mux_v I__1565 (
            .O(N__7730),
            .I(N__7727));
    Sp12to4 I__1564 (
            .O(N__7727),
            .I(N__7724));
    Span12Mux_h I__1563 (
            .O(N__7724),
            .I(N__7719));
    InMux I__1562 (
            .O(N__7723),
            .I(N__7714));
    InMux I__1561 (
            .O(N__7722),
            .I(N__7714));
    Odrv12 I__1560 (
            .O(N__7719),
            .I(TACK_OUTn));
    LocalMux I__1559 (
            .O(N__7714),
            .I(TACK_OUTn));
    CascadeMux I__1558 (
            .O(N__7709),
            .I(N__7703));
    CascadeMux I__1557 (
            .O(N__7708),
            .I(N__7699));
    InMux I__1556 (
            .O(N__7707),
            .I(N__7695));
    InMux I__1555 (
            .O(N__7706),
            .I(N__7692));
    InMux I__1554 (
            .O(N__7703),
            .I(N__7683));
    InMux I__1553 (
            .O(N__7702),
            .I(N__7683));
    InMux I__1552 (
            .O(N__7699),
            .I(N__7683));
    InMux I__1551 (
            .O(N__7698),
            .I(N__7683));
    LocalMux I__1550 (
            .O(N__7695),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1549 (
            .O(N__7692),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1548 (
            .O(N__7683),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    InMux I__1547 (
            .O(N__7676),
            .I(N__7670));
    InMux I__1546 (
            .O(N__7675),
            .I(N__7667));
    InMux I__1545 (
            .O(N__7674),
            .I(N__7662));
    InMux I__1544 (
            .O(N__7673),
            .I(N__7662));
    LocalMux I__1543 (
            .O(N__7670),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1542 (
            .O(N__7667),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1541 (
            .O(N__7662),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    InMux I__1540 (
            .O(N__7655),
            .I(N__7651));
    InMux I__1539 (
            .O(N__7654),
            .I(N__7648));
    LocalMux I__1538 (
            .O(N__7651),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_1_out ));
    LocalMux I__1537 (
            .O(N__7648),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_1_out ));
    InMux I__1536 (
            .O(N__7643),
            .I(N__7640));
    LocalMux I__1535 (
            .O(N__7640),
            .I(N__7636));
    CascadeMux I__1534 (
            .O(N__7639),
            .I(N__7633));
    Span4Mux_h I__1533 (
            .O(N__7636),
            .I(N__7629));
    InMux I__1532 (
            .O(N__7633),
            .I(N__7624));
    InMux I__1531 (
            .O(N__7632),
            .I(N__7624));
    Span4Mux_h I__1530 (
            .O(N__7629),
            .I(N__7619));
    LocalMux I__1529 (
            .O(N__7624),
            .I(N__7619));
    Span4Mux_h I__1528 (
            .O(N__7619),
            .I(N__7616));
    Span4Mux_v I__1527 (
            .O(N__7616),
            .I(N__7613));
    Span4Mux_v I__1526 (
            .O(N__7613),
            .I(N__7610));
    Span4Mux_v I__1525 (
            .O(N__7610),
            .I(N__7607));
    Odrv4 I__1524 (
            .O(N__7607),
            .I(TM_c_0));
    InMux I__1523 (
            .O(N__7604),
            .I(N__7601));
    LocalMux I__1522 (
            .O(N__7601),
            .I(N__7596));
    InMux I__1521 (
            .O(N__7600),
            .I(N__7591));
    InMux I__1520 (
            .O(N__7599),
            .I(N__7591));
    Span4Mux_v I__1519 (
            .O(N__7596),
            .I(N__7588));
    LocalMux I__1518 (
            .O(N__7591),
            .I(N__7585));
    Span4Mux_h I__1517 (
            .O(N__7588),
            .I(N__7580));
    Span4Mux_v I__1516 (
            .O(N__7585),
            .I(N__7580));
    Span4Mux_h I__1515 (
            .O(N__7580),
            .I(N__7577));
    Sp12to4 I__1514 (
            .O(N__7577),
            .I(N__7574));
    Odrv12 I__1513 (
            .O(N__7574),
            .I(TM_c_1));
    InMux I__1512 (
            .O(N__7571),
            .I(N__7566));
    InMux I__1511 (
            .O(N__7570),
            .I(N__7561));
    InMux I__1510 (
            .O(N__7569),
            .I(N__7561));
    LocalMux I__1509 (
            .O(N__7566),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__1508 (
            .O(N__7561),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__1507 (
            .O(N__7556),
            .I(N__7550));
    InMux I__1506 (
            .O(N__7555),
            .I(N__7550));
    LocalMux I__1505 (
            .O(N__7550),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    CascadeMux I__1504 (
            .O(N__7547),
            .I(N__7541));
    InMux I__1503 (
            .O(N__7546),
            .I(N__7537));
    InMux I__1502 (
            .O(N__7545),
            .I(N__7528));
    InMux I__1501 (
            .O(N__7544),
            .I(N__7528));
    InMux I__1500 (
            .O(N__7541),
            .I(N__7528));
    InMux I__1499 (
            .O(N__7540),
            .I(N__7528));
    LocalMux I__1498 (
            .O(N__7537),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__1497 (
            .O(N__7528),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    InMux I__1496 (
            .O(N__7523),
            .I(N__7520));
    LocalMux I__1495 (
            .O(N__7520),
            .I(\U409_TRANSFER_ACK.N_17_mux ));
    CascadeMux I__1494 (
            .O(N__7517),
            .I(N__7512));
    InMux I__1493 (
            .O(N__7516),
            .I(N__7507));
    InMux I__1492 (
            .O(N__7515),
            .I(N__7507));
    InMux I__1491 (
            .O(N__7512),
            .I(N__7504));
    LocalMux I__1490 (
            .O(N__7507),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1489 (
            .O(N__7504),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    InMux I__1488 (
            .O(N__7499),
            .I(N__7496));
    LocalMux I__1487 (
            .O(N__7496),
            .I(N__7493));
    Odrv12 I__1486 (
            .O(N__7493),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1Z0Z_0 ));
    CascadeMux I__1485 (
            .O(N__7490),
            .I(N__7487));
    InMux I__1484 (
            .O(N__7487),
            .I(N__7481));
    InMux I__1483 (
            .O(N__7486),
            .I(N__7481));
    LocalMux I__1482 (
            .O(N__7481),
            .I(N__7477));
    CascadeMux I__1481 (
            .O(N__7480),
            .I(N__7473));
    Span4Mux_v I__1480 (
            .O(N__7477),
            .I(N__7470));
    InMux I__1479 (
            .O(N__7476),
            .I(N__7467));
    InMux I__1478 (
            .O(N__7473),
            .I(N__7464));
    Span4Mux_h I__1477 (
            .O(N__7470),
            .I(N__7455));
    LocalMux I__1476 (
            .O(N__7467),
            .I(N__7455));
    LocalMux I__1475 (
            .O(N__7464),
            .I(N__7455));
    InMux I__1474 (
            .O(N__7463),
            .I(N__7451));
    CascadeMux I__1473 (
            .O(N__7462),
            .I(N__7448));
    Span4Mux_v I__1472 (
            .O(N__7455),
            .I(N__7445));
    InMux I__1471 (
            .O(N__7454),
            .I(N__7442));
    LocalMux I__1470 (
            .O(N__7451),
            .I(N__7438));
    InMux I__1469 (
            .O(N__7448),
            .I(N__7435));
    Span4Mux_v I__1468 (
            .O(N__7445),
            .I(N__7430));
    LocalMux I__1467 (
            .O(N__7442),
            .I(N__7430));
    InMux I__1466 (
            .O(N__7441),
            .I(N__7427));
    Span4Mux_v I__1465 (
            .O(N__7438),
            .I(N__7422));
    LocalMux I__1464 (
            .O(N__7435),
            .I(N__7422));
    Span4Mux_h I__1463 (
            .O(N__7430),
            .I(N__7417));
    LocalMux I__1462 (
            .O(N__7427),
            .I(N__7417));
    Span4Mux_v I__1461 (
            .O(N__7422),
            .I(N__7414));
    Span4Mux_v I__1460 (
            .O(N__7417),
            .I(N__7411));
    Sp12to4 I__1459 (
            .O(N__7414),
            .I(N__7408));
    Span4Mux_v I__1458 (
            .O(N__7411),
            .I(N__7405));
    Span12Mux_v I__1457 (
            .O(N__7408),
            .I(N__7402));
    Span4Mux_v I__1456 (
            .O(N__7405),
            .I(N__7399));
    Span12Mux_h I__1455 (
            .O(N__7402),
            .I(N__7396));
    Span4Mux_h I__1454 (
            .O(N__7399),
            .I(N__7393));
    Odrv12 I__1453 (
            .O(N__7396),
            .I(A_c_22));
    Odrv4 I__1452 (
            .O(N__7393),
            .I(A_c_22));
    InMux I__1451 (
            .O(N__7388),
            .I(N__7381));
    InMux I__1450 (
            .O(N__7387),
            .I(N__7381));
    InMux I__1449 (
            .O(N__7386),
            .I(N__7377));
    LocalMux I__1448 (
            .O(N__7381),
            .I(N__7374));
    InMux I__1447 (
            .O(N__7380),
            .I(N__7371));
    LocalMux I__1446 (
            .O(N__7377),
            .I(N__7367));
    Span4Mux_v I__1445 (
            .O(N__7374),
            .I(N__7362));
    LocalMux I__1444 (
            .O(N__7371),
            .I(N__7362));
    InMux I__1443 (
            .O(N__7370),
            .I(N__7359));
    Span4Mux_v I__1442 (
            .O(N__7367),
            .I(N__7355));
    Span4Mux_v I__1441 (
            .O(N__7362),
            .I(N__7351));
    LocalMux I__1440 (
            .O(N__7359),
            .I(N__7348));
    InMux I__1439 (
            .O(N__7358),
            .I(N__7345));
    Span4Mux_v I__1438 (
            .O(N__7355),
            .I(N__7342));
    InMux I__1437 (
            .O(N__7354),
            .I(N__7339));
    Span4Mux_h I__1436 (
            .O(N__7351),
            .I(N__7334));
    Span4Mux_v I__1435 (
            .O(N__7348),
            .I(N__7334));
    LocalMux I__1434 (
            .O(N__7345),
            .I(N__7331));
    Sp12to4 I__1433 (
            .O(N__7342),
            .I(N__7326));
    LocalMux I__1432 (
            .O(N__7339),
            .I(N__7326));
    Span4Mux_h I__1431 (
            .O(N__7334),
            .I(N__7321));
    Span4Mux_v I__1430 (
            .O(N__7331),
            .I(N__7321));
    Span12Mux_h I__1429 (
            .O(N__7326),
            .I(N__7316));
    Sp12to4 I__1428 (
            .O(N__7321),
            .I(N__7316));
    Odrv12 I__1427 (
            .O(N__7316),
            .I(A_c_23));
    InMux I__1426 (
            .O(N__7313),
            .I(N__7310));
    LocalMux I__1425 (
            .O(N__7310),
            .I(N__7307));
    Odrv4 I__1424 (
            .O(N__7307),
            .I(\U409_TRANSFER_ACK.N_43 ));
    IoInMux I__1423 (
            .O(N__7304),
            .I(N__7301));
    LocalMux I__1422 (
            .O(N__7301),
            .I(N__7298));
    Span4Mux_s3_v I__1421 (
            .O(N__7298),
            .I(N__7295));
    Span4Mux_h I__1420 (
            .O(N__7295),
            .I(N__7292));
    Span4Mux_v I__1419 (
            .O(N__7292),
            .I(N__7289));
    Span4Mux_v I__1418 (
            .O(N__7289),
            .I(N__7286));
    Span4Mux_v I__1417 (
            .O(N__7286),
            .I(N__7282));
    InMux I__1416 (
            .O(N__7285),
            .I(N__7279));
    Odrv4 I__1415 (
            .O(N__7282),
            .I(ROMENn_c));
    LocalMux I__1414 (
            .O(N__7279),
            .I(ROMENn_c));
    InMux I__1413 (
            .O(N__7274),
            .I(N__7271));
    LocalMux I__1412 (
            .O(N__7271),
            .I(N__7267));
    InMux I__1411 (
            .O(N__7270),
            .I(N__7264));
    Span4Mux_h I__1410 (
            .O(N__7267),
            .I(N__7259));
    LocalMux I__1409 (
            .O(N__7264),
            .I(N__7259));
    Odrv4 I__1408 (
            .O(N__7259),
            .I(\U409_TRANSFER_ACK.un1_AUTOVECTOR_0 ));
    InMux I__1407 (
            .O(N__7256),
            .I(N__7253));
    LocalMux I__1406 (
            .O(N__7253),
            .I(N__7249));
    InMux I__1405 (
            .O(N__7252),
            .I(N__7246));
    Span4Mux_v I__1404 (
            .O(N__7249),
            .I(N__7240));
    LocalMux I__1403 (
            .O(N__7246),
            .I(N__7240));
    InMux I__1402 (
            .O(N__7245),
            .I(N__7237));
    Span4Mux_h I__1401 (
            .O(N__7240),
            .I(N__7229));
    LocalMux I__1400 (
            .O(N__7237),
            .I(N__7229));
    InMux I__1399 (
            .O(N__7236),
            .I(N__7226));
    InMux I__1398 (
            .O(N__7235),
            .I(N__7223));
    InMux I__1397 (
            .O(N__7234),
            .I(N__7220));
    Span4Mux_v I__1396 (
            .O(N__7229),
            .I(N__7217));
    LocalMux I__1395 (
            .O(N__7226),
            .I(N__7214));
    LocalMux I__1394 (
            .O(N__7223),
            .I(N__7211));
    LocalMux I__1393 (
            .O(N__7220),
            .I(N__7208));
    Span4Mux_v I__1392 (
            .O(N__7217),
            .I(N__7203));
    Span4Mux_v I__1391 (
            .O(N__7214),
            .I(N__7203));
    Span4Mux_v I__1390 (
            .O(N__7211),
            .I(N__7200));
    Span12Mux_h I__1389 (
            .O(N__7208),
            .I(N__7197));
    Sp12to4 I__1388 (
            .O(N__7203),
            .I(N__7192));
    Sp12to4 I__1387 (
            .O(N__7200),
            .I(N__7192));
    Span12Mux_v I__1386 (
            .O(N__7197),
            .I(N__7189));
    Span12Mux_h I__1385 (
            .O(N__7192),
            .I(N__7186));
    Odrv12 I__1384 (
            .O(N__7189),
            .I(TSn_c));
    Odrv12 I__1383 (
            .O(N__7186),
            .I(TSn_c));
    InMux I__1382 (
            .O(N__7181),
            .I(N__7178));
    LocalMux I__1381 (
            .O(N__7178),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1 ));
    InMux I__1380 (
            .O(N__7175),
            .I(N__7169));
    InMux I__1379 (
            .O(N__7174),
            .I(N__7169));
    LocalMux I__1378 (
            .O(N__7169),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    InMux I__1377 (
            .O(N__7166),
            .I(N__7162));
    InMux I__1376 (
            .O(N__7165),
            .I(N__7159));
    LocalMux I__1375 (
            .O(N__7162),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    LocalMux I__1374 (
            .O(N__7159),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    CascadeMux I__1373 (
            .O(N__7154),
            .I(\U409_TRANSFER_ACK.N_17_mux_cascade_ ));
    CascadeMux I__1372 (
            .O(N__7151),
            .I(\U409_TRANSFER_ACK.N_3_0_cascade_ ));
    CascadeMux I__1371 (
            .O(N__7148),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0_cascade_ ));
    InMux I__1370 (
            .O(N__7145),
            .I(N__7142));
    LocalMux I__1369 (
            .O(N__7142),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0 ));
    InMux I__1368 (
            .O(N__7139),
            .I(N__7136));
    LocalMux I__1367 (
            .O(N__7136),
            .I(\U409_TRANSFER_ACK.N_3_0 ));
    CascadeMux I__1366 (
            .O(N__7133),
            .I(\U409_TRANSFER_ACK.N_6_0_cascade_ ));
    InMux I__1365 (
            .O(N__7130),
            .I(N__7126));
    InMux I__1364 (
            .O(N__7129),
            .I(N__7123));
    LocalMux I__1363 (
            .O(N__7126),
            .I(ATA_BASE_2));
    LocalMux I__1362 (
            .O(N__7123),
            .I(ATA_BASE_2));
    CascadeMux I__1361 (
            .O(N__7118),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2_cascade_ ));
    InMux I__1360 (
            .O(N__7115),
            .I(N__7111));
    InMux I__1359 (
            .O(N__7114),
            .I(N__7108));
    LocalMux I__1358 (
            .O(N__7111),
            .I(N__7105));
    LocalMux I__1357 (
            .O(N__7108),
            .I(ATA_BASE_7));
    Odrv4 I__1356 (
            .O(N__7105),
            .I(ATA_BASE_7));
    InMux I__1355 (
            .O(N__7100),
            .I(N__7097));
    LocalMux I__1354 (
            .O(N__7097),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ));
    InMux I__1353 (
            .O(N__7094),
            .I(N__7091));
    LocalMux I__1352 (
            .O(N__7091),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_0 ));
    CascadeMux I__1351 (
            .O(N__7088),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_5_cascade_ ));
    CascadeMux I__1350 (
            .O(N__7085),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_ ));
    InMux I__1349 (
            .O(N__7082),
            .I(N__7078));
    InMux I__1348 (
            .O(N__7081),
            .I(N__7075));
    LocalMux I__1347 (
            .O(N__7078),
            .I(\U409_AUTOCONFIG.un1_STATE_6_0 ));
    LocalMux I__1346 (
            .O(N__7075),
            .I(\U409_AUTOCONFIG.un1_STATE_6_0 ));
    InMux I__1345 (
            .O(N__7070),
            .I(N__7057));
    InMux I__1344 (
            .O(N__7069),
            .I(N__7054));
    InMux I__1343 (
            .O(N__7068),
            .I(N__7051));
    InMux I__1342 (
            .O(N__7067),
            .I(N__7046));
    InMux I__1341 (
            .O(N__7066),
            .I(N__7046));
    InMux I__1340 (
            .O(N__7065),
            .I(N__7039));
    InMux I__1339 (
            .O(N__7064),
            .I(N__7039));
    InMux I__1338 (
            .O(N__7063),
            .I(N__7039));
    InMux I__1337 (
            .O(N__7062),
            .I(N__7036));
    CascadeMux I__1336 (
            .O(N__7061),
            .I(N__7033));
    InMux I__1335 (
            .O(N__7060),
            .I(N__7028));
    LocalMux I__1334 (
            .O(N__7057),
            .I(N__7025));
    LocalMux I__1333 (
            .O(N__7054),
            .I(N__7017));
    LocalMux I__1332 (
            .O(N__7051),
            .I(N__7017));
    LocalMux I__1331 (
            .O(N__7046),
            .I(N__7017));
    LocalMux I__1330 (
            .O(N__7039),
            .I(N__7011));
    LocalMux I__1329 (
            .O(N__7036),
            .I(N__7011));
    InMux I__1328 (
            .O(N__7033),
            .I(N__7004));
    InMux I__1327 (
            .O(N__7032),
            .I(N__7004));
    InMux I__1326 (
            .O(N__7031),
            .I(N__7004));
    LocalMux I__1325 (
            .O(N__7028),
            .I(N__7001));
    Span4Mux_v I__1324 (
            .O(N__7025),
            .I(N__6998));
    InMux I__1323 (
            .O(N__7024),
            .I(N__6995));
    Span4Mux_v I__1322 (
            .O(N__7017),
            .I(N__6992));
    InMux I__1321 (
            .O(N__7016),
            .I(N__6989));
    Span4Mux_h I__1320 (
            .O(N__7011),
            .I(N__6984));
    LocalMux I__1319 (
            .O(N__7004),
            .I(N__6984));
    Sp12to4 I__1318 (
            .O(N__7001),
            .I(N__6981));
    Sp12to4 I__1317 (
            .O(N__6998),
            .I(N__6972));
    LocalMux I__1316 (
            .O(N__6995),
            .I(N__6972));
    Sp12to4 I__1315 (
            .O(N__6992),
            .I(N__6972));
    LocalMux I__1314 (
            .O(N__6989),
            .I(N__6972));
    Span4Mux_v I__1313 (
            .O(N__6984),
            .I(N__6969));
    Span12Mux_v I__1312 (
            .O(N__6981),
            .I(N__6966));
    Span12Mux_h I__1311 (
            .O(N__6972),
            .I(N__6963));
    Span4Mux_h I__1310 (
            .O(N__6969),
            .I(N__6960));
    Span12Mux_h I__1309 (
            .O(N__6966),
            .I(N__6955));
    Span12Mux_v I__1308 (
            .O(N__6963),
            .I(N__6955));
    Sp12to4 I__1307 (
            .O(N__6960),
            .I(N__6952));
    Odrv12 I__1306 (
            .O(N__6955),
            .I(A_c_1));
    Odrv12 I__1305 (
            .O(N__6952),
            .I(A_c_1));
    InMux I__1304 (
            .O(N__6947),
            .I(N__6944));
    LocalMux I__1303 (
            .O(N__6944),
            .I(N__6940));
    InMux I__1302 (
            .O(N__6943),
            .I(N__6937));
    Span4Mux_v I__1301 (
            .O(N__6940),
            .I(N__6933));
    LocalMux I__1300 (
            .O(N__6937),
            .I(N__6930));
    InMux I__1299 (
            .O(N__6936),
            .I(N__6927));
    Span4Mux_h I__1298 (
            .O(N__6933),
            .I(N__6919));
    Span4Mux_v I__1297 (
            .O(N__6930),
            .I(N__6919));
    LocalMux I__1296 (
            .O(N__6927),
            .I(N__6919));
    InMux I__1295 (
            .O(N__6926),
            .I(N__6916));
    Span4Mux_v I__1294 (
            .O(N__6919),
            .I(N__6912));
    LocalMux I__1293 (
            .O(N__6916),
            .I(N__6909));
    InMux I__1292 (
            .O(N__6915),
            .I(N__6906));
    Span4Mux_v I__1291 (
            .O(N__6912),
            .I(N__6903));
    Span4Mux_v I__1290 (
            .O(N__6909),
            .I(N__6898));
    LocalMux I__1289 (
            .O(N__6906),
            .I(N__6898));
    Span4Mux_v I__1288 (
            .O(N__6903),
            .I(N__6895));
    Sp12to4 I__1287 (
            .O(N__6898),
            .I(N__6892));
    Sp12to4 I__1286 (
            .O(N__6895),
            .I(N__6887));
    Span12Mux_v I__1285 (
            .O(N__6892),
            .I(N__6887));
    Odrv12 I__1284 (
            .O(N__6887),
            .I(A_c_17));
    InMux I__1283 (
            .O(N__6884),
            .I(N__6881));
    LocalMux I__1282 (
            .O(N__6881),
            .I(\U409_ADDRESS_DECODE.un2_ATA_SPACEZ0Z_0 ));
    InMux I__1281 (
            .O(N__6878),
            .I(N__6875));
    LocalMux I__1280 (
            .O(N__6875),
            .I(N__6871));
    InMux I__1279 (
            .O(N__6874),
            .I(N__6868));
    Odrv12 I__1278 (
            .O(N__6871),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn));
    LocalMux I__1277 (
            .O(N__6868),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn));
    CascadeMux I__1276 (
            .O(N__6863),
            .I(U409_ADDRESS_DECODE_PORTSIZE_0_cascade_));
    IoInMux I__1275 (
            .O(N__6860),
            .I(N__6857));
    LocalMux I__1274 (
            .O(N__6857),
            .I(N__6854));
    Span4Mux_s3_v I__1273 (
            .O(N__6854),
            .I(N__6851));
    Span4Mux_h I__1272 (
            .O(N__6851),
            .I(N__6848));
    Sp12to4 I__1271 (
            .O(N__6848),
            .I(N__6845));
    Span12Mux_v I__1270 (
            .O(N__6845),
            .I(N__6842));
    Odrv12 I__1269 (
            .O(N__6842),
            .I(PORTSIZE_0_i));
    CascadeMux I__1268 (
            .O(N__6839),
            .I(N__6835));
    InMux I__1267 (
            .O(N__6838),
            .I(N__6832));
    InMux I__1266 (
            .O(N__6835),
            .I(N__6829));
    LocalMux I__1265 (
            .O(N__6832),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    LocalMux I__1264 (
            .O(N__6829),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    CascadeMux I__1263 (
            .O(N__6824),
            .I(N__6819));
    CascadeMux I__1262 (
            .O(N__6823),
            .I(N__6815));
    CascadeMux I__1261 (
            .O(N__6822),
            .I(N__6812));
    InMux I__1260 (
            .O(N__6819),
            .I(N__6806));
    InMux I__1259 (
            .O(N__6818),
            .I(N__6806));
    InMux I__1258 (
            .O(N__6815),
            .I(N__6799));
    InMux I__1257 (
            .O(N__6812),
            .I(N__6799));
    InMux I__1256 (
            .O(N__6811),
            .I(N__6799));
    LocalMux I__1255 (
            .O(N__6806),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__1254 (
            .O(N__6799),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    CascadeMux I__1253 (
            .O(N__6794),
            .I(N__6791));
    InMux I__1252 (
            .O(N__6791),
            .I(N__6785));
    InMux I__1251 (
            .O(N__6790),
            .I(N__6780));
    InMux I__1250 (
            .O(N__6789),
            .I(N__6780));
    InMux I__1249 (
            .O(N__6788),
            .I(N__6777));
    LocalMux I__1248 (
            .O(N__6785),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1247 (
            .O(N__6780),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1246 (
            .O(N__6777),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__1245 (
            .O(N__6770),
            .I(N__6762));
    InMux I__1244 (
            .O(N__6769),
            .I(N__6755));
    InMux I__1243 (
            .O(N__6768),
            .I(N__6755));
    InMux I__1242 (
            .O(N__6767),
            .I(N__6755));
    InMux I__1241 (
            .O(N__6766),
            .I(N__6752));
    InMux I__1240 (
            .O(N__6765),
            .I(N__6747));
    InMux I__1239 (
            .O(N__6762),
            .I(N__6747));
    LocalMux I__1238 (
            .O(N__6755),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1237 (
            .O(N__6752),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1236 (
            .O(N__6747),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    InMux I__1235 (
            .O(N__6740),
            .I(N__6735));
    InMux I__1234 (
            .O(N__6739),
            .I(N__6730));
    InMux I__1233 (
            .O(N__6738),
            .I(N__6730));
    LocalMux I__1232 (
            .O(N__6735),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__1231 (
            .O(N__6730),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    InMux I__1230 (
            .O(N__6725),
            .I(N__6722));
    LocalMux I__1229 (
            .O(N__6722),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_2 ));
    InMux I__1228 (
            .O(N__6719),
            .I(N__6715));
    InMux I__1227 (
            .O(N__6718),
            .I(N__6710));
    LocalMux I__1226 (
            .O(N__6715),
            .I(N__6707));
    InMux I__1225 (
            .O(N__6714),
            .I(N__6702));
    InMux I__1224 (
            .O(N__6713),
            .I(N__6702));
    LocalMux I__1223 (
            .O(N__6710),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    Odrv4 I__1222 (
            .O(N__6707),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1221 (
            .O(N__6702),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    InMux I__1220 (
            .O(N__6695),
            .I(N__6692));
    LocalMux I__1219 (
            .O(N__6692),
            .I(N__6689));
    Odrv4 I__1218 (
            .O(N__6689),
            .I(\U409_AUTOCONFIG.STATE_d_2 ));
    InMux I__1217 (
            .O(N__6686),
            .I(N__6683));
    LocalMux I__1216 (
            .O(N__6683),
            .I(N__6678));
    InMux I__1215 (
            .O(N__6682),
            .I(N__6675));
    InMux I__1214 (
            .O(N__6681),
            .I(N__6672));
    Span4Mux_v I__1213 (
            .O(N__6678),
            .I(N__6669));
    LocalMux I__1212 (
            .O(N__6675),
            .I(N__6664));
    LocalMux I__1211 (
            .O(N__6672),
            .I(N__6664));
    Sp12to4 I__1210 (
            .O(N__6669),
            .I(N__6661));
    Span4Mux_v I__1209 (
            .O(N__6664),
            .I(N__6658));
    Odrv12 I__1208 (
            .O(N__6661),
            .I(\U409_AUTOCONFIG.un1_AZ0Z_16 ));
    Odrv4 I__1207 (
            .O(N__6658),
            .I(\U409_AUTOCONFIG.un1_AZ0Z_16 ));
    InMux I__1206 (
            .O(N__6653),
            .I(N__6647));
    InMux I__1205 (
            .O(N__6652),
            .I(N__6643));
    InMux I__1204 (
            .O(N__6651),
            .I(N__6638));
    InMux I__1203 (
            .O(N__6650),
            .I(N__6638));
    LocalMux I__1202 (
            .O(N__6647),
            .I(N__6635));
    InMux I__1201 (
            .O(N__6646),
            .I(N__6632));
    LocalMux I__1200 (
            .O(N__6643),
            .I(N__6625));
    LocalMux I__1199 (
            .O(N__6638),
            .I(N__6625));
    Span4Mux_v I__1198 (
            .O(N__6635),
            .I(N__6620));
    LocalMux I__1197 (
            .O(N__6632),
            .I(N__6620));
    InMux I__1196 (
            .O(N__6631),
            .I(N__6617));
    InMux I__1195 (
            .O(N__6630),
            .I(N__6613));
    Span4Mux_v I__1194 (
            .O(N__6625),
            .I(N__6606));
    Span4Mux_v I__1193 (
            .O(N__6620),
            .I(N__6606));
    LocalMux I__1192 (
            .O(N__6617),
            .I(N__6606));
    InMux I__1191 (
            .O(N__6616),
            .I(N__6603));
    LocalMux I__1190 (
            .O(N__6613),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    Odrv4 I__1189 (
            .O(N__6606),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__1188 (
            .O(N__6603),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    CascadeMux I__1187 (
            .O(N__6596),
            .I(N__6593));
    InMux I__1186 (
            .O(N__6593),
            .I(N__6589));
    InMux I__1185 (
            .O(N__6592),
            .I(N__6586));
    LocalMux I__1184 (
            .O(N__6589),
            .I(N__6581));
    LocalMux I__1183 (
            .O(N__6586),
            .I(N__6581));
    Span4Mux_v I__1182 (
            .O(N__6581),
            .I(N__6578));
    Sp12to4 I__1181 (
            .O(N__6578),
            .I(N__6575));
    Span12Mux_h I__1180 (
            .O(N__6575),
            .I(N__6572));
    Span12Mux_v I__1179 (
            .O(N__6572),
            .I(N__6569));
    Odrv12 I__1178 (
            .O(N__6569),
            .I(D_in_4));
    InMux I__1177 (
            .O(N__6566),
            .I(N__6563));
    LocalMux I__1176 (
            .O(N__6563),
            .I(N__6560));
    Span4Mux_v I__1175 (
            .O(N__6560),
            .I(N__6556));
    InMux I__1174 (
            .O(N__6559),
            .I(N__6553));
    Odrv4 I__1173 (
            .O(N__6556),
            .I(BRIDGE_BASE_0));
    LocalMux I__1172 (
            .O(N__6553),
            .I(BRIDGE_BASE_0));
    InMux I__1171 (
            .O(N__6548),
            .I(N__6536));
    InMux I__1170 (
            .O(N__6547),
            .I(N__6536));
    InMux I__1169 (
            .O(N__6546),
            .I(N__6536));
    InMux I__1168 (
            .O(N__6545),
            .I(N__6533));
    InMux I__1167 (
            .O(N__6544),
            .I(N__6530));
    InMux I__1166 (
            .O(N__6543),
            .I(N__6527));
    LocalMux I__1165 (
            .O(N__6536),
            .I(N__6524));
    LocalMux I__1164 (
            .O(N__6533),
            .I(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ));
    LocalMux I__1163 (
            .O(N__6530),
            .I(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ));
    LocalMux I__1162 (
            .O(N__6527),
            .I(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ));
    Odrv12 I__1161 (
            .O(N__6524),
            .I(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ));
    InMux I__1160 (
            .O(N__6515),
            .I(N__6512));
    LocalMux I__1159 (
            .O(N__6512),
            .I(N__6509));
    Span4Mux_v I__1158 (
            .O(N__6509),
            .I(N__6505));
    InMux I__1157 (
            .O(N__6508),
            .I(N__6502));
    Odrv4 I__1156 (
            .O(N__6505),
            .I(BRIDGE_BASE_1));
    LocalMux I__1155 (
            .O(N__6502),
            .I(BRIDGE_BASE_1));
    InMux I__1154 (
            .O(N__6497),
            .I(N__6493));
    InMux I__1153 (
            .O(N__6496),
            .I(N__6488));
    LocalMux I__1152 (
            .O(N__6493),
            .I(N__6485));
    InMux I__1151 (
            .O(N__6492),
            .I(N__6482));
    InMux I__1150 (
            .O(N__6491),
            .I(N__6479));
    LocalMux I__1149 (
            .O(N__6488),
            .I(N__6472));
    Span4Mux_h I__1148 (
            .O(N__6485),
            .I(N__6467));
    LocalMux I__1147 (
            .O(N__6482),
            .I(N__6467));
    LocalMux I__1146 (
            .O(N__6479),
            .I(N__6464));
    InMux I__1145 (
            .O(N__6478),
            .I(N__6459));
    InMux I__1144 (
            .O(N__6477),
            .I(N__6459));
    InMux I__1143 (
            .O(N__6476),
            .I(N__6456));
    InMux I__1142 (
            .O(N__6475),
            .I(N__6453));
    Span4Mux_h I__1141 (
            .O(N__6472),
            .I(N__6448));
    Span4Mux_v I__1140 (
            .O(N__6467),
            .I(N__6448));
    Span4Mux_v I__1139 (
            .O(N__6464),
            .I(N__6445));
    LocalMux I__1138 (
            .O(N__6459),
            .I(N__6442));
    LocalMux I__1137 (
            .O(N__6456),
            .I(N__6437));
    LocalMux I__1136 (
            .O(N__6453),
            .I(N__6437));
    Span4Mux_h I__1135 (
            .O(N__6448),
            .I(N__6434));
    Span4Mux_v I__1134 (
            .O(N__6445),
            .I(N__6431));
    Span4Mux_v I__1133 (
            .O(N__6442),
            .I(N__6428));
    Span4Mux_v I__1132 (
            .O(N__6437),
            .I(N__6425));
    Span4Mux_v I__1131 (
            .O(N__6434),
            .I(N__6422));
    Sp12to4 I__1130 (
            .O(N__6431),
            .I(N__6415));
    Sp12to4 I__1129 (
            .O(N__6428),
            .I(N__6415));
    Sp12to4 I__1128 (
            .O(N__6425),
            .I(N__6415));
    Sp12to4 I__1127 (
            .O(N__6422),
            .I(N__6410));
    Span12Mux_h I__1126 (
            .O(N__6415),
            .I(N__6410));
    Span12Mux_v I__1125 (
            .O(N__6410),
            .I(N__6407));
    Odrv12 I__1124 (
            .O(N__6407),
            .I(A_c_19));
    CascadeMux I__1123 (
            .O(N__6404),
            .I(N__6399));
    InMux I__1122 (
            .O(N__6403),
            .I(N__6395));
    CascadeMux I__1121 (
            .O(N__6402),
            .I(N__6392));
    InMux I__1120 (
            .O(N__6399),
            .I(N__6388));
    InMux I__1119 (
            .O(N__6398),
            .I(N__6385));
    LocalMux I__1118 (
            .O(N__6395),
            .I(N__6382));
    InMux I__1117 (
            .O(N__6392),
            .I(N__6379));
    InMux I__1116 (
            .O(N__6391),
            .I(N__6376));
    LocalMux I__1115 (
            .O(N__6388),
            .I(N__6373));
    LocalMux I__1114 (
            .O(N__6385),
            .I(N__6370));
    Span4Mux_v I__1113 (
            .O(N__6382),
            .I(N__6363));
    LocalMux I__1112 (
            .O(N__6379),
            .I(N__6363));
    LocalMux I__1111 (
            .O(N__6376),
            .I(N__6363));
    Span4Mux_v I__1110 (
            .O(N__6373),
            .I(N__6359));
    Span4Mux_v I__1109 (
            .O(N__6370),
            .I(N__6354));
    Span4Mux_v I__1108 (
            .O(N__6363),
            .I(N__6354));
    InMux I__1107 (
            .O(N__6362),
            .I(N__6351));
    Sp12to4 I__1106 (
            .O(N__6359),
            .I(N__6344));
    Sp12to4 I__1105 (
            .O(N__6354),
            .I(N__6344));
    LocalMux I__1104 (
            .O(N__6351),
            .I(N__6344));
    Span12Mux_h I__1103 (
            .O(N__6344),
            .I(N__6341));
    Span12Mux_v I__1102 (
            .O(N__6341),
            .I(N__6338));
    Odrv12 I__1101 (
            .O(N__6338),
            .I(A_c_18));
    InMux I__1100 (
            .O(N__6335),
            .I(N__6332));
    LocalMux I__1099 (
            .O(N__6332),
            .I(N__6329));
    Odrv12 I__1098 (
            .O(N__6329),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    InMux I__1097 (
            .O(N__6326),
            .I(N__6323));
    LocalMux I__1096 (
            .O(N__6323),
            .I(N__6320));
    Odrv4 I__1095 (
            .O(N__6320),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_11_0 ));
    InMux I__1094 (
            .O(N__6317),
            .I(N__6310));
    InMux I__1093 (
            .O(N__6316),
            .I(N__6303));
    InMux I__1092 (
            .O(N__6315),
            .I(N__6303));
    InMux I__1091 (
            .O(N__6314),
            .I(N__6303));
    InMux I__1090 (
            .O(N__6313),
            .I(N__6300));
    LocalMux I__1089 (
            .O(N__6310),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__1088 (
            .O(N__6303),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__1087 (
            .O(N__6300),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    InMux I__1086 (
            .O(N__6293),
            .I(N__6287));
    InMux I__1085 (
            .O(N__6292),
            .I(N__6282));
    InMux I__1084 (
            .O(N__6291),
            .I(N__6282));
    InMux I__1083 (
            .O(N__6290),
            .I(N__6279));
    LocalMux I__1082 (
            .O(N__6287),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__1081 (
            .O(N__6282),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__1080 (
            .O(N__6279),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    CascadeMux I__1079 (
            .O(N__6272),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_5_cascade_ ));
    InMux I__1078 (
            .O(N__6269),
            .I(N__6266));
    LocalMux I__1077 (
            .O(N__6266),
            .I(N__6263));
    Span4Mux_v I__1076 (
            .O(N__6263),
            .I(N__6259));
    InMux I__1075 (
            .O(N__6262),
            .I(N__6256));
    Odrv4 I__1074 (
            .O(N__6259),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    LocalMux I__1073 (
            .O(N__6256),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    CascadeMux I__1072 (
            .O(N__6251),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_cascade_ ));
    CascadeMux I__1071 (
            .O(N__6248),
            .I(N__6245));
    InMux I__1070 (
            .O(N__6245),
            .I(N__6242));
    LocalMux I__1069 (
            .O(N__6242),
            .I(N__6238));
    InMux I__1068 (
            .O(N__6241),
            .I(N__6235));
    Odrv12 I__1067 (
            .O(N__6238),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    LocalMux I__1066 (
            .O(N__6235),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    InMux I__1065 (
            .O(N__6230),
            .I(N__6227));
    LocalMux I__1064 (
            .O(N__6227),
            .I(N__6218));
    InMux I__1063 (
            .O(N__6226),
            .I(N__6213));
    InMux I__1062 (
            .O(N__6225),
            .I(N__6213));
    InMux I__1061 (
            .O(N__6224),
            .I(N__6208));
    InMux I__1060 (
            .O(N__6223),
            .I(N__6208));
    InMux I__1059 (
            .O(N__6222),
            .I(N__6205));
    InMux I__1058 (
            .O(N__6221),
            .I(N__6202));
    Span4Mux_v I__1057 (
            .O(N__6218),
            .I(N__6199));
    LocalMux I__1056 (
            .O(N__6213),
            .I(N__6196));
    LocalMux I__1055 (
            .O(N__6208),
            .I(N__6189));
    LocalMux I__1054 (
            .O(N__6205),
            .I(N__6189));
    LocalMux I__1053 (
            .O(N__6202),
            .I(N__6189));
    Span4Mux_h I__1052 (
            .O(N__6199),
            .I(N__6184));
    Span4Mux_v I__1051 (
            .O(N__6196),
            .I(N__6184));
    Span12Mux_v I__1050 (
            .O(N__6189),
            .I(N__6179));
    Sp12to4 I__1049 (
            .O(N__6184),
            .I(N__6179));
    Odrv12 I__1048 (
            .O(N__6179),
            .I(A_c_7));
    InMux I__1047 (
            .O(N__6176),
            .I(N__6173));
    LocalMux I__1046 (
            .O(N__6173),
            .I(N__6170));
    Odrv4 I__1045 (
            .O(N__6170),
            .I(\U409_AUTOCONFIG.ATA_BASE11Z0Z_1 ));
    CascadeMux I__1044 (
            .O(N__6167),
            .I(N__6162));
    InMux I__1043 (
            .O(N__6166),
            .I(N__6153));
    InMux I__1042 (
            .O(N__6165),
            .I(N__6153));
    InMux I__1041 (
            .O(N__6162),
            .I(N__6150));
    InMux I__1040 (
            .O(N__6161),
            .I(N__6145));
    InMux I__1039 (
            .O(N__6160),
            .I(N__6140));
    InMux I__1038 (
            .O(N__6159),
            .I(N__6140));
    InMux I__1037 (
            .O(N__6158),
            .I(N__6137));
    LocalMux I__1036 (
            .O(N__6153),
            .I(N__6134));
    LocalMux I__1035 (
            .O(N__6150),
            .I(N__6131));
    InMux I__1034 (
            .O(N__6149),
            .I(N__6128));
    CascadeMux I__1033 (
            .O(N__6148),
            .I(N__6125));
    LocalMux I__1032 (
            .O(N__6145),
            .I(N__6121));
    LocalMux I__1031 (
            .O(N__6140),
            .I(N__6115));
    LocalMux I__1030 (
            .O(N__6137),
            .I(N__6115));
    Span4Mux_v I__1029 (
            .O(N__6134),
            .I(N__6112));
    Span4Mux_h I__1028 (
            .O(N__6131),
            .I(N__6107));
    LocalMux I__1027 (
            .O(N__6128),
            .I(N__6107));
    InMux I__1026 (
            .O(N__6125),
            .I(N__6102));
    InMux I__1025 (
            .O(N__6124),
            .I(N__6102));
    Span4Mux_v I__1024 (
            .O(N__6121),
            .I(N__6099));
    InMux I__1023 (
            .O(N__6120),
            .I(N__6096));
    Span12Mux_v I__1022 (
            .O(N__6115),
            .I(N__6083));
    Sp12to4 I__1021 (
            .O(N__6112),
            .I(N__6083));
    Sp12to4 I__1020 (
            .O(N__6107),
            .I(N__6083));
    LocalMux I__1019 (
            .O(N__6102),
            .I(N__6083));
    Sp12to4 I__1018 (
            .O(N__6099),
            .I(N__6083));
    LocalMux I__1017 (
            .O(N__6096),
            .I(N__6083));
    Odrv12 I__1016 (
            .O(N__6083),
            .I(A_c_5));
    InMux I__1015 (
            .O(N__6080),
            .I(N__6071));
    InMux I__1014 (
            .O(N__6079),
            .I(N__6068));
    InMux I__1013 (
            .O(N__6078),
            .I(N__6063));
    InMux I__1012 (
            .O(N__6077),
            .I(N__6063));
    InMux I__1011 (
            .O(N__6076),
            .I(N__6060));
    InMux I__1010 (
            .O(N__6075),
            .I(N__6057));
    InMux I__1009 (
            .O(N__6074),
            .I(N__6054));
    LocalMux I__1008 (
            .O(N__6071),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    LocalMux I__1007 (
            .O(N__6068),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    LocalMux I__1006 (
            .O(N__6063),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    LocalMux I__1005 (
            .O(N__6060),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    LocalMux I__1004 (
            .O(N__6057),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    LocalMux I__1003 (
            .O(N__6054),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    CascadeMux I__1002 (
            .O(N__6041),
            .I(\U409_AUTOCONFIG.ATA_BASE11_cascade_ ));
    InMux I__1001 (
            .O(N__6038),
            .I(N__6034));
    CascadeMux I__1000 (
            .O(N__6037),
            .I(N__6028));
    LocalMux I__999 (
            .O(N__6034),
            .I(N__6023));
    InMux I__998 (
            .O(N__6033),
            .I(N__6020));
    InMux I__997 (
            .O(N__6032),
            .I(N__6017));
    InMux I__996 (
            .O(N__6031),
            .I(N__6012));
    InMux I__995 (
            .O(N__6028),
            .I(N__6012));
    InMux I__994 (
            .O(N__6027),
            .I(N__6009));
    InMux I__993 (
            .O(N__6026),
            .I(N__6006));
    Span4Mux_v I__992 (
            .O(N__6023),
            .I(N__6001));
    LocalMux I__991 (
            .O(N__6020),
            .I(N__6001));
    LocalMux I__990 (
            .O(N__6017),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__989 (
            .O(N__6012),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__988 (
            .O(N__6009),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__987 (
            .O(N__6006),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    Odrv4 I__986 (
            .O(N__6001),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    InMux I__985 (
            .O(N__5990),
            .I(N__5986));
    CascadeMux I__984 (
            .O(N__5989),
            .I(N__5983));
    LocalMux I__983 (
            .O(N__5986),
            .I(N__5976));
    InMux I__982 (
            .O(N__5983),
            .I(N__5973));
    InMux I__981 (
            .O(N__5982),
            .I(N__5963));
    InMux I__980 (
            .O(N__5981),
            .I(N__5963));
    InMux I__979 (
            .O(N__5980),
            .I(N__5963));
    InMux I__978 (
            .O(N__5979),
            .I(N__5963));
    Span4Mux_v I__977 (
            .O(N__5976),
            .I(N__5960));
    LocalMux I__976 (
            .O(N__5973),
            .I(N__5957));
    InMux I__975 (
            .O(N__5972),
            .I(N__5954));
    LocalMux I__974 (
            .O(N__5963),
            .I(N__5951));
    Odrv4 I__973 (
            .O(N__5960),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ));
    Odrv4 I__972 (
            .O(N__5957),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ));
    LocalMux I__971 (
            .O(N__5954),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ));
    Odrv4 I__970 (
            .O(N__5951),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ));
    InMux I__969 (
            .O(N__5942),
            .I(N__5936));
    InMux I__968 (
            .O(N__5941),
            .I(N__5933));
    InMux I__967 (
            .O(N__5940),
            .I(N__5930));
    CascadeMux I__966 (
            .O(N__5939),
            .I(N__5927));
    LocalMux I__965 (
            .O(N__5936),
            .I(N__5921));
    LocalMux I__964 (
            .O(N__5933),
            .I(N__5916));
    LocalMux I__963 (
            .O(N__5930),
            .I(N__5916));
    InMux I__962 (
            .O(N__5927),
            .I(N__5909));
    InMux I__961 (
            .O(N__5926),
            .I(N__5909));
    InMux I__960 (
            .O(N__5925),
            .I(N__5909));
    InMux I__959 (
            .O(N__5924),
            .I(N__5906));
    Span4Mux_v I__958 (
            .O(N__5921),
            .I(N__5903));
    Span4Mux_v I__957 (
            .O(N__5916),
            .I(N__5900));
    LocalMux I__956 (
            .O(N__5909),
            .I(N__5895));
    LocalMux I__955 (
            .O(N__5906),
            .I(N__5895));
    Odrv4 I__954 (
            .O(N__5903),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_6 ));
    Odrv4 I__953 (
            .O(N__5900),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_6 ));
    Odrv4 I__952 (
            .O(N__5895),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_6 ));
    InMux I__951 (
            .O(N__5888),
            .I(N__5882));
    InMux I__950 (
            .O(N__5887),
            .I(N__5882));
    LocalMux I__949 (
            .O(N__5882),
            .I(ATA_BASE_6));
    CascadeMux I__948 (
            .O(N__5879),
            .I(N__5874));
    InMux I__947 (
            .O(N__5878),
            .I(N__5869));
    InMux I__946 (
            .O(N__5877),
            .I(N__5869));
    InMux I__945 (
            .O(N__5874),
            .I(N__5866));
    LocalMux I__944 (
            .O(N__5869),
            .I(N__5861));
    LocalMux I__943 (
            .O(N__5866),
            .I(N__5861));
    Span4Mux_v I__942 (
            .O(N__5861),
            .I(N__5858));
    Sp12to4 I__941 (
            .O(N__5858),
            .I(N__5855));
    Span12Mux_h I__940 (
            .O(N__5855),
            .I(N__5852));
    Span12Mux_v I__939 (
            .O(N__5852),
            .I(N__5849));
    Odrv12 I__938 (
            .O(N__5849),
            .I(D_in_6));
    CascadeMux I__937 (
            .O(N__5846),
            .I(N__5842));
    CascadeMux I__936 (
            .O(N__5845),
            .I(N__5839));
    InMux I__935 (
            .O(N__5842),
            .I(N__5836));
    InMux I__934 (
            .O(N__5839),
            .I(N__5833));
    LocalMux I__933 (
            .O(N__5836),
            .I(N__5830));
    LocalMux I__932 (
            .O(N__5833),
            .I(BRIDGE_BASE_2));
    Odrv4 I__931 (
            .O(N__5830),
            .I(BRIDGE_BASE_2));
    InMux I__930 (
            .O(N__5825),
            .I(N__5819));
    InMux I__929 (
            .O(N__5824),
            .I(N__5819));
    LocalMux I__928 (
            .O(N__5819),
            .I(N__5814));
    InMux I__927 (
            .O(N__5818),
            .I(N__5811));
    CascadeMux I__926 (
            .O(N__5817),
            .I(N__5805));
    Span4Mux_h I__925 (
            .O(N__5814),
            .I(N__5800));
    LocalMux I__924 (
            .O(N__5811),
            .I(N__5800));
    InMux I__923 (
            .O(N__5810),
            .I(N__5797));
    InMux I__922 (
            .O(N__5809),
            .I(N__5792));
    InMux I__921 (
            .O(N__5808),
            .I(N__5792));
    InMux I__920 (
            .O(N__5805),
            .I(N__5787));
    Span4Mux_h I__919 (
            .O(N__5800),
            .I(N__5782));
    LocalMux I__918 (
            .O(N__5797),
            .I(N__5782));
    LocalMux I__917 (
            .O(N__5792),
            .I(N__5779));
    InMux I__916 (
            .O(N__5791),
            .I(N__5776));
    CascadeMux I__915 (
            .O(N__5790),
            .I(N__5773));
    LocalMux I__914 (
            .O(N__5787),
            .I(N__5770));
    Span4Mux_v I__913 (
            .O(N__5782),
            .I(N__5765));
    Span4Mux_v I__912 (
            .O(N__5779),
            .I(N__5765));
    LocalMux I__911 (
            .O(N__5776),
            .I(N__5762));
    InMux I__910 (
            .O(N__5773),
            .I(N__5759));
    Span12Mux_h I__909 (
            .O(N__5770),
            .I(N__5750));
    Sp12to4 I__908 (
            .O(N__5765),
            .I(N__5750));
    Span12Mux_v I__907 (
            .O(N__5762),
            .I(N__5750));
    LocalMux I__906 (
            .O(N__5759),
            .I(N__5750));
    Odrv12 I__905 (
            .O(N__5750),
            .I(A_c_20));
    InMux I__904 (
            .O(N__5747),
            .I(N__5741));
    InMux I__903 (
            .O(N__5746),
            .I(N__5741));
    LocalMux I__902 (
            .O(N__5741),
            .I(ATA_BASE_4));
    InMux I__901 (
            .O(N__5738),
            .I(N__5732));
    InMux I__900 (
            .O(N__5737),
            .I(N__5725));
    InMux I__899 (
            .O(N__5736),
            .I(N__5725));
    InMux I__898 (
            .O(N__5735),
            .I(N__5725));
    LocalMux I__897 (
            .O(N__5732),
            .I(\U409_AUTOCONFIG.LIDE_CONF_RNIDFPAZ0Z3 ));
    LocalMux I__896 (
            .O(N__5725),
            .I(\U409_AUTOCONFIG.LIDE_CONF_RNIDFPAZ0Z3 ));
    InMux I__895 (
            .O(N__5720),
            .I(N__5714));
    InMux I__894 (
            .O(N__5719),
            .I(N__5714));
    LocalMux I__893 (
            .O(N__5714),
            .I(ATA_BASE_5));
    CascadeMux I__892 (
            .O(N__5711),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ));
    CascadeMux I__891 (
            .O(N__5708),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    InMux I__890 (
            .O(N__5705),
            .I(N__5698));
    InMux I__889 (
            .O(N__5704),
            .I(N__5698));
    InMux I__888 (
            .O(N__5703),
            .I(N__5695));
    LocalMux I__887 (
            .O(N__5698),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ));
    LocalMux I__886 (
            .O(N__5695),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ));
    CascadeMux I__885 (
            .O(N__5690),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_ ));
    InMux I__884 (
            .O(N__5687),
            .I(N__5684));
    LocalMux I__883 (
            .O(N__5684),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5 ));
    IoInMux I__882 (
            .O(N__5681),
            .I(N__5678));
    LocalMux I__881 (
            .O(N__5678),
            .I(N__5675));
    Span12Mux_s8_v I__880 (
            .O(N__5675),
            .I(N__5672));
    Span12Mux_h I__879 (
            .O(N__5672),
            .I(N__5668));
    InMux I__878 (
            .O(N__5671),
            .I(N__5665));
    Odrv12 I__877 (
            .O(N__5668),
            .I(CONFIGENn_c));
    LocalMux I__876 (
            .O(N__5665),
            .I(CONFIGENn_c));
    CascadeMux I__875 (
            .O(N__5660),
            .I(\U409_AUTOCONFIG.STATE_d_2_cascade_ ));
    InMux I__874 (
            .O(N__5657),
            .I(N__5653));
    InMux I__873 (
            .O(N__5656),
            .I(N__5650));
    LocalMux I__872 (
            .O(N__5653),
            .I(N__5646));
    LocalMux I__871 (
            .O(N__5650),
            .I(N__5643));
    InMux I__870 (
            .O(N__5649),
            .I(N__5640));
    Span4Mux_v I__869 (
            .O(N__5646),
            .I(N__5637));
    Span4Mux_v I__868 (
            .O(N__5643),
            .I(N__5634));
    LocalMux I__867 (
            .O(N__5640),
            .I(N__5631));
    Span4Mux_v I__866 (
            .O(N__5637),
            .I(N__5628));
    Span4Mux_v I__865 (
            .O(N__5634),
            .I(N__5625));
    Span12Mux_v I__864 (
            .O(N__5631),
            .I(N__5618));
    Sp12to4 I__863 (
            .O(N__5628),
            .I(N__5618));
    Sp12to4 I__862 (
            .O(N__5625),
            .I(N__5618));
    Odrv12 I__861 (
            .O(N__5618),
            .I(A_c_31));
    InMux I__860 (
            .O(N__5615),
            .I(N__5611));
    InMux I__859 (
            .O(N__5614),
            .I(N__5608));
    LocalMux I__858 (
            .O(N__5611),
            .I(N__5605));
    LocalMux I__857 (
            .O(N__5608),
            .I(N__5602));
    Span4Mux_v I__856 (
            .O(N__5605),
            .I(N__5598));
    Span4Mux_v I__855 (
            .O(N__5602),
            .I(N__5595));
    InMux I__854 (
            .O(N__5601),
            .I(N__5592));
    Span4Mux_v I__853 (
            .O(N__5598),
            .I(N__5589));
    Span4Mux_v I__852 (
            .O(N__5595),
            .I(N__5586));
    LocalMux I__851 (
            .O(N__5592),
            .I(N__5583));
    Span4Mux_h I__850 (
            .O(N__5589),
            .I(N__5580));
    Span4Mux_h I__849 (
            .O(N__5586),
            .I(N__5577));
    Sp12to4 I__848 (
            .O(N__5583),
            .I(N__5574));
    Sp12to4 I__847 (
            .O(N__5580),
            .I(N__5567));
    Sp12to4 I__846 (
            .O(N__5577),
            .I(N__5567));
    Span12Mux_v I__845 (
            .O(N__5574),
            .I(N__5567));
    Odrv12 I__844 (
            .O(N__5567),
            .I(A_c_30));
    CascadeMux I__843 (
            .O(N__5564),
            .I(N__5560));
    InMux I__842 (
            .O(N__5563),
            .I(N__5557));
    InMux I__841 (
            .O(N__5560),
            .I(N__5554));
    LocalMux I__840 (
            .O(N__5557),
            .I(BRIDGE_BASE_3));
    LocalMux I__839 (
            .O(N__5554),
            .I(BRIDGE_BASE_3));
    InMux I__838 (
            .O(N__5549),
            .I(N__5546));
    LocalMux I__837 (
            .O(N__5546),
            .I(N__5541));
    InMux I__836 (
            .O(N__5545),
            .I(N__5538));
    InMux I__835 (
            .O(N__5544),
            .I(N__5535));
    Span4Mux_h I__834 (
            .O(N__5541),
            .I(N__5530));
    LocalMux I__833 (
            .O(N__5538),
            .I(N__5530));
    LocalMux I__832 (
            .O(N__5535),
            .I(N__5525));
    Sp12to4 I__831 (
            .O(N__5530),
            .I(N__5525));
    Span12Mux_v I__830 (
            .O(N__5525),
            .I(N__5522));
    Odrv12 I__829 (
            .O(N__5522),
            .I(A_c_29));
    CascadeMux I__828 (
            .O(N__5519),
            .I(N__5515));
    InMux I__827 (
            .O(N__5518),
            .I(N__5511));
    InMux I__826 (
            .O(N__5515),
            .I(N__5508));
    CascadeMux I__825 (
            .O(N__5514),
            .I(N__5505));
    LocalMux I__824 (
            .O(N__5511),
            .I(N__5500));
    LocalMux I__823 (
            .O(N__5508),
            .I(N__5500));
    InMux I__822 (
            .O(N__5505),
            .I(N__5497));
    Span4Mux_h I__821 (
            .O(N__5500),
            .I(N__5494));
    LocalMux I__820 (
            .O(N__5497),
            .I(N__5491));
    Sp12to4 I__819 (
            .O(N__5494),
            .I(N__5488));
    Span12Mux_v I__818 (
            .O(N__5491),
            .I(N__5485));
    Span12Mux_v I__817 (
            .O(N__5488),
            .I(N__5482));
    Odrv12 I__816 (
            .O(N__5485),
            .I(A_c_28));
    Odrv12 I__815 (
            .O(N__5482),
            .I(A_c_28));
    CascadeMux I__814 (
            .O(N__5477),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2Z0Z_0_cascade_ ));
    InMux I__813 (
            .O(N__5474),
            .I(N__5471));
    LocalMux I__812 (
            .O(N__5471),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_3 ));
    InMux I__811 (
            .O(N__5468),
            .I(N__5465));
    LocalMux I__810 (
            .O(N__5465),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0 ));
    InMux I__809 (
            .O(N__5462),
            .I(N__5458));
    InMux I__808 (
            .O(N__5461),
            .I(N__5455));
    LocalMux I__807 (
            .O(N__5458),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_4 ));
    LocalMux I__806 (
            .O(N__5455),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_4 ));
    CascadeMux I__805 (
            .O(N__5450),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_ ));
    InMux I__804 (
            .O(N__5447),
            .I(N__5444));
    LocalMux I__803 (
            .O(N__5444),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_2_0 ));
    CascadeMux I__802 (
            .O(N__5441),
            .I(N__5438));
    InMux I__801 (
            .O(N__5438),
            .I(N__5434));
    InMux I__800 (
            .O(N__5437),
            .I(N__5431));
    LocalMux I__799 (
            .O(N__5434),
            .I(N__5426));
    LocalMux I__798 (
            .O(N__5431),
            .I(N__5426));
    Span4Mux_v I__797 (
            .O(N__5426),
            .I(N__5423));
    Odrv4 I__796 (
            .O(N__5423),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6 ));
    InMux I__795 (
            .O(N__5420),
            .I(N__5417));
    LocalMux I__794 (
            .O(N__5417),
            .I(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7 ));
    InMux I__793 (
            .O(N__5414),
            .I(N__5411));
    LocalMux I__792 (
            .O(N__5411),
            .I(U409_ADDRESS_DECODE_AUTOVECTOR_8));
    CascadeMux I__791 (
            .O(N__5408),
            .I(U409_ADDRESS_DECODE_AUTOVECTOR_10_cascade_));
    InMux I__790 (
            .O(N__5405),
            .I(N__5402));
    LocalMux I__789 (
            .O(N__5402),
            .I(U409_ADDRESS_DECODE_AUTOVECTOR_9));
    InMux I__788 (
            .O(N__5399),
            .I(N__5396));
    LocalMux I__787 (
            .O(N__5396),
            .I(N__5392));
    InMux I__786 (
            .O(N__5395),
            .I(N__5389));
    Odrv4 I__785 (
            .O(N__5392),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ));
    LocalMux I__784 (
            .O(N__5389),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ));
    CascadeMux I__783 (
            .O(N__5384),
            .I(N__5381));
    InMux I__782 (
            .O(N__5381),
            .I(N__5377));
    InMux I__781 (
            .O(N__5380),
            .I(N__5374));
    LocalMux I__780 (
            .O(N__5377),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ));
    LocalMux I__779 (
            .O(N__5374),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ));
    IoInMux I__778 (
            .O(N__5369),
            .I(N__5366));
    LocalMux I__777 (
            .O(N__5366),
            .I(N__5363));
    Span12Mux_s6_v I__776 (
            .O(N__5363),
            .I(N__5360));
    Odrv12 I__775 (
            .O(N__5360),
            .I(U409_AUTOCONFIG_D_OUT_0_i_1));
    InMux I__774 (
            .O(N__5357),
            .I(N__5353));
    InMux I__773 (
            .O(N__5356),
            .I(N__5350));
    LocalMux I__772 (
            .O(N__5353),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ));
    LocalMux I__771 (
            .O(N__5350),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ));
    InMux I__770 (
            .O(N__5345),
            .I(N__5342));
    LocalMux I__769 (
            .O(N__5342),
            .I(N__5338));
    InMux I__768 (
            .O(N__5341),
            .I(N__5335));
    Odrv4 I__767 (
            .O(N__5338),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2 ));
    LocalMux I__766 (
            .O(N__5335),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2 ));
    IoInMux I__765 (
            .O(N__5330),
            .I(N__5327));
    LocalMux I__764 (
            .O(N__5327),
            .I(N__5324));
    Span12Mux_s7_v I__763 (
            .O(N__5324),
            .I(N__5321));
    Odrv12 I__762 (
            .O(N__5321),
            .I(U409_AUTOCONFIG_D_OUT_0_i_2));
    InMux I__761 (
            .O(N__5318),
            .I(N__5315));
    LocalMux I__760 (
            .O(N__5315),
            .I(N__5311));
    InMux I__759 (
            .O(N__5314),
            .I(N__5308));
    Odrv4 I__758 (
            .O(N__5311),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ));
    LocalMux I__757 (
            .O(N__5308),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ));
    InMux I__756 (
            .O(N__5303),
            .I(N__5300));
    LocalMux I__755 (
            .O(N__5300),
            .I(N__5297));
    Odrv12 I__754 (
            .O(N__5297),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNO_0Z0Z_0 ));
    CascadeMux I__753 (
            .O(N__5294),
            .I(N__5290));
    InMux I__752 (
            .O(N__5293),
            .I(N__5287));
    InMux I__751 (
            .O(N__5290),
            .I(N__5284));
    LocalMux I__750 (
            .O(N__5287),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ));
    LocalMux I__749 (
            .O(N__5284),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ));
    InMux I__748 (
            .O(N__5279),
            .I(N__5276));
    LocalMux I__747 (
            .O(N__5276),
            .I(\U409_AUTOCONFIG.un1_STATE_8_0_0 ));
    InMux I__746 (
            .O(N__5273),
            .I(N__5267));
    InMux I__745 (
            .O(N__5272),
            .I(N__5267));
    LocalMux I__744 (
            .O(N__5267),
            .I(\U409_AUTOCONFIG.STATE4 ));
    InMux I__743 (
            .O(N__5264),
            .I(N__5255));
    InMux I__742 (
            .O(N__5263),
            .I(N__5255));
    InMux I__741 (
            .O(N__5262),
            .I(N__5255));
    LocalMux I__740 (
            .O(N__5255),
            .I(\U409_AUTOCONFIG.un1_STATE_8Z0Z_0 ));
    InMux I__739 (
            .O(N__5252),
            .I(N__5249));
    LocalMux I__738 (
            .O(N__5249),
            .I(N__5246));
    Span4Mux_h I__737 (
            .O(N__5246),
            .I(N__5243));
    Odrv4 I__736 (
            .O(N__5243),
            .I(\U409_AUTOCONFIG.N_248_0 ));
    CascadeMux I__735 (
            .O(N__5240),
            .I(\U409_AUTOCONFIG.un1_STATE_8Z0Z_0_cascade_ ));
    IoInMux I__734 (
            .O(N__5237),
            .I(N__5234));
    LocalMux I__733 (
            .O(N__5234),
            .I(N__5231));
    IoSpan4Mux I__732 (
            .O(N__5231),
            .I(N__5228));
    Span4Mux_s2_h I__731 (
            .O(N__5228),
            .I(N__5225));
    Sp12to4 I__730 (
            .O(N__5225),
            .I(N__5222));
    Span12Mux_s10_h I__729 (
            .O(N__5222),
            .I(N__5219));
    Span12Mux_v I__728 (
            .O(N__5219),
            .I(N__5216));
    Odrv12 I__727 (
            .O(N__5216),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn_i));
    InMux I__726 (
            .O(N__5213),
            .I(N__5210));
    LocalMux I__725 (
            .O(N__5210),
            .I(N__5207));
    Span4Mux_v I__724 (
            .O(N__5207),
            .I(N__5204));
    Sp12to4 I__723 (
            .O(N__5204),
            .I(N__5201));
    Span12Mux_h I__722 (
            .O(N__5201),
            .I(N__5198));
    Odrv12 I__721 (
            .O(N__5198),
            .I(TT_c_1));
    InMux I__720 (
            .O(N__5195),
            .I(N__5192));
    LocalMux I__719 (
            .O(N__5192),
            .I(N__5189));
    Span12Mux_h I__718 (
            .O(N__5189),
            .I(N__5186));
    Span12Mux_v I__717 (
            .O(N__5186),
            .I(N__5183));
    Odrv12 I__716 (
            .O(N__5183),
            .I(TT_c_0));
    IoInMux I__715 (
            .O(N__5180),
            .I(N__5175));
    IoInMux I__714 (
            .O(N__5179),
            .I(N__5172));
    IoInMux I__713 (
            .O(N__5178),
            .I(N__5169));
    LocalMux I__712 (
            .O(N__5175),
            .I(N__5164));
    LocalMux I__711 (
            .O(N__5172),
            .I(N__5164));
    LocalMux I__710 (
            .O(N__5169),
            .I(N__5161));
    Span4Mux_s2_v I__709 (
            .O(N__5164),
            .I(N__5157));
    Span4Mux_s3_v I__708 (
            .O(N__5161),
            .I(N__5154));
    IoInMux I__707 (
            .O(N__5160),
            .I(N__5151));
    Span4Mux_v I__706 (
            .O(N__5157),
            .I(N__5148));
    Span4Mux_h I__705 (
            .O(N__5154),
            .I(N__5145));
    LocalMux I__704 (
            .O(N__5151),
            .I(N__5142));
    Span4Mux_v I__703 (
            .O(N__5148),
            .I(N__5139));
    Sp12to4 I__702 (
            .O(N__5145),
            .I(N__5134));
    Span12Mux_s4_v I__701 (
            .O(N__5142),
            .I(N__5134));
    Odrv4 I__700 (
            .O(N__5139),
            .I(D_1_i));
    Odrv12 I__699 (
            .O(N__5134),
            .I(D_1_i));
    InMux I__698 (
            .O(N__5129),
            .I(N__5126));
    LocalMux I__697 (
            .O(N__5126),
            .I(N__5122));
    InMux I__696 (
            .O(N__5125),
            .I(N__5119));
    Odrv4 I__695 (
            .O(N__5122),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ));
    LocalMux I__694 (
            .O(N__5119),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ));
    IoInMux I__693 (
            .O(N__5114),
            .I(N__5111));
    LocalMux I__692 (
            .O(N__5111),
            .I(N__5108));
    Sp12to4 I__691 (
            .O(N__5108),
            .I(N__5105));
    Span12Mux_v I__690 (
            .O(N__5105),
            .I(N__5102));
    Odrv12 I__689 (
            .O(N__5102),
            .I(U409_AUTOCONFIG_D_OUT_0_i_3));
    CascadeMux I__688 (
            .O(N__5099),
            .I(AUTOCONFIG_SPACE_cascade_));
    InMux I__687 (
            .O(N__5096),
            .I(N__5093));
    LocalMux I__686 (
            .O(N__5093),
            .I(\U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0_a3_0 ));
    CascadeMux I__685 (
            .O(N__5090),
            .I(N__5087));
    InMux I__684 (
            .O(N__5087),
            .I(N__5084));
    LocalMux I__683 (
            .O(N__5084),
            .I(N__5081));
    Span4Mux_v I__682 (
            .O(N__5081),
            .I(N__5077));
    InMux I__681 (
            .O(N__5080),
            .I(N__5074));
    Sp12to4 I__680 (
            .O(N__5077),
            .I(N__5069));
    LocalMux I__679 (
            .O(N__5074),
            .I(N__5069));
    Span12Mux_v I__678 (
            .O(N__5069),
            .I(N__5066));
    Odrv12 I__677 (
            .O(N__5066),
            .I(CPUCONFn_c));
    InMux I__676 (
            .O(N__5063),
            .I(N__5059));
    InMux I__675 (
            .O(N__5062),
            .I(N__5056));
    LocalMux I__674 (
            .O(N__5059),
            .I(\U409_AUTOCONFIG.AC_STARTZ0 ));
    LocalMux I__673 (
            .O(N__5056),
            .I(\U409_AUTOCONFIG.AC_STARTZ0 ));
    CascadeMux I__672 (
            .O(N__5051),
            .I(N__5048));
    InMux I__671 (
            .O(N__5048),
            .I(N__5044));
    InMux I__670 (
            .O(N__5047),
            .I(N__5041));
    LocalMux I__669 (
            .O(N__5044),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ));
    LocalMux I__668 (
            .O(N__5041),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ));
    IoInMux I__667 (
            .O(N__5036),
            .I(N__5033));
    LocalMux I__666 (
            .O(N__5033),
            .I(N__5030));
    Span12Mux_s10_v I__665 (
            .O(N__5030),
            .I(N__5027));
    Odrv12 I__664 (
            .O(N__5027),
            .I(U409_AUTOCONFIG_D_OUT_0_i_0));
    InMux I__663 (
            .O(N__5024),
            .I(N__5021));
    LocalMux I__662 (
            .O(N__5021),
            .I(N__5018));
    Odrv4 I__661 (
            .O(N__5018),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNO_0Z0Z_1 ));
    InMux I__660 (
            .O(N__5015),
            .I(N__5012));
    LocalMux I__659 (
            .O(N__5012),
            .I(N__5009));
    Span4Mux_v I__658 (
            .O(N__5009),
            .I(N__5006));
    Odrv4 I__657 (
            .O(N__5006),
            .I(\U409_AUTOCONFIG.N_265_0 ));
    InMux I__656 (
            .O(N__5003),
            .I(N__4991));
    InMux I__655 (
            .O(N__5002),
            .I(N__4991));
    InMux I__654 (
            .O(N__5001),
            .I(N__4984));
    InMux I__653 (
            .O(N__5000),
            .I(N__4984));
    InMux I__652 (
            .O(N__4999),
            .I(N__4984));
    InMux I__651 (
            .O(N__4998),
            .I(N__4978));
    InMux I__650 (
            .O(N__4997),
            .I(N__4978));
    InMux I__649 (
            .O(N__4996),
            .I(N__4974));
    LocalMux I__648 (
            .O(N__4991),
            .I(N__4966));
    LocalMux I__647 (
            .O(N__4984),
            .I(N__4966));
    InMux I__646 (
            .O(N__4983),
            .I(N__4963));
    LocalMux I__645 (
            .O(N__4978),
            .I(N__4958));
    InMux I__644 (
            .O(N__4977),
            .I(N__4955));
    LocalMux I__643 (
            .O(N__4974),
            .I(N__4952));
    InMux I__642 (
            .O(N__4973),
            .I(N__4945));
    InMux I__641 (
            .O(N__4972),
            .I(N__4945));
    InMux I__640 (
            .O(N__4971),
            .I(N__4945));
    Span4Mux_h I__639 (
            .O(N__4966),
            .I(N__4940));
    LocalMux I__638 (
            .O(N__4963),
            .I(N__4940));
    InMux I__637 (
            .O(N__4962),
            .I(N__4935));
    InMux I__636 (
            .O(N__4961),
            .I(N__4935));
    Span4Mux_v I__635 (
            .O(N__4958),
            .I(N__4930));
    LocalMux I__634 (
            .O(N__4955),
            .I(N__4930));
    Span4Mux_v I__633 (
            .O(N__4952),
            .I(N__4925));
    LocalMux I__632 (
            .O(N__4945),
            .I(N__4925));
    Span4Mux_h I__631 (
            .O(N__4940),
            .I(N__4920));
    LocalMux I__630 (
            .O(N__4935),
            .I(N__4920));
    Span4Mux_v I__629 (
            .O(N__4930),
            .I(N__4917));
    Span4Mux_v I__628 (
            .O(N__4925),
            .I(N__4914));
    Span4Mux_v I__627 (
            .O(N__4920),
            .I(N__4911));
    Sp12to4 I__626 (
            .O(N__4917),
            .I(N__4906));
    Sp12to4 I__625 (
            .O(N__4914),
            .I(N__4906));
    Span4Mux_h I__624 (
            .O(N__4911),
            .I(N__4903));
    Span12Mux_h I__623 (
            .O(N__4906),
            .I(N__4898));
    Sp12to4 I__622 (
            .O(N__4903),
            .I(N__4898));
    Odrv12 I__621 (
            .O(N__4898),
            .I(A_c_2));
    CascadeMux I__620 (
            .O(N__4895),
            .I(\U409_AUTOCONFIG.un1_A_11Z0Z_0_cascade_ ));
    InMux I__619 (
            .O(N__4892),
            .I(N__4889));
    LocalMux I__618 (
            .O(N__4889),
            .I(\U409_AUTOCONFIG.un1_AZ0Z_11 ));
    InMux I__617 (
            .O(N__4886),
            .I(N__4877));
    InMux I__616 (
            .O(N__4885),
            .I(N__4877));
    InMux I__615 (
            .O(N__4884),
            .I(N__4874));
    InMux I__614 (
            .O(N__4883),
            .I(N__4871));
    InMux I__613 (
            .O(N__4882),
            .I(N__4868));
    LocalMux I__612 (
            .O(N__4877),
            .I(N__4863));
    LocalMux I__611 (
            .O(N__4874),
            .I(N__4863));
    LocalMux I__610 (
            .O(N__4871),
            .I(N__4858));
    LocalMux I__609 (
            .O(N__4868),
            .I(N__4858));
    Span4Mux_v I__608 (
            .O(N__4863),
            .I(N__4853));
    Span4Mux_v I__607 (
            .O(N__4858),
            .I(N__4850));
    InMux I__606 (
            .O(N__4857),
            .I(N__4845));
    InMux I__605 (
            .O(N__4856),
            .I(N__4845));
    Sp12to4 I__604 (
            .O(N__4853),
            .I(N__4838));
    Sp12to4 I__603 (
            .O(N__4850),
            .I(N__4838));
    LocalMux I__602 (
            .O(N__4845),
            .I(N__4838));
    Odrv12 I__601 (
            .O(N__4838),
            .I(A_c_6));
    CascadeMux I__600 (
            .O(N__4835),
            .I(N__4831));
    CascadeMux I__599 (
            .O(N__4834),
            .I(N__4827));
    InMux I__598 (
            .O(N__4831),
            .I(N__4820));
    InMux I__597 (
            .O(N__4830),
            .I(N__4815));
    InMux I__596 (
            .O(N__4827),
            .I(N__4815));
    InMux I__595 (
            .O(N__4826),
            .I(N__4809));
    InMux I__594 (
            .O(N__4825),
            .I(N__4809));
    InMux I__593 (
            .O(N__4824),
            .I(N__4806));
    InMux I__592 (
            .O(N__4823),
            .I(N__4803));
    LocalMux I__591 (
            .O(N__4820),
            .I(N__4800));
    LocalMux I__590 (
            .O(N__4815),
            .I(N__4797));
    CascadeMux I__589 (
            .O(N__4814),
            .I(N__4794));
    LocalMux I__588 (
            .O(N__4809),
            .I(N__4791));
    LocalMux I__587 (
            .O(N__4806),
            .I(N__4788));
    LocalMux I__586 (
            .O(N__4803),
            .I(N__4785));
    Span4Mux_v I__585 (
            .O(N__4800),
            .I(N__4778));
    Span4Mux_v I__584 (
            .O(N__4797),
            .I(N__4778));
    InMux I__583 (
            .O(N__4794),
            .I(N__4775));
    Span4Mux_v I__582 (
            .O(N__4791),
            .I(N__4770));
    Span4Mux_v I__581 (
            .O(N__4788),
            .I(N__4770));
    Span4Mux_v I__580 (
            .O(N__4785),
            .I(N__4767));
    InMux I__579 (
            .O(N__4784),
            .I(N__4762));
    InMux I__578 (
            .O(N__4783),
            .I(N__4762));
    Sp12to4 I__577 (
            .O(N__4778),
            .I(N__4751));
    LocalMux I__576 (
            .O(N__4775),
            .I(N__4751));
    Sp12to4 I__575 (
            .O(N__4770),
            .I(N__4751));
    Sp12to4 I__574 (
            .O(N__4767),
            .I(N__4751));
    LocalMux I__573 (
            .O(N__4762),
            .I(N__4751));
    Span12Mux_h I__572 (
            .O(N__4751),
            .I(N__4748));
    Span12Mux_v I__571 (
            .O(N__4748),
            .I(N__4745));
    Odrv12 I__570 (
            .O(N__4745),
            .I(A_c_3));
    InMux I__569 (
            .O(N__4742),
            .I(N__4737));
    InMux I__568 (
            .O(N__4741),
            .I(N__4732));
    InMux I__567 (
            .O(N__4740),
            .I(N__4732));
    LocalMux I__566 (
            .O(N__4737),
            .I(N__4727));
    LocalMux I__565 (
            .O(N__4732),
            .I(N__4724));
    InMux I__564 (
            .O(N__4731),
            .I(N__4721));
    InMux I__563 (
            .O(N__4730),
            .I(N__4718));
    Odrv4 I__562 (
            .O(N__4727),
            .I(\U409_AUTOCONFIG.N_174 ));
    Odrv12 I__561 (
            .O(N__4724),
            .I(\U409_AUTOCONFIG.N_174 ));
    LocalMux I__560 (
            .O(N__4721),
            .I(\U409_AUTOCONFIG.N_174 ));
    LocalMux I__559 (
            .O(N__4718),
            .I(\U409_AUTOCONFIG.N_174 ));
    InMux I__558 (
            .O(N__4709),
            .I(N__4706));
    LocalMux I__557 (
            .O(N__4706),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ));
    InMux I__556 (
            .O(N__4703),
            .I(N__4697));
    InMux I__555 (
            .O(N__4702),
            .I(N__4697));
    LocalMux I__554 (
            .O(N__4697),
            .I(N__4694));
    Odrv12 I__553 (
            .O(N__4694),
            .I(\U409_ADDRESS_DECODE.REG_SPACE_3 ));
    InMux I__552 (
            .O(N__4691),
            .I(N__4685));
    InMux I__551 (
            .O(N__4690),
            .I(N__4685));
    LocalMux I__550 (
            .O(N__4685),
            .I(N__4682));
    Span4Mux_v I__549 (
            .O(N__4682),
            .I(N__4679));
    Sp12to4 I__548 (
            .O(N__4679),
            .I(N__4676));
    Odrv12 I__547 (
            .O(N__4676),
            .I(A_c_25));
    CascadeMux I__546 (
            .O(N__4673),
            .I(\U409_ADDRESS_DECODE.REG_SPACE_3_cascade_ ));
    InMux I__545 (
            .O(N__4670),
            .I(N__4666));
    InMux I__544 (
            .O(N__4669),
            .I(N__4663));
    LocalMux I__543 (
            .O(N__4666),
            .I(N__4660));
    LocalMux I__542 (
            .O(N__4663),
            .I(N__4657));
    Span4Mux_v I__541 (
            .O(N__4660),
            .I(N__4654));
    Span4Mux_v I__540 (
            .O(N__4657),
            .I(N__4651));
    Span4Mux_v I__539 (
            .O(N__4654),
            .I(N__4648));
    Span4Mux_v I__538 (
            .O(N__4651),
            .I(N__4645));
    Sp12to4 I__537 (
            .O(N__4648),
            .I(N__4640));
    Sp12to4 I__536 (
            .O(N__4645),
            .I(N__4640));
    Odrv12 I__535 (
            .O(N__4640),
            .I(A_c_24));
    CascadeMux I__534 (
            .O(N__4637),
            .I(N__4633));
    InMux I__533 (
            .O(N__4636),
            .I(N__4628));
    InMux I__532 (
            .O(N__4633),
            .I(N__4628));
    LocalMux I__531 (
            .O(N__4628),
            .I(N__4625));
    Span12Mux_v I__530 (
            .O(N__4625),
            .I(N__4622));
    Odrv12 I__529 (
            .O(N__4622),
            .I(A_c_27));
    CascadeMux I__528 (
            .O(N__4619),
            .I(N__4616));
    InMux I__527 (
            .O(N__4616),
            .I(N__4610));
    InMux I__526 (
            .O(N__4615),
            .I(N__4610));
    LocalMux I__525 (
            .O(N__4610),
            .I(N__4607));
    Span4Mux_h I__524 (
            .O(N__4607),
            .I(N__4604));
    Sp12to4 I__523 (
            .O(N__4604),
            .I(N__4601));
    Span12Mux_v I__522 (
            .O(N__4601),
            .I(N__4598));
    Odrv12 I__521 (
            .O(N__4598),
            .I(A_c_26));
    InMux I__520 (
            .O(N__4595),
            .I(N__4592));
    LocalMux I__519 (
            .O(N__4592),
            .I(\U409_AUTOCONFIG.N_173 ));
    CascadeMux I__518 (
            .O(N__4589),
            .I(\U409_AUTOCONFIG.N_249_1_cascade_ ));
    InMux I__517 (
            .O(N__4586),
            .I(N__4581));
    InMux I__516 (
            .O(N__4585),
            .I(N__4576));
    InMux I__515 (
            .O(N__4584),
            .I(N__4576));
    LocalMux I__514 (
            .O(N__4581),
            .I(\U409_AUTOCONFIG.N_155_0 ));
    LocalMux I__513 (
            .O(N__4576),
            .I(\U409_AUTOCONFIG.N_155_0 ));
    CascadeMux I__512 (
            .O(N__4571),
            .I(N__4566));
    CascadeMux I__511 (
            .O(N__4570),
            .I(N__4563));
    CascadeMux I__510 (
            .O(N__4569),
            .I(N__4557));
    InMux I__509 (
            .O(N__4566),
            .I(N__4548));
    InMux I__508 (
            .O(N__4563),
            .I(N__4548));
    InMux I__507 (
            .O(N__4562),
            .I(N__4543));
    InMux I__506 (
            .O(N__4561),
            .I(N__4543));
    InMux I__505 (
            .O(N__4560),
            .I(N__4540));
    InMux I__504 (
            .O(N__4557),
            .I(N__4531));
    InMux I__503 (
            .O(N__4556),
            .I(N__4531));
    InMux I__502 (
            .O(N__4555),
            .I(N__4531));
    InMux I__501 (
            .O(N__4554),
            .I(N__4531));
    InMux I__500 (
            .O(N__4553),
            .I(N__4526));
    LocalMux I__499 (
            .O(N__4548),
            .I(N__4521));
    LocalMux I__498 (
            .O(N__4543),
            .I(N__4521));
    LocalMux I__497 (
            .O(N__4540),
            .I(N__4516));
    LocalMux I__496 (
            .O(N__4531),
            .I(N__4516));
    CascadeMux I__495 (
            .O(N__4530),
            .I(N__4513));
    CascadeMux I__494 (
            .O(N__4529),
            .I(N__4510));
    LocalMux I__493 (
            .O(N__4526),
            .I(N__4506));
    Span4Mux_v I__492 (
            .O(N__4521),
            .I(N__4501));
    Span4Mux_v I__491 (
            .O(N__4516),
            .I(N__4498));
    InMux I__490 (
            .O(N__4513),
            .I(N__4495));
    InMux I__489 (
            .O(N__4510),
            .I(N__4492));
    InMux I__488 (
            .O(N__4509),
            .I(N__4489));
    Span4Mux_v I__487 (
            .O(N__4506),
            .I(N__4486));
    InMux I__486 (
            .O(N__4505),
            .I(N__4481));
    InMux I__485 (
            .O(N__4504),
            .I(N__4481));
    Sp12to4 I__484 (
            .O(N__4501),
            .I(N__4466));
    Sp12to4 I__483 (
            .O(N__4498),
            .I(N__4466));
    LocalMux I__482 (
            .O(N__4495),
            .I(N__4466));
    LocalMux I__481 (
            .O(N__4492),
            .I(N__4466));
    LocalMux I__480 (
            .O(N__4489),
            .I(N__4466));
    Sp12to4 I__479 (
            .O(N__4486),
            .I(N__4466));
    LocalMux I__478 (
            .O(N__4481),
            .I(N__4466));
    Odrv12 I__477 (
            .O(N__4466),
            .I(A_c_4));
    CascadeMux I__476 (
            .O(N__4463),
            .I(\U409_AUTOCONFIG.un1_A_19Z0Z_1_cascade_ ));
    IoInMux I__475 (
            .O(N__4460),
            .I(N__4457));
    LocalMux I__474 (
            .O(N__4457),
            .I(N__4454));
    Span12Mux_s2_v I__473 (
            .O(N__4454),
            .I(N__4451));
    Span12Mux_v I__472 (
            .O(N__4451),
            .I(N__4448));
    Span12Mux_h I__471 (
            .O(N__4448),
            .I(N__4445));
    Odrv12 I__470 (
            .O(N__4445),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn_i));
    InMux I__469 (
            .O(N__4442),
            .I(N__4436));
    InMux I__468 (
            .O(N__4441),
            .I(N__4436));
    LocalMux I__467 (
            .O(N__4436),
            .I(N__4433));
    Odrv12 I__466 (
            .O(N__4433),
            .I(\U409_ADDRESS_DECODE.un2_REGSPACEn_0_0 ));
    CascadeMux I__465 (
            .O(N__4430),
            .I(N__4426));
    InMux I__464 (
            .O(N__4429),
            .I(N__4421));
    InMux I__463 (
            .O(N__4426),
            .I(N__4421));
    LocalMux I__462 (
            .O(N__4421),
            .I(N__4418));
    Odrv4 I__461 (
            .O(N__4418),
            .I(\U409_ADDRESS_DECODE.REG_SPACEZ0 ));
    CascadeMux I__460 (
            .O(N__4415),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_ ));
    InMux I__459 (
            .O(N__4412),
            .I(N__4409));
    LocalMux I__458 (
            .O(N__4409),
            .I(\U409_ADDRESS_DECODE.REG_SPACEZ0Z_0 ));
    CascadeMux I__457 (
            .O(N__4406),
            .I(N__4403));
    InMux I__456 (
            .O(N__4403),
            .I(N__4400));
    LocalMux I__455 (
            .O(N__4400),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_0_0 ));
    InMux I__454 (
            .O(N__4397),
            .I(N__4394));
    LocalMux I__453 (
            .O(N__4394),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_1_0 ));
    CascadeMux I__452 (
            .O(N__4391),
            .I(\U409_AUTOCONFIG.N_168_cascade_ ));
    InMux I__451 (
            .O(N__4388),
            .I(N__4385));
    LocalMux I__450 (
            .O(N__4385),
            .I(\U409_AUTOCONFIG.N_167 ));
    CascadeMux I__449 (
            .O(N__4382),
            .I(\U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0_cascade_ ));
    InMux I__448 (
            .O(N__4379),
            .I(N__4370));
    InMux I__447 (
            .O(N__4378),
            .I(N__4370));
    InMux I__446 (
            .O(N__4377),
            .I(N__4370));
    LocalMux I__445 (
            .O(N__4370),
            .I(\U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0 ));
    CascadeMux I__444 (
            .O(N__4367),
            .I(N__4364));
    InMux I__443 (
            .O(N__4364),
            .I(N__4361));
    LocalMux I__442 (
            .O(N__4361),
            .I(N__4358));
    Odrv4 I__441 (
            .O(N__4358),
            .I(\U409_AUTOCONFIG.N_166 ));
    InMux I__440 (
            .O(N__4355),
            .I(N__4352));
    LocalMux I__439 (
            .O(N__4352),
            .I(N__4349));
    Odrv4 I__438 (
            .O(N__4349),
            .I(\U409_AUTOCONFIG.N_213_2 ));
    CascadeMux I__437 (
            .O(N__4346),
            .I(\U409_AUTOCONFIG.N_212_cascade_ ));
    CascadeMux I__436 (
            .O(N__4343),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_3_0_cascade_ ));
    InMux I__435 (
            .O(N__4340),
            .I(N__4337));
    LocalMux I__434 (
            .O(N__4337),
            .I(N__4334));
    Odrv4 I__433 (
            .O(N__4334),
            .I(\U409_AUTOCONFIG.N_165 ));
    CascadeMux I__432 (
            .O(N__4331),
            .I(N__4328));
    InMux I__431 (
            .O(N__4328),
            .I(N__4325));
    LocalMux I__430 (
            .O(N__4325),
            .I(\U409_AUTOCONFIG.un1_A_16Z0Z_2 ));
    InMux I__429 (
            .O(N__4322),
            .I(N__4319));
    LocalMux I__428 (
            .O(N__4319),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_0 ));
    IoInMux I__427 (
            .O(N__4316),
            .I(N__4313));
    LocalMux I__426 (
            .O(N__4313),
            .I(N__4309));
    CascadeMux I__425 (
            .O(N__4312),
            .I(N__4306));
    IoSpan4Mux I__424 (
            .O(N__4309),
            .I(N__4302));
    InMux I__423 (
            .O(N__4306),
            .I(N__4299));
    CascadeMux I__422 (
            .O(N__4305),
            .I(N__4296));
    Span4Mux_s0_h I__421 (
            .O(N__4302),
            .I(N__4293));
    LocalMux I__420 (
            .O(N__4299),
            .I(N__4290));
    InMux I__419 (
            .O(N__4296),
            .I(N__4287));
    Sp12to4 I__418 (
            .O(N__4293),
            .I(N__4284));
    Span4Mux_v I__417 (
            .O(N__4290),
            .I(N__4281));
    LocalMux I__416 (
            .O(N__4287),
            .I(N__4278));
    Span12Mux_v I__415 (
            .O(N__4284),
            .I(N__4275));
    Sp12to4 I__414 (
            .O(N__4281),
            .I(N__4272));
    Span4Mux_h I__413 (
            .O(N__4278),
            .I(N__4269));
    Span12Mux_h I__412 (
            .O(N__4275),
            .I(N__4266));
    Span12Mux_s7_h I__411 (
            .O(N__4272),
            .I(N__4261));
    Sp12to4 I__410 (
            .O(N__4269),
            .I(N__4261));
    Span12Mux_h I__409 (
            .O(N__4266),
            .I(N__4256));
    Span12Mux_v I__408 (
            .O(N__4261),
            .I(N__4256));
    Odrv12 I__407 (
            .O(N__4256),
            .I(A_c_16));
    InMux I__406 (
            .O(N__4253),
            .I(N__4250));
    LocalMux I__405 (
            .O(N__4250),
            .I(\U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0 ));
    CascadeMux I__404 (
            .O(N__4247),
            .I(\U409_AUTOCONFIG.N_167_cascade_ ));
    InMux I__403 (
            .O(N__4244),
            .I(N__4241));
    LocalMux I__402 (
            .O(N__4241),
            .I(N__4238));
    Odrv4 I__401 (
            .O(N__4238),
            .I(\U409_AUTOCONFIG.N_233 ));
    CascadeMux I__400 (
            .O(N__4235),
            .I(\U409_AUTOCONFIG.N_231_cascade_ ));
    InMux I__399 (
            .O(N__4232),
            .I(N__4229));
    LocalMux I__398 (
            .O(N__4229),
            .I(\U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_a5_0_0 ));
    InMux I__397 (
            .O(N__4226),
            .I(N__4223));
    LocalMux I__396 (
            .O(N__4223),
            .I(\U409_AUTOCONFIG.N_212 ));
    CascadeMux I__395 (
            .O(N__4220),
            .I(\U409_AUTOCONFIG.N_213_2_cascade_ ));
    CascadeMux I__394 (
            .O(N__4217),
            .I(\U409_AUTOCONFIG.N_249_cascade_ ));
    InMux I__393 (
            .O(N__4214),
            .I(N__4211));
    LocalMux I__392 (
            .O(N__4211),
            .I(\U409_AUTOCONFIG.N_250_1 ));
    InMux I__391 (
            .O(N__4208),
            .I(N__4205));
    LocalMux I__390 (
            .O(N__4205),
            .I(\U409_AUTOCONFIG.N_249 ));
    CascadeMux I__389 (
            .O(N__4202),
            .I(\U409_AUTOCONFIG.N_250_1_cascade_ ));
    IoInMux I__388 (
            .O(N__4199),
            .I(N__4196));
    LocalMux I__387 (
            .O(N__4196),
            .I(N__4193));
    IoSpan4Mux I__386 (
            .O(N__4193),
            .I(N__4190));
    Span4Mux_s3_h I__385 (
            .O(N__4190),
            .I(N__4187));
    Sp12to4 I__384 (
            .O(N__4187),
            .I(N__4184));
    Span12Mux_h I__383 (
            .O(N__4184),
            .I(N__4181));
    Span12Mux_h I__382 (
            .O(N__4181),
            .I(N__4178));
    Odrv12 I__381 (
            .O(N__4178),
            .I(A_c_15));
    IoInMux I__380 (
            .O(N__4175),
            .I(N__4172));
    LocalMux I__379 (
            .O(N__4172),
            .I(N__4169));
    Span4Mux_s3_h I__378 (
            .O(N__4169),
            .I(N__4166));
    Span4Mux_v I__377 (
            .O(N__4166),
            .I(N__4163));
    Sp12to4 I__376 (
            .O(N__4163),
            .I(N__4160));
    Span12Mux_h I__375 (
            .O(N__4160),
            .I(N__4157));
    Span12Mux_h I__374 (
            .O(N__4157),
            .I(N__4154));
    Odrv12 I__373 (
            .O(N__4154),
            .I(A_c_14));
    ClkMux I__372 (
            .O(N__4151),
            .I(N__4115));
    ClkMux I__371 (
            .O(N__4150),
            .I(N__4115));
    ClkMux I__370 (
            .O(N__4149),
            .I(N__4115));
    ClkMux I__369 (
            .O(N__4148),
            .I(N__4115));
    ClkMux I__368 (
            .O(N__4147),
            .I(N__4115));
    ClkMux I__367 (
            .O(N__4146),
            .I(N__4115));
    ClkMux I__366 (
            .O(N__4145),
            .I(N__4115));
    ClkMux I__365 (
            .O(N__4144),
            .I(N__4115));
    ClkMux I__364 (
            .O(N__4143),
            .I(N__4115));
    ClkMux I__363 (
            .O(N__4142),
            .I(N__4115));
    ClkMux I__362 (
            .O(N__4141),
            .I(N__4115));
    ClkMux I__361 (
            .O(N__4140),
            .I(N__4115));
    GlobalMux I__360 (
            .O(N__4115),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .I(N__4143));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .I(N__4140));
    INV \INVU409_AUTOCONFIG.ATA_BASE_1C  (
            .O(\INVU409_AUTOCONFIG.ATA_BASE_1C_net ),
            .I(N__7943));
    INV \INVU409_TRANSFER_ACK.TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .I(N__4149));
    INV \INVU409_TRANSFER_ACK.TACK_OUTnC  (
            .O(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .I(N__4146));
    INV \INVU409_TRANSFER_ACK.ROMENnC  (
            .O(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .I(N__4144));
    INV \INVU409_TRANSFER_ACK.LASTCLK_0C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .I(N__4142));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__4141));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .I(N__4151));
    INV \INVU409_AUTOCONFIG.LIDE_CONFC  (
            .O(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .I(N__7949));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .I(N__4148));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .I(N__4145));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .I(N__4150));
    INV \INVU409_AUTOCONFIG.ATA_BASE_6C  (
            .O(\INVU409_AUTOCONFIG.ATA_BASE_6C_net ),
            .I(N__7948));
    INV \INVU409_AUTOCONFIG.AC_TACKC  (
            .O(\INVU409_AUTOCONFIG.AC_TACKC_net ),
            .I(N__7951));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .I(N__4147));
    INV \INVU409_AUTOCONFIG.STATE_1C  (
            .O(\INVU409_AUTOCONFIG.STATE_1C_net ),
            .I(N__7956));
    INV \INVU409_AUTOCONFIG.BRIDGE_BASE_3C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net ),
            .I(N__7950));
    INV \INVU409_AUTOCONFIG.LIDE_OUT_1C  (
            .O(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .I(N__7955));
    INV \INVU409_AUTOCONFIG.BRIDGE_OUT_0C  (
            .O(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .I(N__7964));
    defparam IN_MUX_bfv_13_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_6_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_15_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_6_0_));
    defparam IN_MUX_bfv_15_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_7_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_15_7_0_));
    defparam IN_MUX_bfv_15_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_4_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__8900),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_a5_0_2_LC_3_11_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_a5_0_2_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_a5_0_2_LC_3_11_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_a5_0_2_LC_3_11_2  (
            .in0(N__4823),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4983),
            .lcout(\U409_AUTOCONFIG.N_213_2 ),
            .ltout(\U409_AUTOCONFIG.N_213_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_3_1_LC_3_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_3_1_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_3_1_LC_3_11_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_3_1_LC_3_11_3  (
            .in0(N__7062),
            .in1(N__4553),
            .in2(N__4220),
            .in3(N__6120),
            .lcout(\U409_AUTOCONFIG.N_233 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_141_i_a4_LC_3_12_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_141_i_a4_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_141_i_a4_LC_3_12_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_141_i_a4_LC_3_12_1  (
            .in0(N__6161),
            .in1(N__4505),
            .in2(N__7061),
            .in3(N__4962),
            .lcout(\U409_AUTOCONFIG.N_249 ),
            .ltout(\U409_AUTOCONFIG.N_249_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_3_12_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_3_12_2 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_3_12_2  (
            .in0(N__4784),
            .in1(N__4214),
            .in2(N__4217),
            .in3(N__7032),
            .lcout(\U409_AUTOCONFIG.N_265_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_2_0_LC_3_12_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_2_0_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_2_0_LC_3_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_2_0_LC_3_12_3  (
            .in0(_gnd_net_),
            .in1(N__4961),
            .in2(_gnd_net_),
            .in3(N__4504),
            .lcout(\U409_AUTOCONFIG.N_250_1 ),
            .ltout(\U409_AUTOCONFIG.N_250_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_3_12_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_3_12_4 .LUT_INIT=16'b0011001100100011;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_3_12_4  (
            .in0(N__4783),
            .in1(N__4208),
            .in2(N__4202),
            .in3(N__7031),
            .lcout(\U409_AUTOCONFIG.N_248_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_3_12_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_3_12_7 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_3_12_7  (
            .in0(N__4253),
            .in1(N__6492),
            .in2(N__5790),
            .in3(N__6398),
            .lcout(\U409_ADDRESS_DECODE.un2_REGSPACEn_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_3_13_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_3_13_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_3_13_7  (
            .in0(N__7441),
            .in1(N__7358),
            .in2(_gnd_net_),
            .in3(N__8450),
            .lcout(\U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.REG_SPACE_0_LC_5_8_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.REG_SPACE_0_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.REG_SPACE_0_LC_5_8_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.REG_SPACE_0_LC_5_8_2  (
            .in0(N__6475),
            .in1(N__5818),
            .in2(_gnd_net_),
            .in3(N__6915),
            .lcout(\U409_ADDRESS_DECODE.REG_SPACEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_2_LC_5_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_2_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_2_LC_5_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_2_LC_5_10_0  (
            .in0(N__4742),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4226),
            .lcout(\U409_AUTOCONFIG.N_167 ),
            .ltout(\U409_AUTOCONFIG.N_167_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_10_1 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_10_1  (
            .in0(N__4340),
            .in1(N__4560),
            .in2(N__4247),
            .in3(N__4996),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_5_10_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_5_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_5_10_5  (
            .in0(N__6476),
            .in1(N__6362),
            .in2(N__4312),
            .in3(N__6926),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_11_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_11_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_11_1  (
            .in0(N__4999),
            .in1(N__4825),
            .in2(_gnd_net_),
            .in3(N__4555),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_a5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_11_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_11_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_11_2  (
            .in0(N__4556),
            .in1(N__5000),
            .in2(N__6148),
            .in3(N__7064),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.N_231_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_5_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_5_11_3 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_5_11_3  (
            .in0(N__7063),
            .in1(N__4244),
            .in2(N__4235),
            .in3(N__4232),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_85_i_a4_LC_5_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_85_i_a4_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_85_i_a4_LC_5_11_4 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_85_i_a4_LC_5_11_4  (
            .in0(N__4826),
            .in1(N__5001),
            .in2(N__4569),
            .in3(N__7065),
            .lcout(\U409_AUTOCONFIG.N_212 ),
            .ltout(\U409_AUTOCONFIG.N_212_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_5_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_5_11_5 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_5_11_5  (
            .in0(N__4355),
            .in1(N__6124),
            .in2(N__4346),
            .in3(N__4554),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_12_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_12_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_12_1  (
            .in0(N__7066),
            .in1(N__4731),
            .in2(_gnd_net_),
            .in3(N__4971),
            .lcout(\U409_AUTOCONFIG.N_166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_5_12_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_5_12_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_5_12_2  (
            .in0(N__4972),
            .in1(N__6165),
            .in2(N__4814),
            .in3(N__7067),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_5_12_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_5_12_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_5_12_3  (
            .in0(N__4882),
            .in1(N__6225),
            .in2(N__4343),
            .in3(N__4509),
            .lcout(\U409_AUTOCONFIG.N_165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_16_2_LC_5_12_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_16_2_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_16_2_LC_5_12_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_AUTOCONFIG.un1_A_16_2_LC_5_12_5  (
            .in0(N__6166),
            .in1(N__6226),
            .in2(N__4529),
            .in3(N__4973),
            .lcout(\U409_AUTOCONFIG.un1_A_16Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_16_LC_5_13_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_16_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_16_LC_5_13_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_AUTOCONFIG.un1_A_16_LC_5_13_4  (
            .in0(N__4883),
            .in1(N__4824),
            .in2(N__4331),
            .in3(N__7016),
            .lcout(\U409_AUTOCONFIG.un1_AZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_6_LC_5_14_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_6_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_6_LC_5_14_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_6_LC_5_14_0  (
            .in0(N__5545),
            .in1(N__4322),
            .in2(N__5519),
            .in3(N__5601),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_LC_5_14_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_LC_5_14_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(N__5656),
            .in2(_gnd_net_),
            .in3(N__4669),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_6_9_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_6_9_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_6_9_2  (
            .in0(N__4702),
            .in1(N__8825),
            .in2(N__4305),
            .in3(N__5810),
            .lcout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.REG_SPACE_LC_6_9_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.REG_SPACE_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.REG_SPACE_LC_6_9_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.REG_SPACE_LC_6_9_6  (
            .in0(N__4703),
            .in1(N__4412),
            .in2(N__8472),
            .in3(N__6391),
            .lcout(\U409_ADDRESS_DECODE.REG_SPACEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_6_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_6_10_0 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_6_10_0  (
            .in0(N__4397),
            .in1(N__5047),
            .in2(N__4406),
            .in3(N__4377),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_6_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_6_10_1 .LUT_INIT=16'b1111101100000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_6_10_1  (
            .in0(N__4998),
            .in1(N__4741),
            .in2(N__4571),
            .in3(N__4585),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_6_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_6_10_3 .LUT_INIT=16'b1000010000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_6_10_3  (
            .in0(N__4997),
            .in1(N__4740),
            .in2(N__4570),
            .in3(N__7069),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.N_168_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_6_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_6_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_6_10_4 .LUT_INIT=16'b1010101000001100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_6_10_4  (
            .in0(N__5125),
            .in1(N__10919),
            .in2(N__4391),
            .in3(N__4379),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_RNI10V92_LC_6_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_RNI10V92_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.AC_START_RNI10V92_LC_6_10_5 .LUT_INIT=16'b1010001010101010;
    LogicCell40 \U409_AUTOCONFIG.AC_START_RNI10V92_LC_6_10_5  (
            .in0(N__10918),
            .in1(N__5096),
            .in2(N__5090),
            .in3(N__5063),
            .lcout(\U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0 ),
            .ltout(\U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_6_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_6_10_6 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_6_10_6  (
            .in0(N__4388),
            .in1(N__4586),
            .in2(N__4382),
            .in3(N__5341),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_6_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_6_10_7 .LUT_INIT=16'b1010111000000100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_6_10_7  (
            .in0(N__4378),
            .in1(N__4584),
            .in2(N__4367),
            .in3(N__5395),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_3_0_LC_6_11_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_3_0_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_3_0_LC_6_11_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_3_0_LC_6_11_2  (
            .in0(N__6221),
            .in1(N__4857),
            .in2(_gnd_net_),
            .in3(N__6149),
            .lcout(\U409_AUTOCONFIG.N_173 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.ATA_BASE11_1_LC_6_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE11_1_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.ATA_BASE11_1_LC_6_11_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE11_1_LC_6_11_4  (
            .in0(N__4561),
            .in1(N__4856),
            .in2(N__4835),
            .in3(N__5002),
            .lcout(\U409_AUTOCONFIG.ATA_BASE11Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_6_2_LC_6_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_6_2_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_6_2_LC_6_11_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_AUTOCONFIG.un1_A_6_2_LC_6_11_5  (
            .in0(N__5003),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4562),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.N_249_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_o3_0_LC_6_11_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_o3_0_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_o3_0_LC_6_11_6 .LUT_INIT=16'b1100110001001100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_o3_0_LC_6_11_6  (
            .in0(N__4595),
            .in1(N__10917),
            .in2(N__4589),
            .in3(N__7068),
            .lcout(\U409_AUTOCONFIG.N_155_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_19_1_LC_6_12_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_19_1_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_19_1_LC_6_12_0 .LUT_INIT=16'b1111111111101101;
    LogicCell40 \U409_AUTOCONFIG.un1_A_19_1_LC_6_12_0  (
            .in0(N__6158),
            .in1(N__6222),
            .in2(N__4530),
            .in3(N__4884),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.un1_A_19Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_STATE_8_0_LC_6_12_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_STATE_8_0_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_STATE_8_0_LC_6_12_1 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \U409_AUTOCONFIG.un1_STATE_8_0_LC_6_12_1  (
            .in0(N__4892),
            .in1(N__4730),
            .in2(N__4463),
            .in3(N__8252),
            .lcout(\U409_AUTOCONFIG.un1_STATE_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_1_LC_6_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_1_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_1_LC_6_12_2 .LUT_INIT=16'b0000100010000000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_1_LC_6_12_2  (
            .in0(N__5980),
            .in1(N__5925),
            .in2(N__7639),
            .in3(N__7600),
            .lcout(U409_ADDRESS_DECODE_ROMEN_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_12_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_12_3 .LUT_INIT=16'b0011111110111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_12_3  (
            .in0(N__4442),
            .in1(N__5982),
            .in2(N__5939),
            .in3(N__4429),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_12_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_12_4 .LUT_INIT=16'b1010001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_12_4  (
            .in0(N__5981),
            .in1(N__4441),
            .in2(N__4430),
            .in3(N__5926),
            .lcout(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_12_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_12_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_12_6  (
            .in0(N__7632),
            .in1(N__7370),
            .in2(_gnd_net_),
            .in3(N__7599),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ),
            .ltout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_6_12_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_6_12_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_6_12_7  (
            .in0(N__7476),
            .in1(N__5924),
            .in2(N__4415),
            .in3(N__5979),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACE_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_11_0_LC_6_13_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_11_0_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_11_0_LC_6_13_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_AUTOCONFIG.un1_A_11_0_LC_6_13_0  (
            .in0(N__4886),
            .in1(N__7024),
            .in2(_gnd_net_),
            .in3(N__6224),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.un1_A_11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_11_LC_6_13_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_11_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_11_LC_6_13_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_AUTOCONFIG.un1_A_11_LC_6_13_1  (
            .in0(N__4830),
            .in1(N__4977),
            .in2(N__4895),
            .in3(N__6160),
            .lcout(\U409_AUTOCONFIG.un1_AZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_0_0_LC_6_13_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_0_0_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_0_0_LC_6_13_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a2_0_0_LC_6_13_3  (
            .in0(N__6223),
            .in1(N__4885),
            .in2(N__4834),
            .in3(N__6159),
            .lcout(\U409_AUTOCONFIG.N_174 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_4_LC_6_13_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_4_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_4_LC_6_13_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_4_LC_6_13_7  (
            .in0(N__5791),
            .in1(N__4709),
            .in2(N__7480),
            .in3(N__6943),
            .lcout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_6_14_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_6_14_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_6_14_2  (
            .in0(N__10933),
            .in1(N__4636),
            .in2(N__4619),
            .in3(N__4691),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_6_14_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_6_14_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_6_14_3  (
            .in0(N__7354),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7454),
            .lcout(\U409_ADDRESS_DECODE.REG_SPACE_3 ),
            .ltout(\U409_ADDRESS_DECODE.REG_SPACE_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_6_14_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_6_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_6_14_4  (
            .in0(N__5437),
            .in1(N__4690),
            .in2(N__4673),
            .in3(N__4670),
            .lcout(U409_ADDRESS_DECODE_AUTOVECTOR_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_6_14_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_6_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_6_14_7  (
            .in0(N__5544),
            .in1(N__5518),
            .in2(N__4637),
            .in3(N__4615),
            .lcout(U409_ADDRESS_DECODE_AUTOVECTOR_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_8_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_8_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.D_1_i_LC_7_8_3  (
            .in0(N__9070),
            .in1(N__9028),
            .in2(_gnd_net_),
            .in3(N__8261),
            .lcout(D_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIG8DB1_3_LC_7_8_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIG8DB1_3_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIG8DB1_3_LC_7_8_4 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIG8DB1_3_LC_7_8_4  (
            .in0(N__5129),
            .in1(N__5318),
            .in2(N__8360),
            .in3(N__6653),
            .lcout(U409_AUTOCONFIG_D_OUT_0_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_7_9_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_7_9_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_7_9_7  (
            .in0(N__8491),
            .in1(N__6496),
            .in2(N__6402),
            .in3(N__6936),
            .lcout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_7_10_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_7_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__9069),
            .in2(_gnd_net_),
            .in3(N__9027),
            .lcout(),
            .ltout(AUTOCONFIG_SPACE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_LC_7_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_START_LC_7_10_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_AUTOCONFIG.AC_START_LC_7_10_2  (
            .in0(N__7245),
            .in1(N__10888),
            .in2(N__5099),
            .in3(N__8350),
            .lcout(\U409_AUTOCONFIG.AC_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7963),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIBIND1_0_LC_7_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIBIND1_0_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIBIND1_0_LC_7_10_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIBIND1_0_LC_7_10_3  (
            .in0(N__8253),
            .in1(N__6076),
            .in2(_gnd_net_),
            .in3(N__6026),
            .lcout(\U409_AUTOCONFIG.un1_BRIDGE_OUT_8_sqmuxa_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_RNI04BC_LC_7_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_RNI04BC_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.AC_START_RNI04BC_LC_7_10_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_AUTOCONFIG.AC_START_RNI04BC_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(N__5080),
            .in2(_gnd_net_),
            .in3(N__5062),
            .lcout(\U409_AUTOCONFIG.STATE4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIA2DB1_0_LC_7_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIA2DB1_0_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIA2DB1_0_LC_7_10_7 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIA2DB1_0_LC_7_10_7  (
            .in0(N__8351),
            .in1(N__5293),
            .in2(N__5051),
            .in3(N__6652),
            .lcout(U409_AUTOCONFIG_D_OUT_0_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_7_11_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_7_11_1 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_1_LC_7_11_1  (
            .in0(N__5024),
            .in1(N__5380),
            .in2(N__10915),
            .in3(N__5263),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_11_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_11_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_11_2 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_11_2  (
            .in0(N__5264),
            .in1(N__5015),
            .in2(N__10929),
            .in3(N__5314),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_0_LC_7_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_0_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.STATE_0_LC_7_11_3 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \U409_AUTOCONFIG.STATE_0_LC_7_11_3  (
            .in0(N__5273),
            .in1(N__6031),
            .in2(N__10916),
            .in3(N__6078),
            .lcout(\U409_AUTOCONFIG.STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_7_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_7_11_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_7_11_5 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_0_LC_7_11_5  (
            .in0(N__10889),
            .in1(N__5303),
            .in2(N__5294),
            .in3(N__5262),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIILDD3_0_LC_7_11_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIILDD3_0_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIILDD3_0_LC_7_11_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIILDD3_0_LC_7_11_6  (
            .in0(N__6077),
            .in1(N__5279),
            .in2(N__6037),
            .in3(N__5272),
            .lcout(\U409_AUTOCONFIG.un1_STATE_8Z0Z_0 ),
            .ltout(\U409_AUTOCONFIG.un1_STATE_8Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_7_11_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_7_11_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_2_LC_7_11_7  (
            .in0(N__10893),
            .in1(N__5252),
            .in2(N__5240),
            .in3(N__5356),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_7_12_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_7_12_3 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_7_12_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_7_12_3  (
            .in0(N__8053),
            .in1(N__8117),
            .in2(N__5564),
            .in3(N__6545),
            .lcout(BRIDGE_BASE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net ),
            .ce(),
            .sr(N__8573));
    defparam \U409_AUTOCONFIG.ATA_BASE_7_LC_7_12_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_7_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_7_LC_7_12_4 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_7_LC_7_12_4  (
            .in0(N__8116),
            .in1(N__5738),
            .in2(N__8054),
            .in3(N__7114),
            .lcout(ATA_BASE_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.BRIDGE_BASE_3C_net ),
            .ce(),
            .sr(N__8573));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_7_12_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_7_12_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_7_12_5  (
            .in0(N__5462),
            .in1(N__5941),
            .in2(N__5989),
            .in3(N__5468),
            .lcout(U409_ADDRESS_DECODE_un1_RTC_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_7_13_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_7_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_7_13_0  (
            .in0(N__5474),
            .in1(N__5213),
            .in2(N__10934),
            .in3(N__5195),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_3_LC_7_13_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_3_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_3_LC_7_13_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_3_LC_7_13_3  (
            .in0(N__5808),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8473),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACE_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_7_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_7_13_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_7_13_4  (
            .in0(N__8475),
            .in1(N__6497),
            .in2(_gnd_net_),
            .in3(N__6403),
            .lcout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0 ),
            .ltout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_7_13_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_7_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_7_13_5  (
            .in0(N__5940),
            .in1(N__5461),
            .in2(N__5450),
            .in3(N__5972),
            .lcout(U409_ADDRESS_DECODE_un1_RTC_ENn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_13_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_13_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_13_7  (
            .in0(N__5809),
            .in1(N__5447),
            .in2(N__5441),
            .in3(N__8474),
            .lcout(CIA_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_7_14_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_7_14_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_7_14_2  (
            .in0(N__5657),
            .in1(N__5420),
            .in2(_gnd_net_),
            .in3(N__5614),
            .lcout(),
            .ltout(U409_ADDRESS_DECODE_AUTOVECTOR_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_AUTOVECTOR_LC_7_14_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_AUTOVECTOR_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_AUTOVECTOR_LC_7_14_3 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \U409_TRANSFER_ACK.un1_AUTOVECTOR_LC_7_14_3  (
            .in0(N__5414),
            .in1(N__6874),
            .in2(N__5408),
            .in3(N__5405),
            .lcout(\U409_TRANSFER_ACK.un1_AUTOVECTOR_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIC4DB1_1_LC_8_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIC4DB1_1_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIC4DB1_1_LC_8_10_3 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIC4DB1_1_LC_8_10_3  (
            .in0(N__5399),
            .in1(N__6650),
            .in2(N__5384),
            .in3(N__8352),
            .lcout(U409_AUTOCONFIG_D_OUT_0_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIE6DB1_2_LC_8_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIE6DB1_2_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIE6DB1_2_LC_8_10_4 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIE6DB1_2_LC_8_10_4  (
            .in0(N__6651),
            .in1(N__5357),
            .in2(N__8359),
            .in3(N__5345),
            .lcout(U409_AUTOCONFIG_D_OUT_0_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_1_LC_8_10_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_1_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.STATE_1_LC_8_10_7 .LUT_INIT=16'b0001000011000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_1_LC_8_10_7  (
            .in0(N__8259),
            .in1(N__6079),
            .in2(N__10914),
            .in3(N__6032),
            .lcout(\U409_AUTOCONFIG.STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_8_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_8_11_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__6074),
            .in2(_gnd_net_),
            .in3(N__6027),
            .lcout(\U409_AUTOCONFIG.STATE_d_2 ),
            .ltout(\U409_AUTOCONFIG.STATE_d_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_LC_8_11_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_LC_8_11_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_LC_8_11_6  (
            .in0(N__6681),
            .in1(_gnd_net_),
            .in2(N__5660),
            .in3(N__6631),
            .lcout(\U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_2_LC_8_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_2_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_2_LC_8_12_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_2_LC_8_12_1  (
            .in0(N__5649),
            .in1(N__5615),
            .in2(N__5845),
            .in3(N__5563),
            .lcout(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIDFPA3_LC_8_12_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIDFPA3_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIDFPA3_LC_8_12_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIDFPA3_LC_8_12_4  (
            .in0(N__7070),
            .in1(N__7082),
            .in2(_gnd_net_),
            .in3(N__6646),
            .lcout(\U409_AUTOCONFIG.LIDE_CONF_RNIDFPAZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_1_LC_8_13_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_1_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_1_LC_8_13_4 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_1_LC_8_13_4  (
            .in0(N__6515),
            .in1(N__5549),
            .in2(N__5514),
            .in3(N__6566),
            .lcout(\U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_0_LC_9_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_0_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_0_LC_9_8_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_0_LC_9_8_3  (
            .in0(N__5824),
            .in1(N__8492),
            .in2(_gnd_net_),
            .in3(N__6477),
            .lcout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2_0_LC_9_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2_0_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2_0_LC_9_8_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2_0_LC_9_8_6  (
            .in0(N__6478),
            .in1(N__7463),
            .in2(_gnd_net_),
            .in3(N__5825),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_9_8_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_9_8_7 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_9_8_7  (
            .in0(N__7313),
            .in1(N__7386),
            .in2(N__5477),
            .in3(N__8493),
            .lcout(\U409_TRANSFER_ACK.N_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_9_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_9_9_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_9_9_0 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_9_9_0  (
            .in0(N__6292),
            .in1(N__5687),
            .in2(N__6823),
            .in3(N__6316),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__9131));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_9_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_9_9_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_9_9_1  (
            .in0(N__6314),
            .in1(N__6291),
            .in2(N__6248),
            .in3(N__6725),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_6_LC_9_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_6_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_6_LC_9_9_2 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_6_LC_9_9_2  (
            .in0(N__7999),
            .in1(N__7252),
            .in2(N__5711),
            .in3(N__6262),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_9_3 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_9_3 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_9_3  (
            .in0(N__6315),
            .in1(N__5704),
            .in2(N__5708),
            .in3(N__6769),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__9131));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_9_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_9_9_4 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_9_9_4  (
            .in0(N__5705),
            .in1(N__6326),
            .in2(N__6822),
            .in3(N__6740),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__9131));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_9_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_9_9_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_9_9_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_9_9_5  (
            .in0(N__5703),
            .in1(N__6768),
            .in2(_gnd_net_),
            .in3(N__6811),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__9131));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_1_LC_9_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_1_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_1_LC_9_9_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_1_LC_9_9_6  (
            .in0(N__6719),
            .in1(N__7706),
            .in2(N__6794),
            .in3(N__7675),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_6_LC_9_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_6_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_6_LC_9_9_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_6_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5690),
            .in3(N__6767),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_TACK_LC_9_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_TACK_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_TACK_LC_9_10_4 .LUT_INIT=16'b1111111010100000;
    LogicCell40 \U409_AUTOCONFIG.AC_TACK_LC_9_10_4  (
            .in0(N__6080),
            .in1(N__8260),
            .in2(N__7792),
            .in3(N__6038),
            .lcout(AC_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.AC_TACKC_net ),
            .ce(),
            .sr(N__8574));
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_9_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_9_10_5 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_9_10_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_AUTOCONFIG.CONFIGENn_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__5671),
            .in2(_gnd_net_),
            .in3(N__6543),
            .lcout(CONFIGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.AC_TACKC_net ),
            .ce(),
            .sr(N__8574));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0EA21_LC_9_11_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0EA21_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0EA21_LC_9_11_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNI0EA21_LC_9_11_0  (
            .in0(N__6230),
            .in1(N__6176),
            .in2(N__6167),
            .in3(N__6616),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.ATA_BASE11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIDSPQ2_0_LC_9_11_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIDSPQ2_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIDSPQ2_0_LC_9_11_1 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIDSPQ2_0_LC_9_11_1  (
            .in0(N__6682),
            .in1(N__6075),
            .in2(N__6041),
            .in3(N__6033),
            .lcout(\U409_AUTOCONFIG.un1_STATE_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_0_LC_9_12_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_0_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_0_LC_9_12_0 .LUT_INIT=16'b1000000000001000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_0_LC_9_12_0  (
            .in0(N__5990),
            .in1(N__5942),
            .in2(N__7462),
            .in3(N__5887),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.ATA_BASE_6_LC_9_12_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_6_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_6_LC_9_12_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_6_LC_9_12_1  (
            .in0(N__5888),
            .in1(N__5877),
            .in2(N__8115),
            .in3(N__5737),
            .lcout(ATA_BASE_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_6C_net ),
            .ce(),
            .sr(N__8570));
    defparam \U409_AUTOCONFIG.ATA_BASE_2_LC_9_12_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_2_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_2_LC_9_12_3 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_2_LC_9_12_3  (
            .in0(N__8097),
            .in1(N__8130),
            .in2(N__5879),
            .in3(N__7130),
            .lcout(ATA_BASE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_6C_net ),
            .ce(),
            .sr(N__8570));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_12_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_12_4 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_12_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_12_4  (
            .in0(N__5878),
            .in1(N__8107),
            .in2(N__5846),
            .in3(N__6544),
            .lcout(BRIDGE_BASE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_6C_net ),
            .ce(),
            .sr(N__8570));
    defparam \U409_AUTOCONFIG.ATA_BASE_4_LC_9_12_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_4_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_4_LC_9_12_5 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_4_LC_9_12_5  (
            .in0(N__5747),
            .in1(N__6592),
            .in2(N__8113),
            .in3(N__5735),
            .lcout(ATA_BASE_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_6C_net ),
            .ce(),
            .sr(N__8570));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_9_12_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_9_12_6 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_9_12_6  (
            .in0(N__8479),
            .in1(N__5719),
            .in2(N__5817),
            .in3(N__5746),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.ATA_BASE_5_LC_9_12_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_5_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_5_LC_9_12_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_5_LC_9_12_7  (
            .in0(N__5720),
            .in1(N__8190),
            .in2(N__8114),
            .in3(N__5736),
            .lcout(ATA_BASE_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_6C_net ),
            .ce(),
            .sr(N__8570));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_9_13_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_9_13_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_9_13_0 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_9_13_0  (
            .in0(N__6335),
            .in1(N__6838),
            .in2(_gnd_net_),
            .in3(N__6269),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .ce(),
            .sr(N__9127));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_9_14_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_9_14_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_9_14_0  (
            .in0(N__7270),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7235),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_8_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_8_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_8_2  (
            .in0(N__7998),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7256),
            .lcout(\U409_TRANSFER_ACK.N_33_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_7_LC_10_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_7_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_7_LC_10_8_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_7_LC_10_8_3  (
            .in0(N__6293),
            .in1(N__6317),
            .in2(_gnd_net_),
            .in3(N__6766),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_10_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_10_8_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_1_0_LC_10_8_4  (
            .in0(N__8835),
            .in1(N__8854),
            .in2(_gnd_net_),
            .in3(N__8671),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_3_LC_10_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_3_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_3_LC_10_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_3_LC_10_9_0  (
            .in0(N__6789),
            .in1(N__6765),
            .in2(N__7708),
            .in3(N__6313),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_7_LC_10_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_7_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_7_LC_10_9_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_7_LC_10_9_1  (
            .in0(N__6290),
            .in1(N__6739),
            .in2(N__6272),
            .in3(N__6241),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_9_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_9_2 .LUT_INIT=16'b0001010100000101;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_9_2  (
            .in0(N__7702),
            .in1(N__7234),
            .in2(N__6251),
            .in3(N__7997),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__9126));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_1_LC_10_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_1_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_1_LC_10_9_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_1_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__7673),
            .in2(_gnd_net_),
            .in3(N__6713),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_9_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_9_4 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_9_4  (
            .in0(N__7674),
            .in1(_gnd_net_),
            .in2(N__7709),
            .in3(N__6818),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__9126));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_9_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_9_5 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_9_5  (
            .in0(N__7655),
            .in1(N__6790),
            .in2(N__6824),
            .in3(N__6714),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__9126));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_7_LC_10_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_7_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_7_LC_10_9_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_7_LC_10_9_7  (
            .in0(N__6788),
            .in1(N__7698),
            .in2(N__6770),
            .in3(N__6738),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(N__7654),
            .in2(_gnd_net_),
            .in3(N__6718),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__9125));
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_10_11_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_10_11_0 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_LC_10_11_0  (
            .in0(N__6695),
            .in1(N__6686),
            .in2(_gnd_net_),
            .in3(N__6630),
            .lcout(\U409_AUTOCONFIG.LIDE_CONFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__8571));
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_10_11_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_10_11_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_10_11_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U409_AUTOCONFIG.CONFIGURED_LC_10_11_2  (
            .in0(N__6546),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8333),
            .lcout(CONFIGURED),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__8571));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_10_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_10_11_4 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_10_11_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_10_11_4  (
            .in0(N__6547),
            .in1(N__8095),
            .in2(N__6596),
            .in3(N__6559),
            .lcout(BRIDGE_BASE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__8571));
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_10_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_10_11_5 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_10_11_5 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_10_11_5  (
            .in0(N__8096),
            .in1(N__6548),
            .in2(N__8191),
            .in3(N__6508),
            .lcout(BRIDGE_BASE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_CONFC_net ),
            .ce(),
            .sr(N__8571));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_10_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_10_12_1 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_10_12_1  (
            .in0(N__6491),
            .in1(N__8014),
            .in2(N__6404),
            .in3(N__7129),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_5_LC_10_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_5_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_5_LC_10_12_2 .LUT_INIT=16'b0010000000010000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_5_LC_10_12_2  (
            .in0(N__7380),
            .in1(N__6884),
            .in2(N__7118),
            .in3(N__7115),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_10_12_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_10_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_LC_10_12_3  (
            .in0(N__7100),
            .in1(N__7094),
            .in2(N__7088),
            .in3(N__8306),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0 ),
            .ltout(\U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_10_12_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_10_12_4 .LUT_INIT=16'b1010101000100000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_LC_10_12_4  (
            .in0(N__10871),
            .in1(N__8257),
            .in2(N__7085),
            .in3(N__9240),
            .lcout(\U409_ADDRESS_DECODE.ATA_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7947),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIS3FU2_0_LC_10_12_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIS3FU2_0_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIS3FU2_0_LC_10_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIS3FU2_0_LC_10_12_5  (
            .in0(N__7081),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7060),
            .lcout(\U409_AUTOCONFIG.STATE_RNIS3FU2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un2_ATA_SPACE_0_LC_10_13_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un2_ATA_SPACE_0_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un2_ATA_SPACE_0_LC_10_13_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U409_ADDRESS_DECODE.un2_ATA_SPACE_0_LC_10_13_1  (
            .in0(N__6947),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8143),
            .lcout(\U409_ADDRESS_DECODE.un2_ATA_SPACEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_LC_10_13_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_LC_10_13_5 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_LC_10_13_5  (
            .in0(N__9084),
            .in1(N__6878),
            .in2(N__9053),
            .in3(N__9328),
            .lcout(U409_ADDRESS_DECODE_PORTSIZE_0),
            .ltout(U409_ADDRESS_DECODE_PORTSIZE_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNI4345U_LC_10_13_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNI4345U_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNI4345U_LC_10_13_6 .LUT_INIT=16'b1110111110101111;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNI4345U_LC_10_13_6  (
            .in0(N__8539),
            .in1(N__9213),
            .in2(N__6863),
            .in3(N__9241),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_10_13_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_10_13_7 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6839),
            .in3(N__7165),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_14_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_14_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_14_2  (
            .in0(N__7274),
            .in1(N__7236),
            .in2(N__8002),
            .in3(N__7174),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(N__8567));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_14_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_14_4 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_14_4  (
            .in0(N__7181),
            .in1(N__7175),
            .in2(N__8003),
            .in3(N__7166),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(N__8567));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_11_4_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_11_4_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_11_4_1  (
            .in0(N__8000),
            .in1(N__7569),
            .in2(_gnd_net_),
            .in3(N__7555),
            .lcout(\U409_TRANSFER_ACK.N_17_mux ),
            .ltout(\U409_TRANSFER_ACK.N_17_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_4_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_4_2 .LUT_INIT=16'b0001101101011111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_4_2  (
            .in0(N__7540),
            .in1(N__7872),
            .in2(N__7154),
            .in3(N__7889),
            .lcout(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_11_4_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_11_4_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_11_4_3  (
            .in0(_gnd_net_),
            .in1(N__7570),
            .in2(_gnd_net_),
            .in3(N__7556),
            .lcout(\U409_TRANSFER_ACK.N_3_0 ),
            .ltout(\U409_TRANSFER_ACK.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_4_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_4_4 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_4_4  (
            .in0(N__7544),
            .in1(N__7873),
            .in2(N__7151),
            .in3(N__7891),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_4_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_4_5 .LUT_INIT=16'b0000100000101010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_4_5  (
            .in0(N__10816),
            .in1(N__7516),
            .in2(N__7148),
            .in3(N__7145),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_11_4_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_11_4_6 .LUT_INIT=16'b0001000000011111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_11_4_6  (
            .in0(N__7874),
            .in1(N__7890),
            .in2(N__7547),
            .in3(N__7139),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.N_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_4_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_4_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_4_7 .LUT_INIT=16'b0010101000001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_4_7  (
            .in0(N__10817),
            .in1(N__7515),
            .in2(N__7133),
            .in3(N__7545),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_11_5_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_11_5_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_11_5_0  (
            .in0(N__10180),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__8576));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_11_5_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_11_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_11_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7571),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__8576));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_5_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_5_7 .LUT_INIT=16'b0101111100001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_5_7  (
            .in0(N__7546),
            .in1(N__7523),
            .in2(N__7517),
            .in3(N__7810),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_0C_net ),
            .ce(),
            .sr(N__8576));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_0_LC_11_8_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_0_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_0_LC_11_8_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_0_LC_11_8_2  (
            .in0(N__7387),
            .in1(N__8842),
            .in2(_gnd_net_),
            .in3(N__7486),
            .lcout(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_11_8_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_11_8_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_1_LC_11_8_7  (
            .in0(N__8389),
            .in1(N__7499),
            .in2(N__7490),
            .in3(N__7388),
            .lcout(\U409_TRANSFER_ACK.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_LC_11_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_11_9_1 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_11_9_1 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_LC_11_9_1  (
            .in0(N__7285),
            .in1(N__8705),
            .in2(_gnd_net_),
            .in3(N__8774),
            .lcout(ROMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .ce(),
            .sr(N__8572));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_9_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__8730),
            .in2(_gnd_net_),
            .in3(N__8765),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .ce(),
            .sr(N__8572));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_11_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_11_9_4 .LUT_INIT=16'b0110100011001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_11_9_4  (
            .in0(N__8767),
            .in1(N__8673),
            .in2(N__8741),
            .in3(N__8699),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .ce(),
            .sr(N__8572));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_9_5 .LUT_INIT=16'b1101000011110010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_9_5  (
            .in0(N__8639),
            .in1(N__8768),
            .in2(N__7826),
            .in3(N__8737),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .ce(),
            .sr(N__8572));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_9_6 .LUT_INIT=16'b0101101110100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_9_6  (
            .in0(N__8766),
            .in1(N__8672),
            .in2(N__8740),
            .in3(N__8698),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .ce(),
            .sr(N__8572));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_9_7 .LUT_INIT=16'b0011001100100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_9_7  (
            .in0(N__7832),
            .in1(N__8738),
            .in2(N__8794),
            .in3(N__8867),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .ce(),
            .sr(N__8572));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_10_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_10_0  (
            .in0(N__7822),
            .in1(N__7811),
            .in2(N__7796),
            .in3(N__7775),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER6 ),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_10_1 .LUT_INIT=16'b0000000111011101;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_10_1  (
            .in0(N__8627),
            .in1(N__8594),
            .in2(N__7763),
            .in3(N__7722),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_11_10_2 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_11_10_2  (
            .in0(N__7723),
            .in1(_gnd_net_),
            .in2(N__7760),
            .in3(N__10880),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI7S9R_1_LC_11_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI7S9R_1_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI7S9R_1_LC_11_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI7S9R_1_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__7707),
            .in2(_gnd_net_),
            .in3(N__7676),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_1_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_10_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_10_6  (
            .in0(N__8595),
            .in1(N__10879),
            .in2(_gnd_net_),
            .in3(N__8628),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_OUTnC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_11_4 .LUT_INIT=16'b0010000000110000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_11_4  (
            .in0(N__8630),
            .in1(N__8597),
            .in2(N__10913),
            .in3(N__8608),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_11_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_11_12_1 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_11_12_1  (
            .in0(N__7643),
            .in1(N__7604),
            .in2(_gnd_net_),
            .in3(N__8327),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1 ),
            .ltout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_11_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_11_12_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_11_12_2  (
            .in0(N__8300),
            .in1(N__8288),
            .in2(N__8279),
            .in3(N__10884),
            .lcout(U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_11_13_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_11_13_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_11_13_2  (
            .in0(N__8258),
            .in1(N__9091),
            .in2(_gnd_net_),
            .in3(N__9051),
            .lcout(un1_AUTOCONFIG_SPACE),
            .ltout(un1_AUTOCONFIG_SPACE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.ATA_BASE_1_LC_11_13_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_1_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_1_LC_11_13_3 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_1_LC_11_13_3  (
            .in0(N__8192),
            .in1(N__8131),
            .in2(N__8147),
            .in3(N__8144),
            .lcout(ATA_BASE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_1C_net ),
            .ce(),
            .sr(N__8568));
    defparam \U409_AUTOCONFIG.ATA_BASE_3_LC_11_13_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.ATA_BASE_3_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.ATA_BASE_3_LC_11_13_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U409_AUTOCONFIG.ATA_BASE_3_LC_11_13_4  (
            .in0(N__8132),
            .in1(N__8070),
            .in2(N__8038),
            .in3(N__8015),
            .lcout(ATA_BASE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.ATA_BASE_1C_net ),
            .ce(),
            .sr(N__8568));
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_7.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_7.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8001),
            .lcout(GB_BUFFER_CLK40_IN_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_4_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_4_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_4_1  (
            .in0(N__10963),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10793),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__8575));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_4_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7892),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net ),
            .ce(),
            .sr(N__8575));
    defparam \U409_TICK.TICK50_LC_12_6_5 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_12_6_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK50_LC_12_6_5  (
            .in0(N__9836),
            .in1(N__7843),
            .in2(N__9781),
            .in3(N__9884),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10566),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_12_8_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_12_8_6 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_12_8_6  (
            .in0(N__8382),
            .in1(N__8512),
            .in2(_gnd_net_),
            .in3(N__8501),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_12_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_12_9_2 .LUT_INIT=16'b1111111101011010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_12_9_2  (
            .in0(N__8696),
            .in1(_gnd_net_),
            .in2(N__8675),
            .in3(N__8762),
            .lcout(\U409_TRANSFER_ACK.N_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_12_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_12_9_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_12_9_3  (
            .in0(N__8861),
            .in1(N__8663),
            .in2(N__8843),
            .in3(N__8694),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_9_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_9_4  (
            .in0(N__8798),
            .in1(N__8726),
            .in2(N__8777),
            .in3(N__8763),
            .lcout(\U409_TRANSFER_ACK.N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_9_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_9_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_9_5  (
            .in0(N__8764),
            .in1(N__8670),
            .in2(N__8739),
            .in3(N__8697),
            .lcout(\U409_TRANSFER_ACK.N_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_9_6 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_9_6  (
            .in0(N__8695),
            .in1(_gnd_net_),
            .in2(N__8674),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_12_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_12_10_5 .LUT_INIT=16'b0101000011110001;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_LC_12_10_5  (
            .in0(N__8629),
            .in1(N__8609),
            .in2(N__8946),
            .in3(N__8596),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .ce(),
            .sr(N__8569));
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_12_12_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_12_12_3 .LUT_INIT=16'b0101010101010001;
    LogicCell40 \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_12_12_3  (
            .in0(N__8540),
            .in1(N__8519),
            .in2(N__8500),
            .in3(N__8393),
            .lcout(AGNUS_SPACE_0),
            .ltout(AGNUS_SPACE_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_12_12_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_12_12_4 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_12_12_4  (
            .in0(N__10825),
            .in1(_gnd_net_),
            .in2(N__9149),
            .in3(N__9146),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.LV_SPACE_LC_12_13_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.LV_SPACE_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.LV_SPACE_LC_12_13_2 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \U409_ADDRESS_DECODE.LV_SPACE_LC_12_13_2  (
            .in0(N__9092),
            .in1(N__9052),
            .in2(N__8981),
            .in3(N__9224),
            .lcout(BUFENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI2ED4S_LC_12_13_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI2ED4S_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNI2ED4S_LC_12_13_3 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_RNI2ED4S_LC_12_13_3  (
            .in0(N__8990),
            .in1(N__8980),
            .in2(_gnd_net_),
            .in3(N__8947),
            .lcout(TCIn_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_14_2.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_14_2.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_14_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_14_2 (
            .in0(N__10826),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(N__9378),
            .in2(N__9636),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_6_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_13_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_13_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_13_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(N__9412),
            .in2(_gnd_net_),
            .in3(N__8888),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__10564),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_13_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_13_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(N__9571),
            .in2(_gnd_net_),
            .in3(N__8885),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__10564),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3  (
            .in0(_gnd_net_),
            .in1(N__9607),
            .in2(_gnd_net_),
            .in3(N__8882),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_13_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_13_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(N__9649),
            .in2(_gnd_net_),
            .in3(N__9176),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__10564),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9707),
            .in3(N__9173),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_13_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_13_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(N__9256),
            .in2(_gnd_net_),
            .in3(N__9170),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__10564),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(N__9688),
            .in2(_gnd_net_),
            .in3(N__9167),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__9718),
            .in2(_gnd_net_),
            .in3(N__9164),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_13_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_13_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__9274),
            .in2(_gnd_net_),
            .in3(N__9161),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__10565),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_13_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_13_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__9589),
            .in2(_gnd_net_),
            .in3(N__9158),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__10565),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_13_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_13_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__9424),
            .in2(_gnd_net_),
            .in3(N__9155),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__10565),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_13_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_13_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(N__9286),
            .in2(_gnd_net_),
            .in3(N__9152),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__10565),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__9448),
            .in2(_gnd_net_),
            .in3(N__9296),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9668),
            .in3(N__9293),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_13_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_13_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_13_7_7  (
            .in0(_gnd_net_),
            .in1(N__9401),
            .in2(_gnd_net_),
            .in3(N__9290),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10565),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_0  (
            .in0(N__9287),
            .in1(N__9275),
            .in2(N__9263),
            .in3(N__9667),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNI206O6_LC_13_12_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNI206O6_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNI206O6_LC_13_12_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNI206O6_LC_13_12_0  (
            .in0(N__9245),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9220),
            .lcout(U409_ADDRESS_DECODE_un1_ATA_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_14_4_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_14_4_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_14_4_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_14_4_7  (
            .in0(N__9818),
            .in1(N__9883),
            .in2(N__9777),
            .in3(N__10310),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10563),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_14_5_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_14_5_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_14_5_0  (
            .in0(N__10298),
            .in1(N__10631),
            .in2(N__10367),
            .in3(N__10610),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_1_LC_14_5_2 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_1_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_1_LC_14_5_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_CIA.VMA_RNO_1_LC_14_5_2  (
            .in0(N__9999),
            .in1(N__10146),
            .in2(N__10087),
            .in3(N__10126),
            .lcout(),
            .ltout(\U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_14_5_3 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_14_5_3 .LUT_INIT=16'b0010000010000000;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_14_5_3  (
            .in0(N__10027),
            .in1(N__10537),
            .in2(N__9179),
            .in3(N__10509),
            .lcout(),
            .ltout(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_14_5_4 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_14_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_14_5_4 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \U409_CIA.VMA_LC_14_5_4  (
            .in0(N__10510),
            .in1(N__9341),
            .in2(N__9314),
            .in3(N__10950),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9979),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_14_5_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_14_5_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_14_5_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_14_5_6  (
            .in0(N__10349),
            .in1(N__10382),
            .in2(_gnd_net_),
            .in3(N__9944),
            .lcout(\U409_TICK.TICK503_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_14_6_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_14_6_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_14_6_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_14_6_0  (
            .in0(N__9869),
            .in1(N__9815),
            .in2(N__10598),
            .in3(N__9761),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10567),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_14_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_14_6_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_14_6_1  (
            .in0(N__9816),
            .in1(N__9870),
            .in2(N__9775),
            .in3(N__10337),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10567),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_14_6_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_14_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_14_6_2  (
            .in0(N__10328),
            .in1(N__10223),
            .in2(N__10268),
            .in3(N__10652),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_14_6_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_14_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_14_6_3 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_14_6_3  (
            .in0(N__9814),
            .in1(N__9868),
            .in2(N__9311),
            .in3(N__9945),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10567),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_6_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_6_4  (
            .in0(N__10283),
            .in1(N__9923),
            .in2(N__9965),
            .in3(N__10582),
            .lcout(),
            .ltout(\U409_TICK.TICK503_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_14_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_14_6_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_14_6_5  (
            .in0(N__9308),
            .in1(N__10667),
            .in2(N__9302),
            .in3(N__10238),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_14_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_14_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_14_6_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_14_6_6  (
            .in0(N__9817),
            .in1(N__9760),
            .in2(N__9299),
            .in3(N__10619),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10567),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_14_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_14_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_14_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(N__9964),
            .in2(_gnd_net_),
            .in3(N__9946),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10567),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_14_7_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_14_7_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_14_7_0 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_14_7_0  (
            .in0(N__9523),
            .in1(N__9556),
            .in2(N__9637),
            .in3(N__9482),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10568),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_14_7_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_14_7_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_14_7_1  (
            .in0(N__9554),
            .in1(N__9525),
            .in2(N__9493),
            .in3(N__9437),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10568),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_14_7_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_14_7_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_14_7_2  (
            .in0(N__9872),
            .in1(N__9831),
            .in2(N__10253),
            .in3(N__9765),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10568),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_14_7_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_14_7_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_14_7_3  (
            .in0(N__9555),
            .in1(N__9526),
            .in2(N__9494),
            .in3(N__9431),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10568),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_14_7_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_14_7_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_14_7_4  (
            .in0(N__9425),
            .in1(N__9413),
            .in2(N__9383),
            .in3(N__9400),
            .lcout(\U409_TICK.TICK603_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_14_7_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_14_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_14_7_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_14_7_5  (
            .in0(N__9553),
            .in1(N__9524),
            .in2(N__9492),
            .in3(N__9389),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10568),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_14_7_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_14_7_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_14_7_6  (
            .in0(N__9382),
            .in1(_gnd_net_),
            .in2(N__9638),
            .in3(_gnd_net_),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10568),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_14_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_14_7_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_14_7_7  (
            .in0(N__9830),
            .in1(N__9871),
            .in2(N__9776),
            .in3(N__10640),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10568),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_14_8_0 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_14_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_14_8_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK60_LC_14_8_0  (
            .in0(N__9481),
            .in1(N__9352),
            .in2(N__9560),
            .in3(N__9518),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10570),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_14_8_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_14_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_14_8_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_14_8_1  (
            .in0(N__9551),
            .in1(N__9480),
            .in2(N__9527),
            .in3(N__9890),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10570),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_14_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_14_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_14_8_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_14_8_2  (
            .in0(N__9882),
            .in1(N__9832),
            .in2(N__9782),
            .in3(N__10208),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10570),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_8_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_14_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_14_8_3  (
            .in0(N__9719),
            .in1(N__9706),
            .in2(N__9692),
            .in3(N__9449),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_14_8_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_14_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_14_8_4 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_14_8_4  (
            .in0(N__9677),
            .in1(N__9552),
            .in2(N__9671),
            .in3(N__9522),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10570),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_8_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_8_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_8_5  (
            .in0(N__9653),
            .in1(N__9629),
            .in2(_gnd_net_),
            .in3(N__9608),
            .lcout(),
            .ltout(\U409_TICK.TICK603_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_14_8_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_14_8_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_14_8_6  (
            .in0(N__9596),
            .in1(N__9590),
            .in2(N__9578),
            .in3(N__9575),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_14_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_14_8_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_14_8_7  (
            .in0(N__9517),
            .in1(N__9479),
            .in2(N__9458),
            .in3(N__9455),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10570),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_4_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_4_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_4_0  (
            .in0(_gnd_net_),
            .in1(N__10503),
            .in2(N__10127),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_4_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_15_4_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_15_4_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_15_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_15_4_1  (
            .in0(_gnd_net_),
            .in1(N__10145),
            .in2(_gnd_net_),
            .in3(N__9908),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__9980),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_15_4_2 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_15_4_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_15_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_15_4_2  (
            .in0(_gnd_net_),
            .in1(N__9998),
            .in2(_gnd_net_),
            .in3(N__9905),
            .lcout(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_15_4_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_15_4_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_15_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_15_4_3  (
            .in0(_gnd_net_),
            .in1(N__10535),
            .in2(_gnd_net_),
            .in3(N__9902),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__9980),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_15_4_4 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_15_4_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_15_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_15_4_4  (
            .in0(_gnd_net_),
            .in1(N__10082),
            .in2(_gnd_net_),
            .in3(N__9899),
            .lcout(\U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_15_4_5 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_15_4_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_15_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_6_LC_15_4_5  (
            .in0(_gnd_net_),
            .in1(N__10046),
            .in2(_gnd_net_),
            .in3(N__9896),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ),
            .clk(N__9980),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_15_4_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_15_4_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_15_4_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_7_LC_15_4_6  (
            .in0(_gnd_net_),
            .in1(N__10061),
            .in2(_gnd_net_),
            .in3(N__9893),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9980),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_15_4_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_15_4_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_15_4_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_15_4_7  (
            .in0(N__10504),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10122),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9980),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_15_5_0 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_15_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_15_5_0 .LUT_INIT=16'b0000001000010000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_1_LC_15_5_0  (
            .in0(N__10001),
            .in1(N__10148),
            .in2(N__10179),
            .in3(N__10538),
            .lcout(\U409_CIA.CLK_CIA_r_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_15_5_1 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_15_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_15_5_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_15_5_1  (
            .in0(N__10125),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9978),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_15_5_2 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_15_5_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_15_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_0_LC_15_5_2  (
            .in0(N__10045),
            .in1(N__10124),
            .in2(N__10514),
            .in3(N__10060),
            .lcout(),
            .ltout(\U409_CIA.CLK_CIA6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_LC_15_5_3 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_LC_15_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLK_CIA_LC_15_5_3 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \U409_CIA.CLK_CIA_LC_15_5_3  (
            .in0(N__10172),
            .in1(N__10202),
            .in2(N__10196),
            .in3(N__10086),
            .lcout(CLK_CIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9978),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_5_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_5_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_5_4  (
            .in0(N__10000),
            .in1(N__10147),
            .in2(N__10088),
            .in3(N__10123),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_2_0 ),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_15_5_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_15_5_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_15_5_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_15_5_5  (
            .in0(N__10478),
            .in1(N__10028),
            .in2(N__10097),
            .in3(N__10094),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9978),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_15_5_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_15_5_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_15_5_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_15_5_6  (
            .in0(_gnd_net_),
            .in1(N__10059),
            .in2(_gnd_net_),
            .in3(N__10044),
            .lcout(\U409_CIA.CLK_CIA6_4 ),
            .ltout(\U409_CIA.CLK_CIA6_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_15_5_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_15_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_15_5_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_15_5_7  (
            .in0(N__10016),
            .in1(N__10477),
            .in2(N__10010),
            .in3(N__10007),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9978),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_6_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_6_0  (
            .in0(_gnd_net_),
            .in1(N__9960),
            .in2(N__9947),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_6_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_15_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_15_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_15_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_15_6_1  (
            .in0(_gnd_net_),
            .in1(N__9922),
            .in2(_gnd_net_),
            .in3(N__9911),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__10569),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_15_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_15_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_15_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_15_6_2  (
            .in0(_gnd_net_),
            .in1(N__10381),
            .in2(_gnd_net_),
            .in3(N__10370),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__10569),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_15_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_15_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_15_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_15_6_3  (
            .in0(_gnd_net_),
            .in1(N__10363),
            .in2(_gnd_net_),
            .in3(N__10352),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__10569),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_15_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_15_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_15_6_4  (
            .in0(_gnd_net_),
            .in1(N__10348),
            .in2(_gnd_net_),
            .in3(N__10331),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_15_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_15_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_15_6_5  (
            .in0(_gnd_net_),
            .in1(N__10327),
            .in2(_gnd_net_),
            .in3(N__10301),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_15_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_15_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_15_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_15_6_6  (
            .in0(_gnd_net_),
            .in1(N__10297),
            .in2(_gnd_net_),
            .in3(N__10286),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__10569),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_15_6_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_15_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_15_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_15_6_7  (
            .in0(_gnd_net_),
            .in1(N__10282),
            .in2(_gnd_net_),
            .in3(N__10271),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__10569),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_15_7_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_15_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_15_7_0  (
            .in0(_gnd_net_),
            .in1(N__10264),
            .in2(_gnd_net_),
            .in3(N__10241),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_15_7_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_15_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_15_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_15_7_1  (
            .in0(_gnd_net_),
            .in1(N__10237),
            .in2(_gnd_net_),
            .in3(N__10226),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__10571),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_15_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_15_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(N__10219),
            .in2(_gnd_net_),
            .in3(N__10670),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_15_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_15_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_15_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_15_7_3  (
            .in0(_gnd_net_),
            .in1(N__10666),
            .in2(_gnd_net_),
            .in3(N__10655),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__10571),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_15_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_15_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_15_7_4  (
            .in0(_gnd_net_),
            .in1(N__10651),
            .in2(_gnd_net_),
            .in3(N__10634),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_15_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_15_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(N__10630),
            .in2(_gnd_net_),
            .in3(N__10613),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_15_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_15_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_15_7_6  (
            .in0(_gnd_net_),
            .in1(N__10609),
            .in2(_gnd_net_),
            .in3(N__10589),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_15_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_15_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_15_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_15_7_7  (
            .in0(_gnd_net_),
            .in1(N__10583),
            .in2(_gnd_net_),
            .in3(N__10586),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10571),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_16_5_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_16_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_16_5_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_16_5_4  (
            .in0(_gnd_net_),
            .in1(N__10536),
            .in2(_gnd_net_),
            .in3(N__10505),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_24_4_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_24_4_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_24_4_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_24_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_24_4_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_24_4_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_24_4_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_24_4_4  (
            .in0(N__10736),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10426),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS1n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNI692L_0_LC_24_4_5 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNI692L_0_LC_24_4_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNI692L_0_LC_24_4_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_CIA.VMA_RNI692L_0_LC_24_4_5  (
            .in0(N__10967),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10773),
            .lcout(CIA_ENABLE),
            .ltout(CIA_ENABLE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_24_4_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_24_4_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_24_4_6 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_24_4_6  (
            .in0(N__10723),
            .in1(_gnd_net_),
            .in2(N__10688),
            .in3(_gnd_net_),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS0n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Feb 2 2025 09:29:50

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    DMA_LATCH : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__11197\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \N_991_i\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_238_cascade_\ : std_logic;
signal \U712_REG_SM.N_238\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \U712_REG_SM.ASn_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.N_219_cascade_\ : std_logic;
signal \U712_REG_SM.N_304\ : std_logic;
signal \U712_REG_SM.N_304_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_0_i_0_1\ : std_logic;
signal \C3_c\ : std_logic;
signal \C1_c\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \U712_REG_SM.N_307\ : std_logic;
signal \U712_REG_SM.N_219\ : std_logic;
signal \U712_REG_SM.REG_TACK_RNOZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_235\ : std_logic;
signal \U712_CHIP_RAM.un5_DMA_CYCLE_START_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_225\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_1_1_3_cascade_\ : std_logic;
signal \U712_REG_SM.N_259\ : std_logic;
signal \U712_REG_SM.N_259_cascade_\ : std_logic;
signal \U712_REG_SM.N_236\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_i_0_0_3\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \N_40_i\ : std_logic;
signal \U712_REG_SM.N_261\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \N_41_i\ : std_logic;
signal \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_0\ : std_logic;
signal \U712_REG_SM.DS_EN_RNOZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_314\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_2\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \bfn_7_9_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.N_282_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_265_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_i_2_cascade_\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_218\ : std_logic;
signal \U712_CHIP_RAM.N_208_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_245_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a3_0_2\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \U712_BYTE_ENABLE.N_327\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \U712_BYTE_ENABLE.N_319_cascade_\ : std_logic;
signal \N_43_i\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_321\ : std_logic;
signal \A_c_1\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLMBEn_i_0Z0Z_0\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.N_233_i_0_en_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_233_i_0_en_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.N_209_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_359_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_290_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_181_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_a4_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.N_216_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.N_181\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_204_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_279_1\ : std_logic;
signal \U712_CHIP_RAM.N_279_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_398\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_393\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_227_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_226\ : std_logic;
signal \U712_CHIP_RAM.N_245\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_319\ : std_logic;
signal \U712_BYTE_ENABLE.N_322\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_cascade_\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \N_42_i\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_15\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_257\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_205\ : std_logic;
signal \U712_CHIP_RAM.N_205_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_216\ : std_logic;
signal \U712_CHIP_RAM.N_291\ : std_logic;
signal \U712_CHIP_RAM.N_291_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_204\ : std_logic;
signal \U712_CHIP_RAM.N_342_cascade_\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.N_352_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_395\ : std_logic;
signal \U712_CHIP_RAM.N_352\ : std_logic;
signal \U712_CHIP_RAM.N_293_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_99_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_290\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_359\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0\ : std_logic;
signal \U712_CHIP_RAM.N_301\ : std_logic;
signal \U712_CHIP_RAM.N_243\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_209\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_227\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_2\ : std_logic;
signal \U712_CHIP_RAM.N_303\ : std_logic;
signal \U712_CHIP_RAM.N_241\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \N_256\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_289\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_342\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_208\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_a3_0\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_10\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_14\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \un1_LDSn_i_0_0\ : std_logic;
signal \DS_ENm\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \un1_UDSn_i_0_0\ : std_logic;
signal \RASn_c\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10_cascade_\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \DMA_LATCH_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    \RESETn_wire\ <= RESETn;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    DMA_LATCH <= \DMA_LATCH_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__3777\,
            RESETB => \N__6582\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11197\,
            DIN => \N__11196\,
            DOUT => \N__11195\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11197\,
            PADOUT => \N__11196\,
            PADIN => \N__11195\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5469\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11188\,
            DIN => \N__11187\,
            DOUT => \N__11186\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11188\,
            PADOUT => \N__11187\,
            PADIN => \N__11186\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11179\,
            DIN => \N__11178\,
            DOUT => \N__11177\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11179\,
            PADOUT => \N__11178\,
            PADIN => \N__11177\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8322\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11170\,
            DIN => \N__11169\,
            DOUT => \N__11168\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11170\,
            PADOUT => \N__11169\,
            PADIN => \N__11168\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6609\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11161\,
            DIN => \N__11160\,
            DOUT => \N__11159\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11161\,
            PADOUT => \N__11160\,
            PADIN => \N__11159\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11152\,
            DIN => \N__11151\,
            DOUT => \N__11150\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11152\,
            PADOUT => \N__11151\,
            PADIN => \N__11150\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11143\,
            DIN => \N__11142\,
            DOUT => \N__11141\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11143\,
            PADOUT => \N__11142\,
            PADIN => \N__11141\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11134\,
            DIN => \N__11133\,
            DOUT => \N__11132\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11134\,
            PADOUT => \N__11133\,
            PADIN => \N__11132\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11125\,
            DIN => \N__11124\,
            DOUT => \N__11123\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11125\,
            PADOUT => \N__11124\,
            PADIN => \N__11123\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11116\,
            DIN => \N__11115\,
            DOUT => \N__11114\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11116\,
            PADOUT => \N__11115\,
            PADIN => \N__11114\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11107\,
            DIN => \N__11106\,
            DOUT => \N__11105\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11107\,
            PADOUT => \N__11106\,
            PADIN => \N__11105\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11098\,
            DIN => \N__11097\,
            DOUT => \N__11096\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11098\,
            PADOUT => \N__11097\,
            PADIN => \N__11096\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7620\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11089\,
            DIN => \N__11088\,
            DOUT => \N__11087\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11089\,
            PADOUT => \N__11088\,
            PADIN => \N__11087\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11080\,
            DIN => \N__11079\,
            DOUT => \N__11078\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11080\,
            PADOUT => \N__11079\,
            PADIN => \N__11078\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11071\,
            DIN => \N__11070\,
            DOUT => \N__11069\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11071\,
            PADOUT => \N__11070\,
            PADIN => \N__11069\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11062\,
            DIN => \N__11061\,
            DOUT => \N__11060\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11062\,
            PADOUT => \N__11061\,
            PADIN => \N__11060\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5001\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11053\,
            DIN => \N__11052\,
            DOUT => \N__11051\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11053\,
            PADOUT => \N__11052\,
            PADIN => \N__11051\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11044\,
            DIN => \N__11043\,
            DOUT => \N__11042\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11044\,
            PADOUT => \N__11043\,
            PADIN => \N__11042\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11035\,
            DIN => \N__11034\,
            DOUT => \N__11033\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11035\,
            PADOUT => \N__11034\,
            PADIN => \N__11033\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7353\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11026\,
            DIN => \N__11025\,
            DOUT => \N__11024\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11026\,
            PADOUT => \N__11025\,
            PADIN => \N__11024\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11017\,
            DIN => \N__11016\,
            DOUT => \N__11015\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11017\,
            PADOUT => \N__11016\,
            PADIN => \N__11015\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8355\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11008\,
            DIN => \N__11007\,
            DOUT => \N__11006\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11008\,
            PADOUT => \N__11007\,
            PADIN => \N__11006\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10999\,
            DIN => \N__10998\,
            DOUT => \N__10997\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10999\,
            PADOUT => \N__10998\,
            PADIN => \N__10997\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10990\,
            DIN => \N__10989\,
            DOUT => \N__10988\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10990\,
            PADOUT => \N__10989\,
            PADIN => \N__10988\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10981\,
            DIN => \N__10980\,
            DOUT => \N__10979\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10981\,
            PADOUT => \N__10980\,
            PADIN => \N__10979\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10972\,
            DIN => \N__10971\,
            DOUT => \N__10970\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10972\,
            PADOUT => \N__10971\,
            PADIN => \N__10970\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10963\,
            DIN => \N__10962\,
            DOUT => \N__10961\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10963\,
            PADOUT => \N__10962\,
            PADIN => \N__10961\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10954\,
            DIN => \N__10953\,
            DOUT => \N__10952\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10954\,
            PADOUT => \N__10953\,
            PADIN => \N__10952\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10945\,
            DIN => \N__10944\,
            DOUT => \N__10943\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10945\,
            PADOUT => \N__10944\,
            PADIN => \N__10943\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10936\,
            DIN => \N__10935\,
            DOUT => \N__10934\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10936\,
            PADOUT => \N__10935\,
            PADIN => \N__10934\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7368\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10927\,
            DIN => \N__10926\,
            DOUT => \N__10925\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10927\,
            PADOUT => \N__10926\,
            PADIN => \N__10925\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10918\,
            DIN => \N__10917\,
            DOUT => \N__10916\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10918\,
            PADOUT => \N__10917\,
            PADIN => \N__10916\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10909\,
            DIN => \N__10908\,
            DOUT => \N__10907\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10909\,
            PADOUT => \N__10908\,
            PADIN => \N__10907\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10900\,
            DIN => \N__10899\,
            DOUT => \N__10898\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10900\,
            PADOUT => \N__10899\,
            PADIN => \N__10898\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10891\,
            DIN => \N__10890\,
            DOUT => \N__10889\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10891\,
            PADOUT => \N__10890\,
            PADIN => \N__10889\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10882\,
            DIN => \N__10881\,
            DOUT => \N__10880\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10882\,
            PADOUT => \N__10881\,
            PADIN => \N__10880\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8508\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10873\,
            DIN => \N__10872\,
            DOUT => \N__10871\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10873\,
            PADOUT => \N__10872\,
            PADIN => \N__10871\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8766\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10864\,
            DIN => \N__10863\,
            DOUT => \N__10862\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10864\,
            PADOUT => \N__10863\,
            PADIN => \N__10862\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10855\,
            DIN => \N__10854\,
            DOUT => \N__10853\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10855\,
            PADOUT => \N__10854\,
            PADIN => \N__10853\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8376\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10846\,
            DIN => \N__10845\,
            DOUT => \N__10844\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10846\,
            PADOUT => \N__10845\,
            PADIN => \N__10844\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10837\,
            DIN => \N__10836\,
            DOUT => \N__10835\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10837\,
            PADOUT => \N__10836\,
            PADIN => \N__10835\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5910\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10828\,
            DIN => \N__10827\,
            DOUT => \N__10826\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10828\,
            PADOUT => \N__10827\,
            PADIN => \N__10826\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8762\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10819\,
            DIN => \N__10818\,
            DOUT => \N__10817\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10819\,
            PADOUT => \N__10818\,
            PADIN => \N__10817\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3867\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10810\,
            DIN => \N__10809\,
            DOUT => \N__10808\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10810\,
            PADOUT => \N__10809\,
            PADIN => \N__10808\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10801\,
            DIN => \N__10800\,
            DOUT => \N__10799\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10801\,
            PADOUT => \N__10800\,
            PADIN => \N__10799\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3849\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10792\,
            DIN => \N__10791\,
            DOUT => \N__10790\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10792\,
            PADOUT => \N__10791\,
            PADIN => \N__10790\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9120\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10783\,
            DIN => \N__10782\,
            DOUT => \N__10781\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10783\,
            PADOUT => \N__10782\,
            PADIN => \N__10781\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10774\,
            DIN => \N__10773\,
            DOUT => \N__10772\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10774\,
            PADOUT => \N__10773\,
            PADIN => \N__10772\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10765\,
            DIN => \N__10764\,
            DOUT => \N__10763\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10765\,
            PADOUT => \N__10764\,
            PADIN => \N__10763\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__10756\,
            DIN => \N__10755\,
            DOUT => \N__10754\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10756\,
            PADOUT => \N__10755\,
            PADIN => \N__10754\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10747\,
            DIN => \N__10746\,
            DOUT => \N__10745\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10747\,
            PADOUT => \N__10746\,
            PADIN => \N__10745\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8001\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10738\,
            DIN => \N__10737\,
            DOUT => \N__10736\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10738\,
            PADOUT => \N__10737\,
            PADIN => \N__10736\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10729\,
            DIN => \N__10728\,
            DOUT => \N__10727\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10729\,
            PADOUT => \N__10728\,
            PADIN => \N__10727\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8761\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10720\,
            DIN => \N__10719\,
            DOUT => \N__10718\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10720\,
            PADOUT => \N__10719\,
            PADIN => \N__10718\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6507\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10711\,
            DIN => \N__10710\,
            DOUT => \N__10709\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10711\,
            PADOUT => \N__10710\,
            PADIN => \N__10709\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5277\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10702\,
            DIN => \N__10701\,
            DOUT => \N__10700\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10702\,
            PADOUT => \N__10701\,
            PADIN => \N__10700\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4338\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10693\,
            DIN => \N__10692\,
            DOUT => \N__10691\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10693\,
            PADOUT => \N__10692\,
            PADIN => \N__10691\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6537\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10684\,
            DIN => \N__10683\,
            DOUT => \N__10682\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10684\,
            PADOUT => \N__10683\,
            PADIN => \N__10682\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4098\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10675\,
            DIN => \N__10674\,
            DOUT => \N__10673\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10675\,
            PADOUT => \N__10674\,
            PADIN => \N__10673\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10666\,
            DIN => \N__10665\,
            DOUT => \N__10664\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10666\,
            PADOUT => \N__10665\,
            PADIN => \N__10664\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10657\,
            DIN => \N__10656\,
            DOUT => \N__10655\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10657\,
            PADOUT => \N__10656\,
            PADIN => \N__10655\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4221\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10648\,
            DIN => \N__10647\,
            DOUT => \N__10646\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10648\,
            PADOUT => \N__10647\,
            PADIN => \N__10646\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8337\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10639\,
            DIN => \N__10638\,
            DOUT => \N__10637\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10639\,
            PADOUT => \N__10638\,
            PADIN => \N__10637\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5652\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10630\,
            DIN => \N__10629\,
            DOUT => \N__10628\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10630\,
            PADOUT => \N__10629\,
            PADIN => \N__10628\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5337\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10621\,
            DIN => \N__10620\,
            DOUT => \N__10619\,
            PACKAGEPIN => \DMA_LATCH_wire\
        );

    \DMA_LATCH_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10621\,
            PADOUT => \N__10620\,
            PADIN => \N__10619\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10612\,
            DIN => \N__10611\,
            DOUT => \N__10610\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10612\,
            PADOUT => \N__10611\,
            PADIN => \N__10610\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10603\,
            DIN => \N__10602\,
            DOUT => \N__10601\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10603\,
            PADOUT => \N__10602\,
            PADIN => \N__10601\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10594\,
            DIN => \N__10593\,
            DOUT => \N__10592\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10594\,
            PADOUT => \N__10593\,
            PADIN => \N__10592\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10585\,
            DIN => \N__10584\,
            DOUT => \N__10583\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10585\,
            PADOUT => \N__10584\,
            PADIN => \N__10583\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10576\,
            DIN => \N__10575\,
            DOUT => \N__10574\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10576\,
            PADOUT => \N__10575\,
            PADIN => \N__10574\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6492\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10567\,
            DIN => \N__10566\,
            DOUT => \N__10565\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10567\,
            PADOUT => \N__10566\,
            PADIN => \N__10565\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10558\,
            DIN => \N__10557\,
            DOUT => \N__10556\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10558\,
            PADOUT => \N__10557\,
            PADIN => \N__10556\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4929\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10549\,
            DIN => \N__10548\,
            DOUT => \N__10547\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__10549\,
            PADOUT => \N__10548\,
            PADIN => \N__10547\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3885\,
            DIN0 => OPEN,
            DOUT0 => \N__4536\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10540\,
            DIN => \N__10539\,
            DOUT => \N__10538\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10540\,
            PADOUT => \N__10539\,
            PADIN => \N__10538\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7632\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10531\,
            DIN => \N__10530\,
            DOUT => \N__10529\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10531\,
            PADOUT => \N__10530\,
            PADIN => \N__10529\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10522\,
            DIN => \N__10521\,
            DOUT => \N__10520\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10522\,
            PADOUT => \N__10521\,
            PADIN => \N__10520\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10513\,
            DIN => \N__10512\,
            DOUT => \N__10511\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10513\,
            PADOUT => \N__10512\,
            PADIN => \N__10511\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7398\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10504\,
            DIN => \N__10503\,
            DOUT => \N__10502\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10504\,
            PADOUT => \N__10503\,
            PADIN => \N__10502\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10495\,
            DIN => \N__10494\,
            DOUT => \N__10493\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10495\,
            PADOUT => \N__10494\,
            PADIN => \N__10493\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10486\,
            DIN => \N__10485\,
            DOUT => \N__10484\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10486\,
            PADOUT => \N__10485\,
            PADIN => \N__10484\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10477\,
            DIN => \N__10476\,
            DOUT => \N__10475\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10477\,
            PADOUT => \N__10476\,
            PADIN => \N__10475\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10468\,
            DIN => \N__10467\,
            DOUT => \N__10466\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10468\,
            PADOUT => \N__10467\,
            PADIN => \N__10466\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7593\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10459\,
            DIN => \N__10458\,
            DOUT => \N__10457\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10459\,
            PADOUT => \N__10458\,
            PADIN => \N__10457\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8391\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10450\,
            DIN => \N__10449\,
            DOUT => \N__10448\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10450\,
            PADOUT => \N__10449\,
            PADIN => \N__10448\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5217\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10441\,
            DIN => \N__10440\,
            DOUT => \N__10439\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10441\,
            PADOUT => \N__10440\,
            PADIN => \N__10439\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10432\,
            DIN => \N__10431\,
            DOUT => \N__10430\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10432\,
            PADOUT => \N__10431\,
            PADIN => \N__10430\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2541\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10408\
        );

    \I__2540\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10405\
        );

    \I__2539\ : InMux
    port map (
            O => \N__10411\,
            I => \N__10401\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__10408\,
            I => \N__10398\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__10405\,
            I => \N__10395\
        );

    \I__2536\ : InMux
    port map (
            O => \N__10404\,
            I => \N__10392\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__10401\,
            I => \N__10389\
        );

    \I__2534\ : Span4Mux_v
    port map (
            O => \N__10398\,
            I => \N__10382\
        );

    \I__2533\ : Span4Mux_h
    port map (
            O => \N__10395\,
            I => \N__10382\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__10392\,
            I => \N__10382\
        );

    \I__2531\ : Sp12to4
    port map (
            O => \N__10389\,
            I => \N__10379\
        );

    \I__2530\ : Span4Mux_h
    port map (
            O => \N__10382\,
            I => \N__10376\
        );

    \I__2529\ : Span12Mux_v
    port map (
            O => \N__10379\,
            I => \N__10373\
        );

    \I__2528\ : Span4Mux_v
    port map (
            O => \N__10376\,
            I => \N__10370\
        );

    \I__2527\ : Span12Mux_h
    port map (
            O => \N__10373\,
            I => \N__10367\
        );

    \I__2526\ : Sp12to4
    port map (
            O => \N__10370\,
            I => \N__10364\
        );

    \I__2525\ : Odrv12
    port map (
            O => \N__10367\,
            I => \DRA_c_6\
        );

    \I__2524\ : Odrv12
    port map (
            O => \N__10364\,
            I => \DRA_c_6\
        );

    \I__2523\ : InMux
    port map (
            O => \N__10359\,
            I => \N__10354\
        );

    \I__2522\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10348\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__10357\,
            I => \N__10343\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__10354\,
            I => \N__10335\
        );

    \I__2519\ : InMux
    port map (
            O => \N__10353\,
            I => \N__10332\
        );

    \I__2518\ : InMux
    port map (
            O => \N__10352\,
            I => \N__10329\
        );

    \I__2517\ : InMux
    port map (
            O => \N__10351\,
            I => \N__10326\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__10348\,
            I => \N__10323\
        );

    \I__2515\ : InMux
    port map (
            O => \N__10347\,
            I => \N__10320\
        );

    \I__2514\ : InMux
    port map (
            O => \N__10346\,
            I => \N__10317\
        );

    \I__2513\ : InMux
    port map (
            O => \N__10343\,
            I => \N__10308\
        );

    \I__2512\ : InMux
    port map (
            O => \N__10342\,
            I => \N__10308\
        );

    \I__2511\ : InMux
    port map (
            O => \N__10341\,
            I => \N__10308\
        );

    \I__2510\ : InMux
    port map (
            O => \N__10340\,
            I => \N__10308\
        );

    \I__2509\ : InMux
    port map (
            O => \N__10339\,
            I => \N__10305\
        );

    \I__2508\ : InMux
    port map (
            O => \N__10338\,
            I => \N__10300\
        );

    \I__2507\ : Span4Mux_h
    port map (
            O => \N__10335\,
            I => \N__10285\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__10332\,
            I => \N__10285\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__10329\,
            I => \N__10285\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__10326\,
            I => \N__10285\
        );

    \I__2503\ : Span4Mux_v
    port map (
            O => \N__10323\,
            I => \N__10282\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__10320\,
            I => \N__10273\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__10317\,
            I => \N__10273\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__10308\,
            I => \N__10273\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__10305\,
            I => \N__10273\
        );

    \I__2498\ : InMux
    port map (
            O => \N__10304\,
            I => \N__10268\
        );

    \I__2497\ : InMux
    port map (
            O => \N__10303\,
            I => \N__10268\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__10300\,
            I => \N__10265\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10299\,
            I => \N__10260\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10298\,
            I => \N__10260\
        );

    \I__2493\ : InMux
    port map (
            O => \N__10297\,
            I => \N__10257\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10296\,
            I => \N__10252\
        );

    \I__2491\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10252\
        );

    \I__2490\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10249\
        );

    \I__2489\ : Span4Mux_v
    port map (
            O => \N__10285\,
            I => \N__10246\
        );

    \I__2488\ : Span4Mux_h
    port map (
            O => \N__10282\,
            I => \N__10239\
        );

    \I__2487\ : Span4Mux_v
    port map (
            O => \N__10273\,
            I => \N__10239\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__10268\,
            I => \N__10239\
        );

    \I__2485\ : Sp12to4
    port map (
            O => \N__10265\,
            I => \N__10232\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__10260\,
            I => \N__10232\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__10257\,
            I => \N__10232\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__10252\,
            I => \N__10227\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__10249\,
            I => \N__10227\
        );

    \I__2480\ : Sp12to4
    port map (
            O => \N__10246\,
            I => \N__10222\
        );

    \I__2479\ : Sp12to4
    port map (
            O => \N__10239\,
            I => \N__10222\
        );

    \I__2478\ : Span12Mux_h
    port map (
            O => \N__10232\,
            I => \N__10219\
        );

    \I__2477\ : Span12Mux_v
    port map (
            O => \N__10227\,
            I => \N__10216\
        );

    \I__2476\ : Span12Mux_h
    port map (
            O => \N__10222\,
            I => \N__10213\
        );

    \I__2475\ : Span12Mux_v
    port map (
            O => \N__10219\,
            I => \N__10208\
        );

    \I__2474\ : Span12Mux_h
    port map (
            O => \N__10216\,
            I => \N__10208\
        );

    \I__2473\ : Span12Mux_v
    port map (
            O => \N__10213\,
            I => \N__10205\
        );

    \I__2472\ : Odrv12
    port map (
            O => \N__10208\,
            I => \AGNUS_REV_c\
        );

    \I__2471\ : Odrv12
    port map (
            O => \N__10205\,
            I => \AGNUS_REV_c\
        );

    \I__2470\ : InMux
    port map (
            O => \N__10200\,
            I => \N__10195\
        );

    \I__2469\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10192\
        );

    \I__2468\ : InMux
    port map (
            O => \N__10198\,
            I => \N__10189\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__10195\,
            I => \N__10183\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10192\,
            I => \N__10183\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__10189\,
            I => \N__10180\
        );

    \I__2464\ : InMux
    port map (
            O => \N__10188\,
            I => \N__10177\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__10183\,
            I => \N__10174\
        );

    \I__2462\ : Span4Mux_v
    port map (
            O => \N__10180\,
            I => \N__10169\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__10177\,
            I => \N__10169\
        );

    \I__2460\ : Span4Mux_v
    port map (
            O => \N__10174\,
            I => \N__10166\
        );

    \I__2459\ : Span4Mux_v
    port map (
            O => \N__10169\,
            I => \N__10163\
        );

    \I__2458\ : Sp12to4
    port map (
            O => \N__10166\,
            I => \N__10158\
        );

    \I__2457\ : Sp12to4
    port map (
            O => \N__10163\,
            I => \N__10158\
        );

    \I__2456\ : Span12Mux_h
    port map (
            O => \N__10158\,
            I => \N__10155\
        );

    \I__2455\ : Odrv12
    port map (
            O => \N__10155\,
            I => \DRA_c_5\
        );

    \I__2454\ : InMux
    port map (
            O => \N__10152\,
            I => \N__10146\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10151\,
            I => \N__10146\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__10146\,
            I => \N__10143\
        );

    \I__2451\ : Odrv12
    port map (
            O => \N__10143\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2450\ : InMux
    port map (
            O => \N__10140\,
            I => \N__10137\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__10137\,
            I => \N__10125\
        );

    \I__2448\ : ClkMux
    port map (
            O => \N__10136\,
            I => \N__10104\
        );

    \I__2447\ : ClkMux
    port map (
            O => \N__10135\,
            I => \N__10104\
        );

    \I__2446\ : ClkMux
    port map (
            O => \N__10134\,
            I => \N__10104\
        );

    \I__2445\ : ClkMux
    port map (
            O => \N__10133\,
            I => \N__10104\
        );

    \I__2444\ : ClkMux
    port map (
            O => \N__10132\,
            I => \N__10104\
        );

    \I__2443\ : ClkMux
    port map (
            O => \N__10131\,
            I => \N__10104\
        );

    \I__2442\ : ClkMux
    port map (
            O => \N__10130\,
            I => \N__10104\
        );

    \I__2441\ : ClkMux
    port map (
            O => \N__10129\,
            I => \N__10104\
        );

    \I__2440\ : ClkMux
    port map (
            O => \N__10128\,
            I => \N__10104\
        );

    \I__2439\ : Glb2LocalMux
    port map (
            O => \N__10125\,
            I => \N__10104\
        );

    \I__2438\ : GlobalMux
    port map (
            O => \N__10104\,
            I => \N__10101\
        );

    \I__2437\ : gio2CtrlBuf
    port map (
            O => \N__10101\,
            I => \C3_c_g\
        );

    \I__2436\ : CEMux
    port map (
            O => \N__10098\,
            I => \N__10094\
        );

    \I__2435\ : CEMux
    port map (
            O => \N__10097\,
            I => \N__10087\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__10094\,
            I => \N__10083\
        );

    \I__2433\ : CEMux
    port map (
            O => \N__10093\,
            I => \N__10080\
        );

    \I__2432\ : CEMux
    port map (
            O => \N__10092\,
            I => \N__10077\
        );

    \I__2431\ : CEMux
    port map (
            O => \N__10091\,
            I => \N__10074\
        );

    \I__2430\ : CEMux
    port map (
            O => \N__10090\,
            I => \N__10071\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__10087\,
            I => \N__10068\
        );

    \I__2428\ : CEMux
    port map (
            O => \N__10086\,
            I => \N__10065\
        );

    \I__2427\ : Span4Mux_v
    port map (
            O => \N__10083\,
            I => \N__10059\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__10080\,
            I => \N__10059\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__10077\,
            I => \N__10056\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__10074\,
            I => \N__10053\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__10071\,
            I => \N__10046\
        );

    \I__2422\ : Span4Mux_v
    port map (
            O => \N__10068\,
            I => \N__10046\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__10065\,
            I => \N__10046\
        );

    \I__2420\ : CEMux
    port map (
            O => \N__10064\,
            I => \N__10043\
        );

    \I__2419\ : Span4Mux_h
    port map (
            O => \N__10059\,
            I => \N__10038\
        );

    \I__2418\ : Span4Mux_h
    port map (
            O => \N__10056\,
            I => \N__10038\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__10053\,
            I => \N__10035\
        );

    \I__2416\ : Span4Mux_h
    port map (
            O => \N__10046\,
            I => \N__10032\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__10043\,
            I => \N__10029\
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__10038\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\
        );

    \I__2413\ : Odrv4
    port map (
            O => \N__10035\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\
        );

    \I__2412\ : Odrv4
    port map (
            O => \N__10032\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\
        );

    \I__2411\ : Odrv12
    port map (
            O => \N__10029\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10012\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10019\,
            I => \N__10009\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10018\,
            I => \N__10006\
        );

    \I__2407\ : InMux
    port map (
            O => \N__10017\,
            I => \N__10003\
        );

    \I__2406\ : InMux
    port map (
            O => \N__10016\,
            I => \N__9998\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10015\,
            I => \N__9998\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10012\,
            I => \N__9991\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__10009\,
            I => \N__9983\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__10006\,
            I => \N__9975\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__10003\,
            I => \N__9965\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__9998\,
            I => \N__9943\
        );

    \I__2399\ : SRMux
    port map (
            O => \N__9997\,
            I => \N__9852\
        );

    \I__2398\ : SRMux
    port map (
            O => \N__9996\,
            I => \N__9852\
        );

    \I__2397\ : SRMux
    port map (
            O => \N__9995\,
            I => \N__9852\
        );

    \I__2396\ : SRMux
    port map (
            O => \N__9994\,
            I => \N__9852\
        );

    \I__2395\ : Glb2LocalMux
    port map (
            O => \N__9991\,
            I => \N__9852\
        );

    \I__2394\ : SRMux
    port map (
            O => \N__9990\,
            I => \N__9852\
        );

    \I__2393\ : SRMux
    port map (
            O => \N__9989\,
            I => \N__9852\
        );

    \I__2392\ : SRMux
    port map (
            O => \N__9988\,
            I => \N__9852\
        );

    \I__2391\ : SRMux
    port map (
            O => \N__9987\,
            I => \N__9852\
        );

    \I__2390\ : SRMux
    port map (
            O => \N__9986\,
            I => \N__9852\
        );

    \I__2389\ : Glb2LocalMux
    port map (
            O => \N__9983\,
            I => \N__9852\
        );

    \I__2388\ : SRMux
    port map (
            O => \N__9982\,
            I => \N__9852\
        );

    \I__2387\ : SRMux
    port map (
            O => \N__9981\,
            I => \N__9852\
        );

    \I__2386\ : SRMux
    port map (
            O => \N__9980\,
            I => \N__9852\
        );

    \I__2385\ : SRMux
    port map (
            O => \N__9979\,
            I => \N__9852\
        );

    \I__2384\ : SRMux
    port map (
            O => \N__9978\,
            I => \N__9852\
        );

    \I__2383\ : Glb2LocalMux
    port map (
            O => \N__9975\,
            I => \N__9852\
        );

    \I__2382\ : SRMux
    port map (
            O => \N__9974\,
            I => \N__9852\
        );

    \I__2381\ : SRMux
    port map (
            O => \N__9973\,
            I => \N__9852\
        );

    \I__2380\ : SRMux
    port map (
            O => \N__9972\,
            I => \N__9852\
        );

    \I__2379\ : SRMux
    port map (
            O => \N__9971\,
            I => \N__9852\
        );

    \I__2378\ : SRMux
    port map (
            O => \N__9970\,
            I => \N__9852\
        );

    \I__2377\ : SRMux
    port map (
            O => \N__9969\,
            I => \N__9852\
        );

    \I__2376\ : SRMux
    port map (
            O => \N__9968\,
            I => \N__9852\
        );

    \I__2375\ : Glb2LocalMux
    port map (
            O => \N__9965\,
            I => \N__9852\
        );

    \I__2374\ : SRMux
    port map (
            O => \N__9964\,
            I => \N__9852\
        );

    \I__2373\ : SRMux
    port map (
            O => \N__9963\,
            I => \N__9852\
        );

    \I__2372\ : SRMux
    port map (
            O => \N__9962\,
            I => \N__9852\
        );

    \I__2371\ : SRMux
    port map (
            O => \N__9961\,
            I => \N__9852\
        );

    \I__2370\ : SRMux
    port map (
            O => \N__9960\,
            I => \N__9852\
        );

    \I__2369\ : SRMux
    port map (
            O => \N__9959\,
            I => \N__9852\
        );

    \I__2368\ : SRMux
    port map (
            O => \N__9958\,
            I => \N__9852\
        );

    \I__2367\ : SRMux
    port map (
            O => \N__9957\,
            I => \N__9852\
        );

    \I__2366\ : SRMux
    port map (
            O => \N__9956\,
            I => \N__9852\
        );

    \I__2365\ : SRMux
    port map (
            O => \N__9955\,
            I => \N__9852\
        );

    \I__2364\ : SRMux
    port map (
            O => \N__9954\,
            I => \N__9852\
        );

    \I__2363\ : SRMux
    port map (
            O => \N__9953\,
            I => \N__9852\
        );

    \I__2362\ : SRMux
    port map (
            O => \N__9952\,
            I => \N__9852\
        );

    \I__2361\ : SRMux
    port map (
            O => \N__9951\,
            I => \N__9852\
        );

    \I__2360\ : SRMux
    port map (
            O => \N__9950\,
            I => \N__9852\
        );

    \I__2359\ : SRMux
    port map (
            O => \N__9949\,
            I => \N__9852\
        );

    \I__2358\ : SRMux
    port map (
            O => \N__9948\,
            I => \N__9852\
        );

    \I__2357\ : SRMux
    port map (
            O => \N__9947\,
            I => \N__9852\
        );

    \I__2356\ : SRMux
    port map (
            O => \N__9946\,
            I => \N__9852\
        );

    \I__2355\ : Glb2LocalMux
    port map (
            O => \N__9943\,
            I => \N__9852\
        );

    \I__2354\ : GlobalMux
    port map (
            O => \N__9852\,
            I => \N__9849\
        );

    \I__2353\ : gio2CtrlBuf
    port map (
            O => \N__9849\,
            I => \RESETn_c_i_g\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__9846\,
            I => \N__9843\
        );

    \I__2351\ : InMux
    port map (
            O => \N__9843\,
            I => \N__9840\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__9840\,
            I => \N__9837\
        );

    \I__2349\ : Span4Mux_h
    port map (
            O => \N__9837\,
            I => \N__9834\
        );

    \I__2348\ : Odrv4
    port map (
            O => \N__9834\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2347\ : InMux
    port map (
            O => \N__9831\,
            I => \N__9823\
        );

    \I__2346\ : InMux
    port map (
            O => \N__9830\,
            I => \N__9823\
        );

    \I__2345\ : InMux
    port map (
            O => \N__9829\,
            I => \N__9820\
        );

    \I__2344\ : InMux
    port map (
            O => \N__9828\,
            I => \N__9817\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__9823\,
            I => \N__9814\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__9820\,
            I => \N__9809\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__9817\,
            I => \N__9809\
        );

    \I__2340\ : Span4Mux_v
    port map (
            O => \N__9814\,
            I => \N__9806\
        );

    \I__2339\ : Span4Mux_v
    port map (
            O => \N__9809\,
            I => \N__9803\
        );

    \I__2338\ : Span4Mux_h
    port map (
            O => \N__9806\,
            I => \N__9800\
        );

    \I__2337\ : Sp12to4
    port map (
            O => \N__9803\,
            I => \N__9797\
        );

    \I__2336\ : Sp12to4
    port map (
            O => \N__9800\,
            I => \N__9792\
        );

    \I__2335\ : Span12Mux_h
    port map (
            O => \N__9797\,
            I => \N__9792\
        );

    \I__2334\ : Odrv12
    port map (
            O => \N__9792\,
            I => \DRA_c_7\
        );

    \I__2333\ : InMux
    port map (
            O => \N__9789\,
            I => \N__9786\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__9786\,
            I => \N__9783\
        );

    \I__2331\ : Span4Mux_h
    port map (
            O => \N__9783\,
            I => \N__9780\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__9780\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2329\ : InMux
    port map (
            O => \N__9777\,
            I => \N__9774\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__9774\,
            I => \N__9771\
        );

    \I__2327\ : Odrv4
    port map (
            O => \N__9771\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2326\ : InMux
    port map (
            O => \N__9768\,
            I => \N__9765\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__9765\,
            I => \N__9759\
        );

    \I__2324\ : InMux
    port map (
            O => \N__9764\,
            I => \N__9756\
        );

    \I__2323\ : InMux
    port map (
            O => \N__9763\,
            I => \N__9751\
        );

    \I__2322\ : InMux
    port map (
            O => \N__9762\,
            I => \N__9751\
        );

    \I__2321\ : Span4Mux_h
    port map (
            O => \N__9759\,
            I => \N__9746\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__9756\,
            I => \N__9746\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__9751\,
            I => \N__9741\
        );

    \I__2318\ : Sp12to4
    port map (
            O => \N__9746\,
            I => \N__9741\
        );

    \I__2317\ : Span12Mux_v
    port map (
            O => \N__9741\,
            I => \N__9738\
        );

    \I__2316\ : Span12Mux_h
    port map (
            O => \N__9738\,
            I => \N__9735\
        );

    \I__2315\ : Odrv12
    port map (
            O => \N__9735\,
            I => \DRA_c_3\
        );

    \I__2314\ : InMux
    port map (
            O => \N__9732\,
            I => \N__9729\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__9729\,
            I => \N__9726\
        );

    \I__2312\ : Odrv4
    port map (
            O => \N__9726\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2311\ : InMux
    port map (
            O => \N__9723\,
            I => \N__9717\
        );

    \I__2310\ : InMux
    port map (
            O => \N__9722\,
            I => \N__9714\
        );

    \I__2309\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9709\
        );

    \I__2308\ : InMux
    port map (
            O => \N__9720\,
            I => \N__9709\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__9717\,
            I => \N__9704\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__9714\,
            I => \N__9704\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__9709\,
            I => \N__9701\
        );

    \I__2304\ : Span4Mux_v
    port map (
            O => \N__9704\,
            I => \N__9698\
        );

    \I__2303\ : Span4Mux_h
    port map (
            O => \N__9701\,
            I => \N__9695\
        );

    \I__2302\ : Span4Mux_v
    port map (
            O => \N__9698\,
            I => \N__9692\
        );

    \I__2301\ : Span4Mux_v
    port map (
            O => \N__9695\,
            I => \N__9689\
        );

    \I__2300\ : Sp12to4
    port map (
            O => \N__9692\,
            I => \N__9684\
        );

    \I__2299\ : Sp12to4
    port map (
            O => \N__9689\,
            I => \N__9684\
        );

    \I__2298\ : Span12Mux_h
    port map (
            O => \N__9684\,
            I => \N__9681\
        );

    \I__2297\ : Odrv12
    port map (
            O => \N__9681\,
            I => \DRA_c_4\
        );

    \I__2296\ : InMux
    port map (
            O => \N__9678\,
            I => \N__9675\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__9675\,
            I => \N__9672\
        );

    \I__2294\ : Span4Mux_h
    port map (
            O => \N__9672\,
            I => \N__9669\
        );

    \I__2293\ : Odrv4
    port map (
            O => \N__9669\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__9666\,
            I => \N__9663\
        );

    \I__2291\ : InMux
    port map (
            O => \N__9663\,
            I => \N__9659\
        );

    \I__2290\ : InMux
    port map (
            O => \N__9662\,
            I => \N__9656\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__9659\,
            I => \N__9651\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__9656\,
            I => \N__9651\
        );

    \I__2287\ : Span12Mux_h
    port map (
            O => \N__9651\,
            I => \N__9648\
        );

    \I__2286\ : Span12Mux_v
    port map (
            O => \N__9648\,
            I => \N__9645\
        );

    \I__2285\ : Odrv12
    port map (
            O => \N__9645\,
            I => \DRA_c_0\
        );

    \I__2284\ : InMux
    port map (
            O => \N__9642\,
            I => \N__9639\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__9639\,
            I => \N__9636\
        );

    \I__2282\ : Span4Mux_h
    port map (
            O => \N__9636\,
            I => \N__9633\
        );

    \I__2281\ : Odrv4
    port map (
            O => \N__9633\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2280\ : InMux
    port map (
            O => \N__9630\,
            I => \N__9625\
        );

    \I__2279\ : InMux
    port map (
            O => \N__9629\,
            I => \N__9622\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__9628\,
            I => \N__9619\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__9625\,
            I => \N__9615\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__9622\,
            I => \N__9612\
        );

    \I__2275\ : InMux
    port map (
            O => \N__9619\,
            I => \N__9609\
        );

    \I__2274\ : InMux
    port map (
            O => \N__9618\,
            I => \N__9606\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__9615\,
            I => \N__9603\
        );

    \I__2272\ : Span4Mux_v
    port map (
            O => \N__9612\,
            I => \N__9596\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__9609\,
            I => \N__9596\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__9606\,
            I => \N__9596\
        );

    \I__2269\ : Span4Mux_v
    port map (
            O => \N__9603\,
            I => \N__9593\
        );

    \I__2268\ : Span4Mux_v
    port map (
            O => \N__9596\,
            I => \N__9590\
        );

    \I__2267\ : Sp12to4
    port map (
            O => \N__9593\,
            I => \N__9585\
        );

    \I__2266\ : Sp12to4
    port map (
            O => \N__9590\,
            I => \N__9585\
        );

    \I__2265\ : Span12Mux_h
    port map (
            O => \N__9585\,
            I => \N__9582\
        );

    \I__2264\ : Span12Mux_v
    port map (
            O => \N__9582\,
            I => \N__9579\
        );

    \I__2263\ : Odrv12
    port map (
            O => \N__9579\,
            I => \DRA_c_9\
        );

    \I__2262\ : InMux
    port map (
            O => \N__9576\,
            I => \N__9571\
        );

    \I__2261\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9568\
        );

    \I__2260\ : InMux
    port map (
            O => \N__9574\,
            I => \N__9565\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__9571\,
            I => \N__9562\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__9568\,
            I => \N__9557\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__9565\,
            I => \N__9557\
        );

    \I__2256\ : Span4Mux_v
    port map (
            O => \N__9562\,
            I => \N__9553\
        );

    \I__2255\ : Span4Mux_v
    port map (
            O => \N__9557\,
            I => \N__9550\
        );

    \I__2254\ : InMux
    port map (
            O => \N__9556\,
            I => \N__9547\
        );

    \I__2253\ : Span4Mux_h
    port map (
            O => \N__9553\,
            I => \N__9544\
        );

    \I__2252\ : Span4Mux_h
    port map (
            O => \N__9550\,
            I => \N__9541\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__9547\,
            I => \N__9538\
        );

    \I__2250\ : Sp12to4
    port map (
            O => \N__9544\,
            I => \N__9531\
        );

    \I__2249\ : Sp12to4
    port map (
            O => \N__9541\,
            I => \N__9531\
        );

    \I__2248\ : Span12Mux_h
    port map (
            O => \N__9538\,
            I => \N__9531\
        );

    \I__2247\ : Odrv12
    port map (
            O => \N__9531\,
            I => \DRA_c_8\
        );

    \I__2246\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__9525\,
            I => \N__9522\
        );

    \I__2244\ : Span12Mux_v
    port map (
            O => \N__9522\,
            I => \N__9519\
        );

    \I__2243\ : Odrv12
    port map (
            O => \N__9519\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9516\,
            I => \N__9509\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9515\,
            I => \N__9509\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9514\,
            I => \N__9505\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__9509\,
            I => \N__9502\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9508\,
            I => \N__9499\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__9505\,
            I => \N__9492\
        );

    \I__2236\ : Span4Mux_h
    port map (
            O => \N__9502\,
            I => \N__9492\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__9499\,
            I => \N__9492\
        );

    \I__2234\ : Span4Mux_v
    port map (
            O => \N__9492\,
            I => \N__9489\
        );

    \I__2233\ : Sp12to4
    port map (
            O => \N__9489\,
            I => \N__9486\
        );

    \I__2232\ : Span12Mux_h
    port map (
            O => \N__9486\,
            I => \N__9483\
        );

    \I__2231\ : Span12Mux_v
    port map (
            O => \N__9483\,
            I => \N__9480\
        );

    \I__2230\ : Odrv12
    port map (
            O => \N__9480\,
            I => \DRA_c_2\
        );

    \I__2229\ : InMux
    port map (
            O => \N__9477\,
            I => \N__9474\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__9474\,
            I => \N__9469\
        );

    \I__2227\ : InMux
    port map (
            O => \N__9473\,
            I => \N__9466\
        );

    \I__2226\ : InMux
    port map (
            O => \N__9472\,
            I => \N__9462\
        );

    \I__2225\ : Span4Mux_v
    port map (
            O => \N__9469\,
            I => \N__9459\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__9466\,
            I => \N__9456\
        );

    \I__2223\ : InMux
    port map (
            O => \N__9465\,
            I => \N__9453\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__9462\,
            I => \N__9450\
        );

    \I__2221\ : Sp12to4
    port map (
            O => \N__9459\,
            I => \N__9447\
        );

    \I__2220\ : Sp12to4
    port map (
            O => \N__9456\,
            I => \N__9442\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__9453\,
            I => \N__9442\
        );

    \I__2218\ : Span12Mux_h
    port map (
            O => \N__9450\,
            I => \N__9439\
        );

    \I__2217\ : Span12Mux_h
    port map (
            O => \N__9447\,
            I => \N__9436\
        );

    \I__2216\ : Span12Mux_v
    port map (
            O => \N__9442\,
            I => \N__9433\
        );

    \I__2215\ : Span12Mux_v
    port map (
            O => \N__9439\,
            I => \N__9430\
        );

    \I__2214\ : Span12Mux_v
    port map (
            O => \N__9436\,
            I => \N__9425\
        );

    \I__2213\ : Span12Mux_h
    port map (
            O => \N__9433\,
            I => \N__9425\
        );

    \I__2212\ : Odrv12
    port map (
            O => \N__9430\,
            I => \DRA_c_1\
        );

    \I__2211\ : Odrv12
    port map (
            O => \N__9425\,
            I => \DRA_c_1\
        );

    \I__2210\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9414\
        );

    \I__2209\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9414\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__9414\,
            I => \N__9411\
        );

    \I__2207\ : Odrv12
    port map (
            O => \N__9411\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2206\ : InMux
    port map (
            O => \N__9408\,
            I => \N__9405\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__9405\,
            I => \N__9402\
        );

    \I__2204\ : Span4Mux_h
    port map (
            O => \N__9402\,
            I => \N__9399\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__9399\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9396\,
            I => \N__9393\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__9393\,
            I => \N__9390\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__9390\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2199\ : InMux
    port map (
            O => \N__9387\,
            I => \N__9384\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__9384\,
            I => \N__9381\
        );

    \I__2197\ : Span4Mux_h
    port map (
            O => \N__9381\,
            I => \N__9378\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__9378\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9375\,
            I => \N__9372\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__9372\,
            I => \N__9369\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__9369\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9366\,
            I => \N__9363\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__9363\,
            I => \N__9360\
        );

    \I__2190\ : Odrv4
    port map (
            O => \N__9360\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2189\ : InMux
    port map (
            O => \N__9357\,
            I => \N__9354\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__9354\,
            I => \N__9351\
        );

    \I__2187\ : Span4Mux_h
    port map (
            O => \N__9351\,
            I => \N__9348\
        );

    \I__2186\ : Odrv4
    port map (
            O => \N__9348\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9345\,
            I => \N__9342\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__9342\,
            I => \N__9339\
        );

    \I__2183\ : Span4Mux_h
    port map (
            O => \N__9339\,
            I => \N__9336\
        );

    \I__2182\ : Span4Mux_h
    port map (
            O => \N__9336\,
            I => \N__9333\
        );

    \I__2181\ : Odrv4
    port map (
            O => \N__9333\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9330\,
            I => \N__9327\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9327\,
            I => \N__9324\
        );

    \I__2178\ : Span4Mux_h
    port map (
            O => \N__9324\,
            I => \N__9321\
        );

    \I__2177\ : Odrv4
    port map (
            O => \N__9321\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2176\ : InMux
    port map (
            O => \N__9318\,
            I => \N__9315\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__9315\,
            I => \N__9312\
        );

    \I__2174\ : Span4Mux_h
    port map (
            O => \N__9312\,
            I => \N__9309\
        );

    \I__2173\ : Odrv4
    port map (
            O => \N__9309\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2172\ : CEMux
    port map (
            O => \N__9306\,
            I => \N__9302\
        );

    \I__2171\ : CEMux
    port map (
            O => \N__9305\,
            I => \N__9299\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9302\,
            I => \N__9296\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__9299\,
            I => \N__9293\
        );

    \I__2168\ : Span4Mux_v
    port map (
            O => \N__9296\,
            I => \N__9287\
        );

    \I__2167\ : Span12Mux_h
    port map (
            O => \N__9293\,
            I => \N__9284\
        );

    \I__2166\ : CEMux
    port map (
            O => \N__9292\,
            I => \N__9281\
        );

    \I__2165\ : CEMux
    port map (
            O => \N__9291\,
            I => \N__9278\
        );

    \I__2164\ : CEMux
    port map (
            O => \N__9290\,
            I => \N__9275\
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__9287\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\
        );

    \I__2162\ : Odrv12
    port map (
            O => \N__9284\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__9281\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__9278\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__9275\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9264\,
            I => \N__9261\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9261\,
            I => \N__9257\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9254\
        );

    \I__2155\ : Span4Mux_v
    port map (
            O => \N__9257\,
            I => \N__9251\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9254\,
            I => \N__9248\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__9251\,
            I => \N__9243\
        );

    \I__2152\ : Span4Mux_v
    port map (
            O => \N__9248\,
            I => \N__9243\
        );

    \I__2151\ : Sp12to4
    port map (
            O => \N__9243\,
            I => \N__9240\
        );

    \I__2150\ : Span12Mux_h
    port map (
            O => \N__9240\,
            I => \N__9237\
        );

    \I__2149\ : Odrv12
    port map (
            O => \N__9237\,
            I => \RAS0n_c\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9231\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__9231\,
            I => \N__9228\
        );

    \I__2146\ : Span4Mux_h
    port map (
            O => \N__9228\,
            I => \N__9225\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__9225\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9214\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9211\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9206\
        );

    \I__2141\ : InMux
    port map (
            O => \N__9219\,
            I => \N__9206\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9218\,
            I => \N__9201\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9201\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9214\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9211\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9206\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__9201\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2134\ : CascadeMux
    port map (
            O => \N__9192\,
            I => \N__9185\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__9191\,
            I => \N__9182\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__9190\,
            I => \N__9179\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__9189\,
            I => \N__9174\
        );

    \I__2130\ : CascadeMux
    port map (
            O => \N__9188\,
            I => \N__9171\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9166\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9166\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9179\,
            I => \N__9163\
        );

    \I__2126\ : CascadeMux
    port map (
            O => \N__9178\,
            I => \N__9159\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9177\,
            I => \N__9156\
        );

    \I__2124\ : InMux
    port map (
            O => \N__9174\,
            I => \N__9153\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9171\,
            I => \N__9150\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9166\,
            I => \N__9147\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__9163\,
            I => \N__9144\
        );

    \I__2120\ : InMux
    port map (
            O => \N__9162\,
            I => \N__9139\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9159\,
            I => \N__9139\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9156\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9153\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__9150\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__9147\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2114\ : Odrv4
    port map (
            O => \N__9144\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__9139\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__2112\ : InMux
    port map (
            O => \N__9126\,
            I => \N__9123\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__9123\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__2110\ : IoInMux
    port map (
            O => \N__9120\,
            I => \N__9117\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__9117\,
            I => \N__9114\
        );

    \I__2108\ : Span12Mux_s7_h
    port map (
            O => \N__9114\,
            I => \N__9111\
        );

    \I__2107\ : Span12Mux_v
    port map (
            O => \N__9111\,
            I => \N__9108\
        );

    \I__2106\ : Odrv12
    port map (
            O => \N__9108\,
            I => \CMA_c_3\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9105\,
            I => \N__9102\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9102\,
            I => \N__9072\
        );

    \I__2103\ : ClkMux
    port map (
            O => \N__9101\,
            I => \N__8997\
        );

    \I__2102\ : ClkMux
    port map (
            O => \N__9100\,
            I => \N__8997\
        );

    \I__2101\ : ClkMux
    port map (
            O => \N__9099\,
            I => \N__8997\
        );

    \I__2100\ : ClkMux
    port map (
            O => \N__9098\,
            I => \N__8997\
        );

    \I__2099\ : ClkMux
    port map (
            O => \N__9097\,
            I => \N__8997\
        );

    \I__2098\ : ClkMux
    port map (
            O => \N__9096\,
            I => \N__8997\
        );

    \I__2097\ : ClkMux
    port map (
            O => \N__9095\,
            I => \N__8997\
        );

    \I__2096\ : ClkMux
    port map (
            O => \N__9094\,
            I => \N__8997\
        );

    \I__2095\ : ClkMux
    port map (
            O => \N__9093\,
            I => \N__8997\
        );

    \I__2094\ : ClkMux
    port map (
            O => \N__9092\,
            I => \N__8997\
        );

    \I__2093\ : ClkMux
    port map (
            O => \N__9091\,
            I => \N__8997\
        );

    \I__2092\ : ClkMux
    port map (
            O => \N__9090\,
            I => \N__8997\
        );

    \I__2091\ : ClkMux
    port map (
            O => \N__9089\,
            I => \N__8997\
        );

    \I__2090\ : ClkMux
    port map (
            O => \N__9088\,
            I => \N__8997\
        );

    \I__2089\ : ClkMux
    port map (
            O => \N__9087\,
            I => \N__8997\
        );

    \I__2088\ : ClkMux
    port map (
            O => \N__9086\,
            I => \N__8997\
        );

    \I__2087\ : ClkMux
    port map (
            O => \N__9085\,
            I => \N__8997\
        );

    \I__2086\ : ClkMux
    port map (
            O => \N__9084\,
            I => \N__8997\
        );

    \I__2085\ : ClkMux
    port map (
            O => \N__9083\,
            I => \N__8997\
        );

    \I__2084\ : ClkMux
    port map (
            O => \N__9082\,
            I => \N__8997\
        );

    \I__2083\ : ClkMux
    port map (
            O => \N__9081\,
            I => \N__8997\
        );

    \I__2082\ : ClkMux
    port map (
            O => \N__9080\,
            I => \N__8997\
        );

    \I__2081\ : ClkMux
    port map (
            O => \N__9079\,
            I => \N__8997\
        );

    \I__2080\ : ClkMux
    port map (
            O => \N__9078\,
            I => \N__8997\
        );

    \I__2079\ : ClkMux
    port map (
            O => \N__9077\,
            I => \N__8997\
        );

    \I__2078\ : ClkMux
    port map (
            O => \N__9076\,
            I => \N__8997\
        );

    \I__2077\ : ClkMux
    port map (
            O => \N__9075\,
            I => \N__8997\
        );

    \I__2076\ : Glb2LocalMux
    port map (
            O => \N__9072\,
            I => \N__8997\
        );

    \I__2075\ : ClkMux
    port map (
            O => \N__9071\,
            I => \N__8997\
        );

    \I__2074\ : ClkMux
    port map (
            O => \N__9070\,
            I => \N__8997\
        );

    \I__2073\ : ClkMux
    port map (
            O => \N__9069\,
            I => \N__8997\
        );

    \I__2072\ : ClkMux
    port map (
            O => \N__9068\,
            I => \N__8997\
        );

    \I__2071\ : ClkMux
    port map (
            O => \N__9067\,
            I => \N__8997\
        );

    \I__2070\ : ClkMux
    port map (
            O => \N__9066\,
            I => \N__8997\
        );

    \I__2069\ : GlobalMux
    port map (
            O => \N__8997\,
            I => \CLK80_PLL\
        );

    \I__2068\ : CEMux
    port map (
            O => \N__8994\,
            I => \N__8990\
        );

    \I__2067\ : CEMux
    port map (
            O => \N__8993\,
            I => \N__8985\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__8990\,
            I => \N__8980\
        );

    \I__2065\ : CEMux
    port map (
            O => \N__8989\,
            I => \N__8977\
        );

    \I__2064\ : CEMux
    port map (
            O => \N__8988\,
            I => \N__8974\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__8985\,
            I => \N__8971\
        );

    \I__2062\ : CEMux
    port map (
            O => \N__8984\,
            I => \N__8968\
        );

    \I__2061\ : CEMux
    port map (
            O => \N__8983\,
            I => \N__8965\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__8980\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__8977\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__8974\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__8971\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__8968\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__8965\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2054\ : InMux
    port map (
            O => \N__8952\,
            I => \N__8948\
        );

    \I__2053\ : InMux
    port map (
            O => \N__8951\,
            I => \N__8945\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__8948\,
            I => \N__8942\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__8945\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2050\ : Odrv4
    port map (
            O => \N__8942\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2049\ : InMux
    port map (
            O => \N__8937\,
            I => \N__8934\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__8934\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__8931\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10_cascade_\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__8928\,
            I => \N__8925\
        );

    \I__2045\ : InMux
    port map (
            O => \N__8925\,
            I => \N__8918\
        );

    \I__2044\ : InMux
    port map (
            O => \N__8924\,
            I => \N__8918\
        );

    \I__2043\ : InMux
    port map (
            O => \N__8923\,
            I => \N__8915\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__8918\,
            I => \N__8912\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__8915\,
            I => \N__8908\
        );

    \I__2040\ : Span4Mux_v
    port map (
            O => \N__8912\,
            I => \N__8905\
        );

    \I__2039\ : InMux
    port map (
            O => \N__8911\,
            I => \N__8902\
        );

    \I__2038\ : Span4Mux_h
    port map (
            O => \N__8908\,
            I => \N__8899\
        );

    \I__2037\ : Sp12to4
    port map (
            O => \N__8905\,
            I => \N__8894\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__8902\,
            I => \N__8894\
        );

    \I__2035\ : Sp12to4
    port map (
            O => \N__8899\,
            I => \N__8889\
        );

    \I__2034\ : Span12Mux_h
    port map (
            O => \N__8894\,
            I => \N__8889\
        );

    \I__2033\ : Span12Mux_v
    port map (
            O => \N__8889\,
            I => \N__8886\
        );

    \I__2032\ : Odrv12
    port map (
            O => \N__8886\,
            I => \DBRn_c\
        );

    \I__2031\ : InMux
    port map (
            O => \N__8883\,
            I => \N__8877\
        );

    \I__2030\ : InMux
    port map (
            O => \N__8882\,
            I => \N__8874\
        );

    \I__2029\ : InMux
    port map (
            O => \N__8881\,
            I => \N__8869\
        );

    \I__2028\ : InMux
    port map (
            O => \N__8880\,
            I => \N__8869\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__8877\,
            I => \N__8859\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__8874\,
            I => \N__8856\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__8869\,
            I => \N__8853\
        );

    \I__2024\ : ClkMux
    port map (
            O => \N__8868\,
            I => \N__8832\
        );

    \I__2023\ : ClkMux
    port map (
            O => \N__8867\,
            I => \N__8832\
        );

    \I__2022\ : ClkMux
    port map (
            O => \N__8866\,
            I => \N__8832\
        );

    \I__2021\ : ClkMux
    port map (
            O => \N__8865\,
            I => \N__8832\
        );

    \I__2020\ : ClkMux
    port map (
            O => \N__8864\,
            I => \N__8832\
        );

    \I__2019\ : ClkMux
    port map (
            O => \N__8863\,
            I => \N__8832\
        );

    \I__2018\ : ClkMux
    port map (
            O => \N__8862\,
            I => \N__8832\
        );

    \I__2017\ : Glb2LocalMux
    port map (
            O => \N__8859\,
            I => \N__8832\
        );

    \I__2016\ : Glb2LocalMux
    port map (
            O => \N__8856\,
            I => \N__8832\
        );

    \I__2015\ : Glb2LocalMux
    port map (
            O => \N__8853\,
            I => \N__8832\
        );

    \I__2014\ : GlobalMux
    port map (
            O => \N__8832\,
            I => \N__8829\
        );

    \I__2013\ : gio2CtrlBuf
    port map (
            O => \N__8829\,
            I => \C1_c_g\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__8826\,
            I => \N__8822\
        );

    \I__2011\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8818\
        );

    \I__2010\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8814\
        );

    \I__2009\ : InMux
    port map (
            O => \N__8821\,
            I => \N__8811\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__8818\,
            I => \N__8808\
        );

    \I__2007\ : InMux
    port map (
            O => \N__8817\,
            I => \N__8805\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__8814\,
            I => \N__8802\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__8811\,
            I => \N__8799\
        );

    \I__2004\ : Span4Mux_v
    port map (
            O => \N__8808\,
            I => \N__8796\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__8805\,
            I => \N__8793\
        );

    \I__2002\ : Span4Mux_v
    port map (
            O => \N__8802\,
            I => \N__8790\
        );

    \I__2001\ : Span4Mux_v
    port map (
            O => \N__8799\,
            I => \N__8785\
        );

    \I__2000\ : Span4Mux_h
    port map (
            O => \N__8796\,
            I => \N__8785\
        );

    \I__1999\ : Span4Mux_v
    port map (
            O => \N__8793\,
            I => \N__8780\
        );

    \I__1998\ : Span4Mux_v
    port map (
            O => \N__8790\,
            I => \N__8780\
        );

    \I__1997\ : Span4Mux_v
    port map (
            O => \N__8785\,
            I => \N__8777\
        );

    \I__1996\ : Sp12to4
    port map (
            O => \N__8780\,
            I => \N__8774\
        );

    \I__1995\ : Sp12to4
    port map (
            O => \N__8777\,
            I => \N__8769\
        );

    \I__1994\ : Span12Mux_h
    port map (
            O => \N__8774\,
            I => \N__8769\
        );

    \I__1993\ : Odrv12
    port map (
            O => \N__8769\,
            I => \CLK40_PLL_i\
        );

    \I__1992\ : IoInMux
    port map (
            O => \N__8766\,
            I => \N__8763\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__8763\,
            I => \N__8758\
        );

    \I__1990\ : IoInMux
    port map (
            O => \N__8762\,
            I => \N__8755\
        );

    \I__1989\ : IoInMux
    port map (
            O => \N__8761\,
            I => \N__8752\
        );

    \I__1988\ : Span4Mux_s3_v
    port map (
            O => \N__8758\,
            I => \N__8749\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__8755\,
            I => \N__8746\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__8752\,
            I => \N__8743\
        );

    \I__1985\ : Span4Mux_h
    port map (
            O => \N__8749\,
            I => \N__8740\
        );

    \I__1984\ : Span4Mux_s3_v
    port map (
            O => \N__8746\,
            I => \N__8737\
        );

    \I__1983\ : Span4Mux_s3_h
    port map (
            O => \N__8743\,
            I => \N__8734\
        );

    \I__1982\ : Sp12to4
    port map (
            O => \N__8740\,
            I => \N__8729\
        );

    \I__1981\ : Sp12to4
    port map (
            O => \N__8737\,
            I => \N__8729\
        );

    \I__1980\ : Span4Mux_h
    port map (
            O => \N__8734\,
            I => \N__8726\
        );

    \I__1979\ : Span12Mux_h
    port map (
            O => \N__8729\,
            I => \N__8723\
        );

    \I__1978\ : Span4Mux_h
    port map (
            O => \N__8726\,
            I => \N__8720\
        );

    \I__1977\ : Span12Mux_v
    port map (
            O => \N__8723\,
            I => \N__8717\
        );

    \I__1976\ : Span4Mux_h
    port map (
            O => \N__8720\,
            I => \N__8714\
        );

    \I__1975\ : Odrv12
    port map (
            O => \N__8717\,
            I => \CLK40_PLL_i_i\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__8714\,
            I => \CLK40_PLL_i_i\
        );

    \I__1973\ : InMux
    port map (
            O => \N__8709\,
            I => \N__8696\
        );

    \I__1972\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8693\
        );

    \I__1971\ : InMux
    port map (
            O => \N__8707\,
            I => \N__8688\
        );

    \I__1970\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8688\
        );

    \I__1969\ : InMux
    port map (
            O => \N__8705\,
            I => \N__8685\
        );

    \I__1968\ : InMux
    port map (
            O => \N__8704\,
            I => \N__8682\
        );

    \I__1967\ : InMux
    port map (
            O => \N__8703\,
            I => \N__8677\
        );

    \I__1966\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8671\
        );

    \I__1965\ : InMux
    port map (
            O => \N__8701\,
            I => \N__8666\
        );

    \I__1964\ : InMux
    port map (
            O => \N__8700\,
            I => \N__8666\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8699\,
            I => \N__8663\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__8696\,
            I => \N__8655\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__8693\,
            I => \N__8655\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__8688\,
            I => \N__8655\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__8685\,
            I => \N__8652\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__8682\,
            I => \N__8649\
        );

    \I__1957\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8644\
        );

    \I__1956\ : InMux
    port map (
            O => \N__8680\,
            I => \N__8644\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__8677\,
            I => \N__8641\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8636\
        );

    \I__1953\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8636\
        );

    \I__1952\ : InMux
    port map (
            O => \N__8674\,
            I => \N__8633\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__8671\,
            I => \N__8628\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__8666\,
            I => \N__8628\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__8663\,
            I => \N__8625\
        );

    \I__1948\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8622\
        );

    \I__1947\ : Span4Mux_v
    port map (
            O => \N__8655\,
            I => \N__8617\
        );

    \I__1946\ : Span4Mux_v
    port map (
            O => \N__8652\,
            I => \N__8617\
        );

    \I__1945\ : Span4Mux_v
    port map (
            O => \N__8649\,
            I => \N__8614\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__8644\,
            I => \N__8611\
        );

    \I__1943\ : Span4Mux_v
    port map (
            O => \N__8641\,
            I => \N__8606\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__8636\,
            I => \N__8606\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__8633\,
            I => \N__8603\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__8628\,
            I => \N__8600\
        );

    \I__1939\ : Span4Mux_h
    port map (
            O => \N__8625\,
            I => \N__8595\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__8622\,
            I => \N__8595\
        );

    \I__1937\ : Span4Mux_h
    port map (
            O => \N__8617\,
            I => \N__8584\
        );

    \I__1936\ : Span4Mux_v
    port map (
            O => \N__8614\,
            I => \N__8584\
        );

    \I__1935\ : Span4Mux_v
    port map (
            O => \N__8611\,
            I => \N__8584\
        );

    \I__1934\ : Span4Mux_v
    port map (
            O => \N__8606\,
            I => \N__8584\
        );

    \I__1933\ : Span4Mux_v
    port map (
            O => \N__8603\,
            I => \N__8584\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__8600\,
            I => \N__8579\
        );

    \I__1931\ : Span4Mux_v
    port map (
            O => \N__8595\,
            I => \N__8579\
        );

    \I__1930\ : Sp12to4
    port map (
            O => \N__8584\,
            I => \N__8574\
        );

    \I__1929\ : Sp12to4
    port map (
            O => \N__8579\,
            I => \N__8574\
        );

    \I__1928\ : Span12Mux_h
    port map (
            O => \N__8574\,
            I => \N__8571\
        );

    \I__1927\ : Odrv12
    port map (
            O => \N__8571\,
            I => \RESETn_c\
        );

    \I__1926\ : IoInMux
    port map (
            O => \N__8568\,
            I => \N__8565\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__8565\,
            I => \N__8562\
        );

    \I__1924\ : Span12Mux_s3_v
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__1923\ : Odrv12
    port map (
            O => \N__8559\,
            I => \RESETn_c_i\
        );

    \I__1922\ : InMux
    port map (
            O => \N__8556\,
            I => \N__8552\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8555\,
            I => \N__8549\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__8552\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__8549\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1918\ : InMux
    port map (
            O => \N__8544\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__1917\ : InMux
    port map (
            O => \N__8541\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__8538\,
            I => \N__8535\
        );

    \I__1915\ : InMux
    port map (
            O => \N__8535\,
            I => \N__8532\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__8532\,
            I => \N__8528\
        );

    \I__1913\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8525\
        );

    \I__1912\ : Span4Mux_h
    port map (
            O => \N__8528\,
            I => \N__8522\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__8525\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__8522\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1909\ : SRMux
    port map (
            O => \N__8517\,
            I => \N__8514\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8514\,
            I => \N__8511\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__8511\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1906\ : IoInMux
    port map (
            O => \N__8508\,
            I => \N__8505\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__8505\,
            I => \N__8502\
        );

    \I__1904\ : Span4Mux_s2_v
    port map (
            O => \N__8502\,
            I => \N__8499\
        );

    \I__1903\ : Sp12to4
    port map (
            O => \N__8499\,
            I => \N__8496\
        );

    \I__1902\ : Span12Mux_h
    port map (
            O => \N__8496\,
            I => \N__8493\
        );

    \I__1901\ : Odrv12
    port map (
            O => \N__8493\,
            I => \un1_LDSn_i_0_0\
        );

    \I__1900\ : InMux
    port map (
            O => \N__8490\,
            I => \N__8486\
        );

    \I__1899\ : InMux
    port map (
            O => \N__8489\,
            I => \N__8483\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__8486\,
            I => \N__8478\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__8483\,
            I => \N__8478\
        );

    \I__1896\ : Span4Mux_v
    port map (
            O => \N__8478\,
            I => \N__8475\
        );

    \I__1895\ : Span4Mux_h
    port map (
            O => \N__8475\,
            I => \N__8471\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8468\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__8471\,
            I => \DS_ENm\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__8468\,
            I => \DS_ENm\
        );

    \I__1891\ : InMux
    port map (
            O => \N__8463\,
            I => \N__8459\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8456\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__8459\,
            I => \N__8448\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8456\,
            I => \N__8448\
        );

    \I__1887\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8441\
        );

    \I__1886\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8441\
        );

    \I__1885\ : InMux
    port map (
            O => \N__8453\,
            I => \N__8441\
        );

    \I__1884\ : Span4Mux_v
    port map (
            O => \N__8448\,
            I => \N__8438\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__8441\,
            I => \N__8435\
        );

    \I__1882\ : Span4Mux_h
    port map (
            O => \N__8438\,
            I => \N__8430\
        );

    \I__1881\ : Span4Mux_v
    port map (
            O => \N__8435\,
            I => \N__8430\
        );

    \I__1880\ : Sp12to4
    port map (
            O => \N__8430\,
            I => \N__8427\
        );

    \I__1879\ : Odrv12
    port map (
            O => \N__8427\,
            I => \A_c_0\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8424\,
            I => \N__8420\
        );

    \I__1877\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8417\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8420\,
            I => \N__8414\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8417\,
            I => \N__8408\
        );

    \I__1874\ : Span4Mux_v
    port map (
            O => \N__8414\,
            I => \N__8408\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8413\,
            I => \N__8405\
        );

    \I__1872\ : Span4Mux_h
    port map (
            O => \N__8408\,
            I => \N__8400\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8405\,
            I => \N__8400\
        );

    \I__1870\ : Sp12to4
    port map (
            O => \N__8400\,
            I => \N__8397\
        );

    \I__1869\ : Span12Mux_v
    port map (
            O => \N__8397\,
            I => \N__8394\
        );

    \I__1868\ : Odrv12
    port map (
            O => \N__8394\,
            I => \SIZ_c_0\
        );

    \I__1867\ : IoInMux
    port map (
            O => \N__8391\,
            I => \N__8388\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__8388\,
            I => \N__8385\
        );

    \I__1865\ : Span12Mux_s5_v
    port map (
            O => \N__8385\,
            I => \N__8382\
        );

    \I__1864\ : Span12Mux_h
    port map (
            O => \N__8382\,
            I => \N__8379\
        );

    \I__1863\ : Odrv12
    port map (
            O => \N__8379\,
            I => \un1_UDSn_i_0_0\
        );

    \I__1862\ : IoInMux
    port map (
            O => \N__8376\,
            I => \N__8373\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8373\,
            I => \N__8370\
        );

    \I__1860\ : Span4Mux_s0_v
    port map (
            O => \N__8370\,
            I => \N__8367\
        );

    \I__1859\ : Span4Mux_v
    port map (
            O => \N__8367\,
            I => \N__8364\
        );

    \I__1858\ : Span4Mux_v
    port map (
            O => \N__8364\,
            I => \N__8361\
        );

    \I__1857\ : Sp12to4
    port map (
            O => \N__8361\,
            I => \N__8358\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__8358\,
            I => \RASn_c\
        );

    \I__1855\ : IoInMux
    port map (
            O => \N__8355\,
            I => \N__8352\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8352\,
            I => \N__8349\
        );

    \I__1853\ : Span4Mux_s2_v
    port map (
            O => \N__8349\,
            I => \N__8346\
        );

    \I__1852\ : Sp12to4
    port map (
            O => \N__8346\,
            I => \N__8343\
        );

    \I__1851\ : Span12Mux_h
    port map (
            O => \N__8343\,
            I => \N__8340\
        );

    \I__1850\ : Odrv12
    port map (
            O => \N__8340\,
            I => \CRCSn_c\
        );

    \I__1849\ : IoInMux
    port map (
            O => \N__8337\,
            I => \N__8334\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8334\,
            I => \N__8331\
        );

    \I__1847\ : Span12Mux_s4_h
    port map (
            O => \N__8331\,
            I => \N__8328\
        );

    \I__1846\ : Span12Mux_h
    port map (
            O => \N__8328\,
            I => \N__8325\
        );

    \I__1845\ : Odrv12
    port map (
            O => \N__8325\,
            I => \WEn_c\
        );

    \I__1844\ : IoInMux
    port map (
            O => \N__8322\,
            I => \N__8319\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__8319\,
            I => \N__8316\
        );

    \I__1842\ : Span12Mux_s3_v
    port map (
            O => \N__8316\,
            I => \N__8313\
        );

    \I__1841\ : Span12Mux_h
    port map (
            O => \N__8313\,
            I => \N__8310\
        );

    \I__1840\ : Odrv12
    port map (
            O => \N__8310\,
            I => \CASn_c\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__8307\,
            I => \N__8301\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8306\,
            I => \N__8297\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8305\,
            I => \N__8294\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8304\,
            I => \N__8291\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8286\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8300\,
            I => \N__8286\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__8297\,
            I => \N__8283\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8294\,
            I => \N__8279\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__8291\,
            I => \N__8274\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8286\,
            I => \N__8274\
        );

    \I__1829\ : Span4Mux_v
    port map (
            O => \N__8283\,
            I => \N__8271\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8282\,
            I => \N__8268\
        );

    \I__1827\ : Span12Mux_h
    port map (
            O => \N__8279\,
            I => \N__8265\
        );

    \I__1826\ : Span4Mux_v
    port map (
            O => \N__8274\,
            I => \N__8262\
        );

    \I__1825\ : Span4Mux_v
    port map (
            O => \N__8271\,
            I => \N__8257\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__8268\,
            I => \N__8257\
        );

    \I__1823\ : Odrv12
    port map (
            O => \N__8265\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__8262\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__8257\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8250\,
            I => \N__8247\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8247\,
            I => \N__8243\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8246\,
            I => \N__8240\
        );

    \I__1817\ : Span4Mux_h
    port map (
            O => \N__8243\,
            I => \N__8232\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8240\,
            I => \N__8232\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__8239\,
            I => \N__8228\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__8238\,
            I => \N__8225\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__8237\,
            I => \N__8222\
        );

    \I__1812\ : Span4Mux_v
    port map (
            O => \N__8232\,
            I => \N__8216\
        );

    \I__1811\ : InMux
    port map (
            O => \N__8231\,
            I => \N__8213\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8208\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8225\,
            I => \N__8208\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8222\,
            I => \N__8200\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8221\,
            I => \N__8197\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__8220\,
            I => \N__8194\
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__8219\,
            I => \N__8188\
        );

    \I__1804\ : Sp12to4
    port map (
            O => \N__8216\,
            I => \N__8180\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8213\,
            I => \N__8180\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8208\,
            I => \N__8180\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8207\,
            I => \N__8177\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8206\,
            I => \N__8174\
        );

    \I__1799\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8169\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8204\,
            I => \N__8169\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8203\,
            I => \N__8166\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8200\,
            I => \N__8159\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__8197\,
            I => \N__8156\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8194\,
            I => \N__8151\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8193\,
            I => \N__8151\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8192\,
            I => \N__8148\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8141\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8188\,
            I => \N__8141\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8187\,
            I => \N__8141\
        );

    \I__1788\ : Span12Mux_h
    port map (
            O => \N__8180\,
            I => \N__8137\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__8177\,
            I => \N__8132\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8174\,
            I => \N__8132\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__8169\,
            I => \N__8127\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__8166\,
            I => \N__8127\
        );

    \I__1783\ : InMux
    port map (
            O => \N__8165\,
            I => \N__8118\
        );

    \I__1782\ : InMux
    port map (
            O => \N__8164\,
            I => \N__8118\
        );

    \I__1781\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8118\
        );

    \I__1780\ : InMux
    port map (
            O => \N__8162\,
            I => \N__8118\
        );

    \I__1779\ : Span4Mux_v
    port map (
            O => \N__8159\,
            I => \N__8107\
        );

    \I__1778\ : Span4Mux_h
    port map (
            O => \N__8156\,
            I => \N__8107\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__8151\,
            I => \N__8107\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__8148\,
            I => \N__8107\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__8141\,
            I => \N__8107\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8140\,
            I => \N__8104\
        );

    \I__1773\ : Odrv12
    port map (
            O => \N__8137\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1772\ : Odrv4
    port map (
            O => \N__8132\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1771\ : Odrv12
    port map (
            O => \N__8127\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8118\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__8107\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8104\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__8091\,
            I => \N__8087\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8090\,
            I => \N__8084\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8087\,
            I => \N__8081\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8084\,
            I => \N__8075\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__8081\,
            I => \N__8075\
        );

    \I__1762\ : InMux
    port map (
            O => \N__8080\,
            I => \N__8072\
        );

    \I__1761\ : Span12Mux_v
    port map (
            O => \N__8075\,
            I => \N__8068\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__8072\,
            I => \N__8065\
        );

    \I__1759\ : InMux
    port map (
            O => \N__8071\,
            I => \N__8062\
        );

    \I__1758\ : Odrv12
    port map (
            O => \N__8068\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__8065\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8062\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8055\,
            I => \N__8052\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8052\,
            I => \N__8049\
        );

    \I__1753\ : Span4Mux_v
    port map (
            O => \N__8049\,
            I => \N__8043\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8048\,
            I => \N__8040\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8047\,
            I => \N__8035\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8046\,
            I => \N__8035\
        );

    \I__1749\ : Sp12to4
    port map (
            O => \N__8043\,
            I => \N__8029\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8040\,
            I => \N__8029\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8035\,
            I => \N__8025\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__8034\,
            I => \N__8022\
        );

    \I__1745\ : Span12Mux_h
    port map (
            O => \N__8029\,
            I => \N__8019\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8028\,
            I => \N__8016\
        );

    \I__1743\ : Span4Mux_h
    port map (
            O => \N__8025\,
            I => \N__8013\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8022\,
            I => \N__8010\
        );

    \I__1741\ : Odrv12
    port map (
            O => \N__8019\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__8016\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__8013\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8010\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1737\ : IoInMux
    port map (
            O => \N__8001\,
            I => \N__7998\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__7998\,
            I => \N__7995\
        );

    \I__1735\ : Span4Mux_s0_v
    port map (
            O => \N__7995\,
            I => \N__7992\
        );

    \I__1734\ : Sp12to4
    port map (
            O => \N__7992\,
            I => \N__7989\
        );

    \I__1733\ : Span12Mux_h
    port map (
            O => \N__7989\,
            I => \N__7986\
        );

    \I__1732\ : Odrv12
    port map (
            O => \N__7986\,
            I => \CMA_c_10\
        );

    \I__1731\ : InMux
    port map (
            O => \N__7983\,
            I => \N__7979\
        );

    \I__1730\ : InMux
    port map (
            O => \N__7982\,
            I => \N__7976\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__7979\,
            I => \N__7971\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__7976\,
            I => \N__7971\
        );

    \I__1727\ : Span4Mux_h
    port map (
            O => \N__7971\,
            I => \N__7966\
        );

    \I__1726\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7961\
        );

    \I__1725\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7961\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__7966\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__7961\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1722\ : InMux
    port map (
            O => \N__7956\,
            I => \N__7950\
        );

    \I__1721\ : InMux
    port map (
            O => \N__7955\,
            I => \N__7950\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__7950\,
            I => \N__7947\
        );

    \I__1719\ : Span4Mux_v
    port map (
            O => \N__7947\,
            I => \N__7944\
        );

    \I__1718\ : Sp12to4
    port map (
            O => \N__7944\,
            I => \N__7941\
        );

    \I__1717\ : Span12Mux_h
    port map (
            O => \N__7941\,
            I => \N__7938\
        );

    \I__1716\ : Span12Mux_v
    port map (
            O => \N__7938\,
            I => \N__7935\
        );

    \I__1715\ : Odrv12
    port map (
            O => \N__7935\,
            I => \A_c_14\
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__7932\,
            I => \N__7927\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__7931\,
            I => \N__7916\
        );

    \I__1712\ : InMux
    port map (
            O => \N__7930\,
            I => \N__7906\
        );

    \I__1711\ : InMux
    port map (
            O => \N__7927\,
            I => \N__7906\
        );

    \I__1710\ : InMux
    port map (
            O => \N__7926\,
            I => \N__7906\
        );

    \I__1709\ : InMux
    port map (
            O => \N__7925\,
            I => \N__7903\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__7924\,
            I => \N__7899\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__7923\,
            I => \N__7896\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__7922\,
            I => \N__7893\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__7921\,
            I => \N__7890\
        );

    \I__1704\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7885\
        );

    \I__1703\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7882\
        );

    \I__1702\ : InMux
    port map (
            O => \N__7916\,
            I => \N__7877\
        );

    \I__1701\ : InMux
    port map (
            O => \N__7915\,
            I => \N__7874\
        );

    \I__1700\ : InMux
    port map (
            O => \N__7914\,
            I => \N__7869\
        );

    \I__1699\ : InMux
    port map (
            O => \N__7913\,
            I => \N__7869\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__7906\,
            I => \N__7864\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__7903\,
            I => \N__7864\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__7902\,
            I => \N__7861\
        );

    \I__1695\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7858\
        );

    \I__1694\ : InMux
    port map (
            O => \N__7896\,
            I => \N__7849\
        );

    \I__1693\ : InMux
    port map (
            O => \N__7893\,
            I => \N__7849\
        );

    \I__1692\ : InMux
    port map (
            O => \N__7890\,
            I => \N__7849\
        );

    \I__1691\ : InMux
    port map (
            O => \N__7889\,
            I => \N__7846\
        );

    \I__1690\ : InMux
    port map (
            O => \N__7888\,
            I => \N__7841\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__7885\,
            I => \N__7838\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__7882\,
            I => \N__7835\
        );

    \I__1687\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7830\
        );

    \I__1686\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7830\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__7877\,
            I => \N__7825\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__7874\,
            I => \N__7825\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__7869\,
            I => \N__7822\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__7864\,
            I => \N__7819\
        );

    \I__1681\ : InMux
    port map (
            O => \N__7861\,
            I => \N__7816\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__7858\,
            I => \N__7813\
        );

    \I__1679\ : InMux
    port map (
            O => \N__7857\,
            I => \N__7808\
        );

    \I__1678\ : InMux
    port map (
            O => \N__7856\,
            I => \N__7808\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__7849\,
            I => \N__7803\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__7846\,
            I => \N__7803\
        );

    \I__1675\ : InMux
    port map (
            O => \N__7845\,
            I => \N__7798\
        );

    \I__1674\ : InMux
    port map (
            O => \N__7844\,
            I => \N__7798\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__7841\,
            I => \N__7793\
        );

    \I__1672\ : Span4Mux_h
    port map (
            O => \N__7838\,
            I => \N__7793\
        );

    \I__1671\ : Span4Mux_h
    port map (
            O => \N__7835\,
            I => \N__7784\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__7830\,
            I => \N__7784\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__7825\,
            I => \N__7784\
        );

    \I__1668\ : Span4Mux_h
    port map (
            O => \N__7822\,
            I => \N__7784\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__7819\,
            I => \CPU_CYCLEm\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__7816\,
            I => \CPU_CYCLEm\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__7813\,
            I => \CPU_CYCLEm\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__7808\,
            I => \CPU_CYCLEm\
        );

    \I__1663\ : Odrv4
    port map (
            O => \N__7803\,
            I => \CPU_CYCLEm\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7798\,
            I => \CPU_CYCLEm\
        );

    \I__1661\ : Odrv4
    port map (
            O => \N__7793\,
            I => \CPU_CYCLEm\
        );

    \I__1660\ : Odrv4
    port map (
            O => \N__7784\,
            I => \CPU_CYCLEm\
        );

    \I__1659\ : InMux
    port map (
            O => \N__7767\,
            I => \N__7764\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__7764\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1657\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7758\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__7758\,
            I => \N__7755\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__7755\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7752\,
            I => \N__7748\
        );

    \I__1653\ : InMux
    port map (
            O => \N__7751\,
            I => \N__7745\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__7748\,
            I => \N__7740\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__7745\,
            I => \N__7740\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__7740\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__1649\ : InMux
    port map (
            O => \N__7737\,
            I => \bfn_11_11_0_\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7734\,
            I => \N__7730\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7727\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__7730\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__7727\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__1644\ : InMux
    port map (
            O => \N__7722\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__1643\ : InMux
    port map (
            O => \N__7719\,
            I => \N__7715\
        );

    \I__1642\ : InMux
    port map (
            O => \N__7718\,
            I => \N__7712\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7715\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__7712\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__1639\ : InMux
    port map (
            O => \N__7707\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__1638\ : InMux
    port map (
            O => \N__7704\,
            I => \N__7701\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__7701\,
            I => \N__7697\
        );

    \I__1636\ : InMux
    port map (
            O => \N__7700\,
            I => \N__7694\
        );

    \I__1635\ : Span4Mux_h
    port map (
            O => \N__7697\,
            I => \N__7691\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__7694\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1633\ : Odrv4
    port map (
            O => \N__7691\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1632\ : InMux
    port map (
            O => \N__7686\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__7683\,
            I => \N__7679\
        );

    \I__1630\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7676\
        );

    \I__1629\ : InMux
    port map (
            O => \N__7679\,
            I => \N__7673\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__7676\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__7673\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1626\ : InMux
    port map (
            O => \N__7668\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__1625\ : InMux
    port map (
            O => \N__7665\,
            I => \N__7661\
        );

    \I__1624\ : InMux
    port map (
            O => \N__7664\,
            I => \N__7658\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7661\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__7658\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1621\ : InMux
    port map (
            O => \N__7653\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__1620\ : InMux
    port map (
            O => \N__7650\,
            I => \N__7647\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7647\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i\
        );

    \I__1618\ : InMux
    port map (
            O => \N__7644\,
            I => \N__7641\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__7641\,
            I => \N__7638\
        );

    \I__1616\ : Span4Mux_h
    port map (
            O => \N__7638\,
            I => \N__7635\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__7635\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1614\ : IoInMux
    port map (
            O => \N__7632\,
            I => \N__7629\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__7629\,
            I => \N__7626\
        );

    \I__1612\ : Span12Mux_s4_v
    port map (
            O => \N__7626\,
            I => \N__7623\
        );

    \I__1611\ : Odrv12
    port map (
            O => \N__7623\,
            I => \CMA_c_2\
        );

    \I__1610\ : IoInMux
    port map (
            O => \N__7620\,
            I => \N__7617\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__7617\,
            I => \N__7614\
        );

    \I__1608\ : IoSpan4Mux
    port map (
            O => \N__7614\,
            I => \N__7611\
        );

    \I__1607\ : Sp12to4
    port map (
            O => \N__7611\,
            I => \N__7608\
        );

    \I__1606\ : Span12Mux_s7_h
    port map (
            O => \N__7608\,
            I => \N__7605\
        );

    \I__1605\ : Span12Mux_v
    port map (
            O => \N__7605\,
            I => \N__7602\
        );

    \I__1604\ : Odrv12
    port map (
            O => \N__7602\,
            I => \CMA_c_7\
        );

    \I__1603\ : InMux
    port map (
            O => \N__7599\,
            I => \N__7596\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__7596\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__1601\ : IoInMux
    port map (
            O => \N__7593\,
            I => \N__7590\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7590\,
            I => \N__7587\
        );

    \I__1599\ : IoSpan4Mux
    port map (
            O => \N__7587\,
            I => \N__7584\
        );

    \I__1598\ : IoSpan4Mux
    port map (
            O => \N__7584\,
            I => \N__7581\
        );

    \I__1597\ : Span4Mux_s3_h
    port map (
            O => \N__7581\,
            I => \N__7578\
        );

    \I__1596\ : Sp12to4
    port map (
            O => \N__7578\,
            I => \N__7575\
        );

    \I__1595\ : Span12Mux_h
    port map (
            O => \N__7575\,
            I => \N__7572\
        );

    \I__1594\ : Odrv12
    port map (
            O => \N__7572\,
            I => \CMA_c_5\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7566\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__7566\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7563\,
            I => \N__7560\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__7560\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1589\ : InMux
    port map (
            O => \N__7557\,
            I => \N__7554\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__7554\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7551\,
            I => \N__7548\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__7548\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1585\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7542\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7542\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7539\,
            I => \N__7536\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7536\,
            I => \N__7533\
        );

    \I__1581\ : Odrv12
    port map (
            O => \N__7533\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7530\,
            I => \N__7527\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__7527\,
            I => \N__7524\
        );

    \I__1578\ : Span4Mux_v
    port map (
            O => \N__7524\,
            I => \N__7521\
        );

    \I__1577\ : Sp12to4
    port map (
            O => \N__7521\,
            I => \N__7518\
        );

    \I__1576\ : Span12Mux_h
    port map (
            O => \N__7518\,
            I => \N__7515\
        );

    \I__1575\ : Odrv12
    port map (
            O => \N__7515\,
            I => \A_c_10\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7509\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7509\,
            I => \N__7506\
        );

    \I__1572\ : Span12Mux_v
    port map (
            O => \N__7506\,
            I => \N__7503\
        );

    \I__1571\ : Span12Mux_h
    port map (
            O => \N__7503\,
            I => \N__7500\
        );

    \I__1570\ : Odrv12
    port map (
            O => \N__7500\,
            I => \A_c_3\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7497\,
            I => \N__7494\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7494\,
            I => \N__7491\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__7491\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\
        );

    \I__1566\ : InMux
    port map (
            O => \N__7488\,
            I => \N__7485\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__7485\,
            I => \N__7482\
        );

    \I__1564\ : Span12Mux_v
    port map (
            O => \N__7482\,
            I => \N__7479\
        );

    \I__1563\ : Span12Mux_h
    port map (
            O => \N__7479\,
            I => \N__7476\
        );

    \I__1562\ : Odrv12
    port map (
            O => \N__7476\,
            I => \A_c_12\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7473\,
            I => \N__7470\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__7470\,
            I => \N__7467\
        );

    \I__1559\ : Span4Mux_h
    port map (
            O => \N__7467\,
            I => \N__7464\
        );

    \I__1558\ : Span4Mux_v
    port map (
            O => \N__7464\,
            I => \N__7461\
        );

    \I__1557\ : Sp12to4
    port map (
            O => \N__7461\,
            I => \N__7458\
        );

    \I__1556\ : Odrv12
    port map (
            O => \N__7458\,
            I => \A_c_5\
        );

    \I__1555\ : InMux
    port map (
            O => \N__7455\,
            I => \N__7452\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__7452\,
            I => \N__7449\
        );

    \I__1553\ : Span4Mux_v
    port map (
            O => \N__7449\,
            I => \N__7446\
        );

    \I__1552\ : Sp12to4
    port map (
            O => \N__7446\,
            I => \N__7443\
        );

    \I__1551\ : Span12Mux_h
    port map (
            O => \N__7443\,
            I => \N__7440\
        );

    \I__1550\ : Span12Mux_v
    port map (
            O => \N__7440\,
            I => \N__7437\
        );

    \I__1549\ : Odrv12
    port map (
            O => \N__7437\,
            I => \A_c_2\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7434\,
            I => \N__7431\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7431\,
            I => \N__7428\
        );

    \I__1546\ : Span12Mux_h
    port map (
            O => \N__7428\,
            I => \N__7425\
        );

    \I__1545\ : Odrv12
    port map (
            O => \N__7425\,
            I => \A_c_9\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7422\,
            I => \N__7419\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__7419\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7416\,
            I => \N__7413\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__7413\,
            I => \N__7410\
        );

    \I__1540\ : Sp12to4
    port map (
            O => \N__7410\,
            I => \N__7407\
        );

    \I__1539\ : Span12Mux_v
    port map (
            O => \N__7407\,
            I => \N__7404\
        );

    \I__1538\ : Span12Mux_h
    port map (
            O => \N__7404\,
            I => \N__7401\
        );

    \I__1537\ : Odrv12
    port map (
            O => \N__7401\,
            I => \A_c_17\
        );

    \I__1536\ : IoInMux
    port map (
            O => \N__7398\,
            I => \N__7395\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__7395\,
            I => \N__7392\
        );

    \I__1534\ : IoSpan4Mux
    port map (
            O => \N__7392\,
            I => \N__7389\
        );

    \I__1533\ : IoSpan4Mux
    port map (
            O => \N__7389\,
            I => \N__7386\
        );

    \I__1532\ : Span4Mux_s2_h
    port map (
            O => \N__7386\,
            I => \N__7383\
        );

    \I__1531\ : Sp12to4
    port map (
            O => \N__7383\,
            I => \N__7380\
        );

    \I__1530\ : Span12Mux_s9_h
    port map (
            O => \N__7380\,
            I => \N__7377\
        );

    \I__1529\ : Odrv12
    port map (
            O => \N__7377\,
            I => \CMA_c_8\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7371\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7371\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1526\ : IoInMux
    port map (
            O => \N__7368\,
            I => \N__7365\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__7365\,
            I => \N__7362\
        );

    \I__1524\ : Span12Mux_s5_h
    port map (
            O => \N__7362\,
            I => \N__7359\
        );

    \I__1523\ : Span12Mux_h
    port map (
            O => \N__7359\,
            I => \N__7356\
        );

    \I__1522\ : Odrv12
    port map (
            O => \N__7356\,
            I => \CMA_c_6\
        );

    \I__1521\ : IoInMux
    port map (
            O => \N__7353\,
            I => \N__7350\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7350\,
            I => \N__7347\
        );

    \I__1519\ : Span4Mux_s3_v
    port map (
            O => \N__7347\,
            I => \N__7344\
        );

    \I__1518\ : Span4Mux_v
    port map (
            O => \N__7344\,
            I => \N__7341\
        );

    \I__1517\ : Span4Mux_v
    port map (
            O => \N__7341\,
            I => \N__7338\
        );

    \I__1516\ : Span4Mux_h
    port map (
            O => \N__7338\,
            I => \N__7335\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__7335\,
            I => \CMA_c_0\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7329\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7329\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7326\,
            I => \N__7323\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7323\,
            I => \N__7320\
        );

    \I__1510\ : Span4Mux_h
    port map (
            O => \N__7320\,
            I => \N__7317\
        );

    \I__1509\ : Span4Mux_v
    port map (
            O => \N__7317\,
            I => \N__7314\
        );

    \I__1508\ : Sp12to4
    port map (
            O => \N__7314\,
            I => \N__7311\
        );

    \I__1507\ : Odrv12
    port map (
            O => \N__7311\,
            I => \A_c_7\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__7308\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7305\,
            I => \N__7302\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7302\,
            I => \U712_CHIP_RAM.N_289\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7299\,
            I => \N__7296\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7296\,
            I => \N__7293\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__7293\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7290\,
            I => \N__7287\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__7287\,
            I => \N__7281\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7286\,
            I => \N__7276\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7285\,
            I => \N__7276\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7284\,
            I => \N__7272\
        );

    \I__1495\ : Span4Mux_h
    port map (
            O => \N__7281\,
            I => \N__7269\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7276\,
            I => \N__7266\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7275\,
            I => \N__7263\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7272\,
            I => \U712_CHIP_RAM.N_342\
        );

    \I__1491\ : Odrv4
    port map (
            O => \N__7269\,
            I => \U712_CHIP_RAM.N_342\
        );

    \I__1490\ : Odrv4
    port map (
            O => \N__7266\,
            I => \U712_CHIP_RAM.N_342\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7263\,
            I => \U712_CHIP_RAM.N_342\
        );

    \I__1488\ : CascadeMux
    port map (
            O => \N__7254\,
            I => \N__7247\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__7253\,
            I => \N__7240\
        );

    \I__1486\ : CascadeMux
    port map (
            O => \N__7252\,
            I => \N__7234\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__7251\,
            I => \N__7231\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7227\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7247\,
            I => \N__7224\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7246\,
            I => \N__7221\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7245\,
            I => \N__7218\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7244\,
            I => \N__7209\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7243\,
            I => \N__7209\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7240\,
            I => \N__7209\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7239\,
            I => \N__7204\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7204\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7237\,
            I => \N__7197\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7234\,
            I => \N__7197\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7231\,
            I => \N__7197\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7230\,
            I => \N__7194\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7227\,
            I => \N__7191\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7224\,
            I => \N__7184\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7221\,
            I => \N__7184\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7218\,
            I => \N__7184\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7217\,
            I => \N__7181\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7216\,
            I => \N__7174\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7209\,
            I => \N__7169\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7204\,
            I => \N__7169\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7197\,
            I => \N__7164\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7194\,
            I => \N__7164\
        );

    \I__1461\ : Span4Mux_v
    port map (
            O => \N__7191\,
            I => \N__7157\
        );

    \I__1460\ : Span4Mux_v
    port map (
            O => \N__7184\,
            I => \N__7157\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7181\,
            I => \N__7157\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7180\,
            I => \N__7154\
        );

    \I__1457\ : InMux
    port map (
            O => \N__7179\,
            I => \N__7149\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7178\,
            I => \N__7149\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7177\,
            I => \N__7146\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7174\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__7169\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__7164\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__7157\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7154\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7149\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7146\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7131\,
            I => \N__7125\
        );

    \I__1446\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7122\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7129\,
            I => \N__7119\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7128\,
            I => \N__7116\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7125\,
            I => \N__7109\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__7122\,
            I => \N__7104\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7119\,
            I => \N__7104\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__7116\,
            I => \N__7101\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7115\,
            I => \N__7098\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7114\,
            I => \N__7092\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7113\,
            I => \N__7092\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7112\,
            I => \N__7089\
        );

    \I__1435\ : Span4Mux_h
    port map (
            O => \N__7109\,
            I => \N__7086\
        );

    \I__1434\ : Span4Mux_h
    port map (
            O => \N__7104\,
            I => \N__7083\
        );

    \I__1433\ : Span4Mux_h
    port map (
            O => \N__7101\,
            I => \N__7078\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7098\,
            I => \N__7078\
        );

    \I__1431\ : InMux
    port map (
            O => \N__7097\,
            I => \N__7075\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__7092\,
            I => \U712_CHIP_RAM.N_208\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7089\,
            I => \U712_CHIP_RAM.N_208\
        );

    \I__1428\ : Odrv4
    port map (
            O => \N__7086\,
            I => \U712_CHIP_RAM.N_208\
        );

    \I__1427\ : Odrv4
    port map (
            O => \N__7083\,
            I => \U712_CHIP_RAM.N_208\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__7078\,
            I => \U712_CHIP_RAM.N_208\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7075\,
            I => \U712_CHIP_RAM.N_208\
        );

    \I__1424\ : CEMux
    port map (
            O => \N__7062\,
            I => \N__7059\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__7059\,
            I => \N__7056\
        );

    \I__1422\ : Span4Mux_h
    port map (
            O => \N__7056\,
            I => \N__7053\
        );

    \I__1421\ : Odrv4
    port map (
            O => \N__7053\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0\
        );

    \I__1420\ : CascadeMux
    port map (
            O => \N__7050\,
            I => \N__7045\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7049\,
            I => \N__7035\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7048\,
            I => \N__7032\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7045\,
            I => \N__7026\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7044\,
            I => \N__7022\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7043\,
            I => \N__7010\
        );

    \I__1414\ : InMux
    port map (
            O => \N__7042\,
            I => \N__7010\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7010\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7040\,
            I => \N__7010\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7039\,
            I => \N__7010\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7038\,
            I => \N__7005\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__7035\,
            I => \N__7000\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__7032\,
            I => \N__7000\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7031\,
            I => \N__6997\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7030\,
            I => \N__6992\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7029\,
            I => \N__6992\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7026\,
            I => \N__6987\
        );

    \I__1403\ : InMux
    port map (
            O => \N__7025\,
            I => \N__6984\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__7022\,
            I => \N__6981\
        );

    \I__1401\ : InMux
    port map (
            O => \N__7021\,
            I => \N__6978\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7010\,
            I => \N__6975\
        );

    \I__1399\ : InMux
    port map (
            O => \N__7009\,
            I => \N__6972\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7008\,
            I => \N__6969\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__7005\,
            I => \N__6960\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__7000\,
            I => \N__6960\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__6997\,
            I => \N__6960\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6992\,
            I => \N__6960\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6991\,
            I => \N__6955\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6990\,
            I => \N__6955\
        );

    \I__1391\ : Span4Mux_v
    port map (
            O => \N__6987\,
            I => \N__6950\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6984\,
            I => \N__6950\
        );

    \I__1389\ : Odrv4
    port map (
            O => \N__6981\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__6978\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__6975\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__6972\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__6969\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1384\ : Odrv4
    port map (
            O => \N__6960\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__6955\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1382\ : Odrv4
    port map (
            O => \N__6950\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__6933\,
            I => \N__6926\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6921\
        );

    \I__1379\ : InMux
    port map (
            O => \N__6931\,
            I => \N__6917\
        );

    \I__1378\ : InMux
    port map (
            O => \N__6930\,
            I => \N__6914\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6929\,
            I => \N__6907\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6926\,
            I => \N__6900\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6900\
        );

    \I__1374\ : InMux
    port map (
            O => \N__6924\,
            I => \N__6900\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__6921\,
            I => \N__6897\
        );

    \I__1372\ : InMux
    port map (
            O => \N__6920\,
            I => \N__6894\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__6917\,
            I => \N__6891\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__6914\,
            I => \N__6888\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6913\,
            I => \N__6885\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__6912\,
            I => \N__6881\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__6911\,
            I => \N__6877\
        );

    \I__1366\ : InMux
    port map (
            O => \N__6910\,
            I => \N__6874\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__6907\,
            I => \N__6869\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__6900\,
            I => \N__6869\
        );

    \I__1363\ : Span4Mux_v
    port map (
            O => \N__6897\,
            I => \N__6858\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__6894\,
            I => \N__6858\
        );

    \I__1361\ : Span4Mux_v
    port map (
            O => \N__6891\,
            I => \N__6858\
        );

    \I__1360\ : Span4Mux_h
    port map (
            O => \N__6888\,
            I => \N__6858\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__6885\,
            I => \N__6858\
        );

    \I__1358\ : InMux
    port map (
            O => \N__6884\,
            I => \N__6853\
        );

    \I__1357\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6853\
        );

    \I__1356\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6848\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6877\,
            I => \N__6848\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6874\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__6869\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1352\ : Odrv4
    port map (
            O => \N__6858\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6853\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6848\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1349\ : InMux
    port map (
            O => \N__6837\,
            I => \N__6834\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__6834\,
            I => \N__6831\
        );

    \I__1347\ : Span4Mux_h
    port map (
            O => \N__6831\,
            I => \N__6828\
        );

    \I__1346\ : Odrv4
    port map (
            O => \N__6828\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_a3_0\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6825\,
            I => \N__6822\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__6822\,
            I => \N__6819\
        );

    \I__1343\ : Span12Mux_v
    port map (
            O => \N__6819\,
            I => \N__6816\
        );

    \I__1342\ : Span12Mux_h
    port map (
            O => \N__6816\,
            I => \N__6813\
        );

    \I__1341\ : Odrv12
    port map (
            O => \N__6813\,
            I => \A_c_16\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6810\,
            I => \N__6807\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__6807\,
            I => \N__6804\
        );

    \I__1338\ : Span12Mux_v
    port map (
            O => \N__6804\,
            I => \N__6801\
        );

    \I__1337\ : Span12Mux_h
    port map (
            O => \N__6801\,
            I => \N__6798\
        );

    \I__1336\ : Odrv12
    port map (
            O => \N__6798\,
            I => \A_c_18\
        );

    \I__1335\ : InMux
    port map (
            O => \N__6795\,
            I => \N__6791\
        );

    \I__1334\ : InMux
    port map (
            O => \N__6794\,
            I => \N__6788\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__6791\,
            I => \U712_CHIP_RAM.N_303\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6788\,
            I => \U712_CHIP_RAM.N_303\
        );

    \I__1331\ : InMux
    port map (
            O => \N__6783\,
            I => \N__6777\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6770\
        );

    \I__1329\ : InMux
    port map (
            O => \N__6781\,
            I => \N__6770\
        );

    \I__1328\ : InMux
    port map (
            O => \N__6780\,
            I => \N__6770\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__6777\,
            I => \U712_CHIP_RAM.N_241\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__6770\,
            I => \U712_CHIP_RAM.N_241\
        );

    \I__1325\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6761\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6764\,
            I => \N__6758\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__6761\,
            I => \N__6751\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6758\,
            I => \N__6748\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6757\,
            I => \N__6745\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6756\,
            I => \N__6742\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6755\,
            I => \N__6739\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6754\,
            I => \N__6736\
        );

    \I__1317\ : Span4Mux_v
    port map (
            O => \N__6751\,
            I => \N__6727\
        );

    \I__1316\ : Span4Mux_h
    port map (
            O => \N__6748\,
            I => \N__6727\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__6745\,
            I => \N__6727\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__6742\,
            I => \N__6727\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6739\,
            I => \N__6724\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6736\,
            I => \N__6720\
        );

    \I__1311\ : Span4Mux_v
    port map (
            O => \N__6727\,
            I => \N__6717\
        );

    \I__1310\ : Span4Mux_h
    port map (
            O => \N__6724\,
            I => \N__6714\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6711\
        );

    \I__1308\ : Odrv12
    port map (
            O => \N__6720\,
            I => \DMA_CYCLEm\
        );

    \I__1307\ : Odrv4
    port map (
            O => \N__6717\,
            I => \DMA_CYCLEm\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__6714\,
            I => \DMA_CYCLEm\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6711\,
            I => \DMA_CYCLEm\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6702\,
            I => \N__6698\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6701\,
            I => \N__6695\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__6698\,
            I => \N__6692\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__6695\,
            I => \N__6689\
        );

    \I__1300\ : Span4Mux_v
    port map (
            O => \N__6692\,
            I => \N__6685\
        );

    \I__1299\ : Span4Mux_v
    port map (
            O => \N__6689\,
            I => \N__6682\
        );

    \I__1298\ : InMux
    port map (
            O => \N__6688\,
            I => \N__6679\
        );

    \I__1297\ : Span4Mux_v
    port map (
            O => \N__6685\,
            I => \N__6676\
        );

    \I__1296\ : Span4Mux_v
    port map (
            O => \N__6682\,
            I => \N__6671\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__6679\,
            I => \N__6671\
        );

    \I__1294\ : Span4Mux_v
    port map (
            O => \N__6676\,
            I => \N__6668\
        );

    \I__1293\ : Span4Mux_v
    port map (
            O => \N__6671\,
            I => \N__6665\
        );

    \I__1292\ : Sp12to4
    port map (
            O => \N__6668\,
            I => \N__6660\
        );

    \I__1291\ : Sp12to4
    port map (
            O => \N__6665\,
            I => \N__6660\
        );

    \I__1290\ : Span12Mux_h
    port map (
            O => \N__6660\,
            I => \N__6657\
        );

    \I__1289\ : Odrv12
    port map (
            O => \N__6657\,
            I => \AWEn_c\
        );

    \I__1288\ : InMux
    port map (
            O => \N__6654\,
            I => \N__6651\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__6651\,
            I => \N__6646\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6650\,
            I => \N__6643\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6649\,
            I => \N__6640\
        );

    \I__1284\ : Span4Mux_v
    port map (
            O => \N__6646\,
            I => \N__6632\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6643\,
            I => \N__6632\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__6640\,
            I => \N__6632\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6639\,
            I => \N__6629\
        );

    \I__1280\ : Span4Mux_v
    port map (
            O => \N__6632\,
            I => \N__6626\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6629\,
            I => \N__6623\
        );

    \I__1278\ : Span4Mux_v
    port map (
            O => \N__6626\,
            I => \N__6618\
        );

    \I__1277\ : Span4Mux_v
    port map (
            O => \N__6623\,
            I => \N__6618\
        );

    \I__1276\ : Sp12to4
    port map (
            O => \N__6618\,
            I => \N__6615\
        );

    \I__1275\ : Span12Mux_h
    port map (
            O => \N__6615\,
            I => \N__6612\
        );

    \I__1274\ : Odrv12
    port map (
            O => \N__6612\,
            I => \RnW_c\
        );

    \I__1273\ : IoInMux
    port map (
            O => \N__6609\,
            I => \N__6606\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6606\,
            I => \N__6603\
        );

    \I__1271\ : IoSpan4Mux
    port map (
            O => \N__6603\,
            I => \N__6600\
        );

    \I__1270\ : Sp12to4
    port map (
            O => \N__6600\,
            I => \N__6597\
        );

    \I__1269\ : Span12Mux_s7_h
    port map (
            O => \N__6597\,
            I => \N__6594\
        );

    \I__1268\ : Span12Mux_h
    port map (
            O => \N__6594\,
            I => \N__6591\
        );

    \I__1267\ : Odrv12
    port map (
            O => \N__6591\,
            I => \N_256\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6588\,
            I => \N__6585\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6585\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1264\ : IoInMux
    port map (
            O => \N__6582\,
            I => \N__6579\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__6579\,
            I => \N__6576\
        );

    \I__1262\ : IoSpan4Mux
    port map (
            O => \N__6576\,
            I => \N__6573\
        );

    \I__1261\ : Span4Mux_s2_v
    port map (
            O => \N__6573\,
            I => \N__6570\
        );

    \I__1260\ : Span4Mux_v
    port map (
            O => \N__6570\,
            I => \N__6567\
        );

    \I__1259\ : Span4Mux_v
    port map (
            O => \N__6567\,
            I => \N__6563\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6566\,
            I => \N__6560\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__6563\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__6560\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6552\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6552\,
            I => \N__6549\
        );

    \I__1253\ : Span4Mux_h
    port map (
            O => \N__6549\,
            I => \N__6546\
        );

    \I__1252\ : Sp12to4
    port map (
            O => \N__6546\,
            I => \N__6543\
        );

    \I__1251\ : Span12Mux_v
    port map (
            O => \N__6543\,
            I => \N__6540\
        );

    \I__1250\ : Odrv12
    port map (
            O => \N__6540\,
            I => \A_c_19\
        );

    \I__1249\ : IoInMux
    port map (
            O => \N__6537\,
            I => \N__6534\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6534\,
            I => \N__6531\
        );

    \I__1247\ : IoSpan4Mux
    port map (
            O => \N__6531\,
            I => \N__6528\
        );

    \I__1246\ : Span4Mux_s1_h
    port map (
            O => \N__6528\,
            I => \N__6525\
        );

    \I__1245\ : Span4Mux_v
    port map (
            O => \N__6525\,
            I => \N__6522\
        );

    \I__1244\ : Sp12to4
    port map (
            O => \N__6522\,
            I => \N__6519\
        );

    \I__1243\ : Span12Mux_s10_h
    port map (
            O => \N__6519\,
            I => \N__6516\
        );

    \I__1242\ : Odrv12
    port map (
            O => \N__6516\,
            I => \CMA_c_9\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6513\,
            I => \N__6510\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__6510\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1239\ : IoInMux
    port map (
            O => \N__6507\,
            I => \N__6504\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6504\,
            I => \N__6501\
        );

    \I__1237\ : Span12Mux_s6_h
    port map (
            O => \N__6501\,
            I => \N__6498\
        );

    \I__1236\ : Span12Mux_h
    port map (
            O => \N__6498\,
            I => \N__6495\
        );

    \I__1235\ : Odrv12
    port map (
            O => \N__6495\,
            I => \CMA_c_4\
        );

    \I__1234\ : IoInMux
    port map (
            O => \N__6492\,
            I => \N__6489\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6489\,
            I => \N__6486\
        );

    \I__1232\ : Span4Mux_s3_v
    port map (
            O => \N__6486\,
            I => \N__6483\
        );

    \I__1231\ : Sp12to4
    port map (
            O => \N__6483\,
            I => \N__6480\
        );

    \I__1230\ : Span12Mux_h
    port map (
            O => \N__6480\,
            I => \N__6477\
        );

    \I__1229\ : Odrv12
    port map (
            O => \N__6477\,
            I => \CMA_c_1\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6471\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6471\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__1226\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6465\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6465\,
            I => \N__6462\
        );

    \I__1224\ : Span4Mux_h
    port map (
            O => \N__6462\,
            I => \N__6458\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6461\,
            I => \N__6455\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__6458\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__6455\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__6450\,
            I => \N__6447\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6447\,
            I => \N__6444\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6444\,
            I => \N__6441\
        );

    \I__1217\ : Span4Mux_h
    port map (
            O => \N__6441\,
            I => \N__6437\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6440\,
            I => \N__6434\
        );

    \I__1215\ : Odrv4
    port map (
            O => \N__6437\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6434\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6429\,
            I => \N__6426\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6426\,
            I => \N__6422\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6425\,
            I => \N__6419\
        );

    \I__1210\ : Span4Mux_v
    port map (
            O => \N__6422\,
            I => \N__6413\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6419\,
            I => \N__6413\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6410\
        );

    \I__1207\ : Span4Mux_h
    port map (
            O => \N__6413\,
            I => \N__6407\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__6410\,
            I => \N__6404\
        );

    \I__1205\ : Odrv4
    port map (
            O => \N__6407\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1204\ : Odrv4
    port map (
            O => \N__6404\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6399\,
            I => \N__6396\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__6396\,
            I => \N__6392\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6395\,
            I => \N__6387\
        );

    \I__1200\ : Span4Mux_h
    port map (
            O => \N__6392\,
            I => \N__6384\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6391\,
            I => \N__6379\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6379\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6387\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__6384\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__6379\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__6372\,
            I => \N__6369\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6369\,
            I => \N__6365\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6362\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__6365\,
            I => \N__6359\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__6362\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1189\ : Odrv4
    port map (
            O => \N__6359\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6354\,
            I => \N__6351\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__6351\,
            I => \N__6348\
        );

    \I__1186\ : Span4Mux_v
    port map (
            O => \N__6348\,
            I => \N__6345\
        );

    \I__1185\ : Sp12to4
    port map (
            O => \N__6345\,
            I => \N__6342\
        );

    \I__1184\ : Span12Mux_h
    port map (
            O => \N__6342\,
            I => \N__6339\
        );

    \I__1183\ : Odrv12
    port map (
            O => \N__6339\,
            I => \RAS1n_c\
        );

    \I__1182\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6330\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6330\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6330\,
            I => \U712_CHIP_RAM.REFRESH_SYNCZ0Z_0\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6324\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6324\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__6321\,
            I => \N__6318\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6318\,
            I => \N__6315\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6315\,
            I => \N__6312\
        );

    \I__1174\ : Odrv4
    port map (
            O => \N__6312\,
            I => \U712_CHIP_RAM.N_301\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6309\,
            I => \N__6306\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6306\,
            I => \N__6303\
        );

    \I__1171\ : Span4Mux_h
    port map (
            O => \N__6303\,
            I => \N__6300\
        );

    \I__1170\ : Odrv4
    port map (
            O => \N__6300\,
            I => \U712_CHIP_RAM.N_243\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6297\,
            I => \N__6294\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6294\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6288\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6288\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0\
        );

    \I__1165\ : CEMux
    port map (
            O => \N__6285\,
            I => \N__6281\
        );

    \I__1164\ : CEMux
    port map (
            O => \N__6284\,
            I => \N__6278\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6281\,
            I => \N__6275\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__6278\,
            I => \N__6272\
        );

    \I__1161\ : Span4Mux_v
    port map (
            O => \N__6275\,
            I => \N__6269\
        );

    \I__1160\ : Span4Mux_v
    port map (
            O => \N__6272\,
            I => \N__6266\
        );

    \I__1159\ : Span4Mux_h
    port map (
            O => \N__6269\,
            I => \N__6263\
        );

    \I__1158\ : Span4Mux_h
    port map (
            O => \N__6266\,
            I => \N__6260\
        );

    \I__1157\ : Odrv4
    port map (
            O => \N__6263\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\
        );

    \I__1156\ : Odrv4
    port map (
            O => \N__6260\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__6255\,
            I => \N__6249\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__6254\,
            I => \N__6246\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__6253\,
            I => \N__6242\
        );

    \I__1152\ : InMux
    port map (
            O => \N__6252\,
            I => \N__6235\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6226\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6226\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6245\,
            I => \N__6226\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6242\,
            I => \N__6226\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6221\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6240\,
            I => \N__6221\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6239\,
            I => \N__6217\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6238\,
            I => \N__6214\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6235\,
            I => \N__6209\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__6226\,
            I => \N__6209\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__6221\,
            I => \N__6206\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6220\,
            I => \N__6203\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6217\,
            I => \N__6197\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__6214\,
            I => \N__6188\
        );

    \I__1137\ : Span4Mux_v
    port map (
            O => \N__6209\,
            I => \N__6188\
        );

    \I__1136\ : Span4Mux_v
    port map (
            O => \N__6206\,
            I => \N__6188\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6203\,
            I => \N__6188\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6181\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6181\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6200\,
            I => \N__6181\
        );

    \I__1131\ : Odrv12
    port map (
            O => \N__6197\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1130\ : Odrv4
    port map (
            O => \N__6188\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6181\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1128\ : CascadeMux
    port map (
            O => \N__6174\,
            I => \N__6171\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6167\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6164\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6167\,
            I => \N__6158\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6164\,
            I => \N__6158\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6163\,
            I => \N__6155\
        );

    \I__1122\ : Span4Mux_v
    port map (
            O => \N__6158\,
            I => \N__6152\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6155\,
            I => \U712_CHIP_RAM.N_209\
        );

    \I__1120\ : Odrv4
    port map (
            O => \N__6152\,
            I => \U712_CHIP_RAM.N_209\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6147\,
            I => \N__6144\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6144\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_1\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__6141\,
            I => \N__6136\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__6140\,
            I => \N__6133\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__6139\,
            I => \N__6130\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6136\,
            I => \N__6122\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6111\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6130\,
            I => \N__6111\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__6129\,
            I => \N__6108\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6128\,
            I => \N__6104\
        );

    \I__1109\ : InMux
    port map (
            O => \N__6127\,
            I => \N__6099\
        );

    \I__1108\ : InMux
    port map (
            O => \N__6126\,
            I => \N__6099\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6125\,
            I => \N__6096\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6122\,
            I => \N__6093\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6121\,
            I => \N__6090\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6120\,
            I => \N__6083\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6119\,
            I => \N__6083\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6118\,
            I => \N__6083\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__6117\,
            I => \N__6078\
        );

    \I__1100\ : InMux
    port map (
            O => \N__6116\,
            I => \N__6074\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6111\,
            I => \N__6071\
        );

    \I__1098\ : InMux
    port map (
            O => \N__6108\,
            I => \N__6068\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6107\,
            I => \N__6065\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__6104\,
            I => \N__6060\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__6099\,
            I => \N__6060\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6096\,
            I => \N__6055\
        );

    \I__1093\ : Span4Mux_v
    port map (
            O => \N__6093\,
            I => \N__6055\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__6090\,
            I => \N__6050\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__6083\,
            I => \N__6050\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6047\
        );

    \I__1089\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6044\
        );

    \I__1088\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6039\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6039\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__6074\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__6071\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__6068\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__6065\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__6060\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__6055\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1080\ : Odrv4
    port map (
            O => \N__6050\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6047\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6044\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__6039\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6018\,
            I => \N__6015\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6015\,
            I => \U712_CHIP_RAM.N_227\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6012\,
            I => \N__6009\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__6009\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_2\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__6006\,
            I => \U712_CHIP_RAM.N_342_cascade_\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6003\,
            I => \N__6000\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__6000\,
            I => \N__5997\
        );

    \I__1069\ : Span4Mux_v
    port map (
            O => \N__5997\,
            I => \N__5994\
        );

    \I__1068\ : Span4Mux_v
    port map (
            O => \N__5994\,
            I => \N__5991\
        );

    \I__1067\ : Span4Mux_h
    port map (
            O => \N__5991\,
            I => \N__5988\
        );

    \I__1066\ : Sp12to4
    port map (
            O => \N__5988\,
            I => \N__5985\
        );

    \I__1065\ : Odrv12
    port map (
            O => \N__5985\,
            I => \A_c_20\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__5982\,
            I => \U712_CHIP_RAM.N_352_cascade_\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5979\,
            I => \N__5972\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5978\,
            I => \N__5972\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5977\,
            I => \N__5969\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__5972\,
            I => \U712_CHIP_RAM.N_395\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5969\,
            I => \U712_CHIP_RAM.N_395\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5964\,
            I => \N__5959\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5963\,
            I => \N__5956\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5962\,
            I => \N__5953\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__5959\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5956\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__5953\,
            I => \U712_CHIP_RAM.N_352\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__5946\,
            I => \U712_CHIP_RAM.N_293_cascade_\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5943\,
            I => \N__5938\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5935\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5932\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5938\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5935\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__5932\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__5925\,
            I => \U712_CHIP_RAM.N_99_cascade_\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5922\,
            I => \N__5918\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5921\,
            I => \N__5915\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5918\,
            I => \U712_CHIP_RAM.N_290\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5915\,
            I => \U712_CHIP_RAM.N_290\
        );

    \I__1040\ : IoInMux
    port map (
            O => \N__5910\,
            I => \N__5907\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__5907\,
            I => \N__5904\
        );

    \I__1038\ : Span4Mux_s3_v
    port map (
            O => \N__5904\,
            I => \N__5901\
        );

    \I__1037\ : Span4Mux_v
    port map (
            O => \N__5901\,
            I => \N__5898\
        );

    \I__1036\ : Span4Mux_v
    port map (
            O => \N__5898\,
            I => \N__5895\
        );

    \I__1035\ : Span4Mux_h
    port map (
            O => \N__5895\,
            I => \N__5891\
        );

    \I__1034\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5888\
        );

    \I__1033\ : Odrv4
    port map (
            O => \N__5891\,
            I => \BANK0_c\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5888\,
            I => \BANK0_c\
        );

    \I__1031\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5880\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5880\,
            I => \N__5876\
        );

    \I__1029\ : InMux
    port map (
            O => \N__5879\,
            I => \N__5873\
        );

    \I__1028\ : Span4Mux_v
    port map (
            O => \N__5876\,
            I => \N__5870\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5873\,
            I => \N__5867\
        );

    \I__1026\ : Span4Mux_h
    port map (
            O => \N__5870\,
            I => \N__5862\
        );

    \I__1025\ : Span4Mux_v
    port map (
            O => \N__5867\,
            I => \N__5862\
        );

    \I__1024\ : Sp12to4
    port map (
            O => \N__5862\,
            I => \N__5859\
        );

    \I__1023\ : Span12Mux_h
    port map (
            O => \N__5859\,
            I => \N__5856\
        );

    \I__1022\ : Span12Mux_v
    port map (
            O => \N__5856\,
            I => \N__5853\
        );

    \I__1021\ : Odrv12
    port map (
            O => \N__5853\,
            I => \TSn_c\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5850\,
            I => \N__5847\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5847\,
            I => \N__5844\
        );

    \I__1018\ : Span4Mux_v
    port map (
            O => \N__5844\,
            I => \N__5841\
        );

    \I__1017\ : Sp12to4
    port map (
            O => \N__5841\,
            I => \N__5838\
        );

    \I__1016\ : Span12Mux_h
    port map (
            O => \N__5838\,
            I => \N__5835\
        );

    \I__1015\ : Span12Mux_v
    port map (
            O => \N__5835\,
            I => \N__5832\
        );

    \I__1014\ : Odrv12
    port map (
            O => \N__5832\,
            I => \RAMSPACEn_c\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5829\,
            I => \N__5824\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5828\,
            I => \N__5821\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5827\,
            I => \N__5818\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__5824\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__5821\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5818\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5811\,
            I => \N__5806\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5810\,
            I => \N__5803\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5809\,
            I => \N__5800\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__5806\,
            I => \N__5797\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5803\,
            I => \N__5794\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__5800\,
            I => \N__5789\
        );

    \I__1001\ : Span4Mux_v
    port map (
            O => \N__5797\,
            I => \N__5786\
        );

    \I__1000\ : Span4Mux_h
    port map (
            O => \N__5794\,
            I => \N__5783\
        );

    \I__999\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5780\
        );

    \I__998\ : InMux
    port map (
            O => \N__5792\,
            I => \N__5777\
        );

    \I__997\ : Odrv4
    port map (
            O => \N__5789\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__996\ : Odrv4
    port map (
            O => \N__5786\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__995\ : Odrv4
    port map (
            O => \N__5783\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5780\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5777\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__5766\,
            I => \N__5763\
        );

    \I__991\ : InMux
    port map (
            O => \N__5763\,
            I => \N__5751\
        );

    \I__990\ : InMux
    port map (
            O => \N__5762\,
            I => \N__5751\
        );

    \I__989\ : InMux
    port map (
            O => \N__5761\,
            I => \N__5746\
        );

    \I__988\ : InMux
    port map (
            O => \N__5760\,
            I => \N__5746\
        );

    \I__987\ : InMux
    port map (
            O => \N__5759\,
            I => \N__5741\
        );

    \I__986\ : InMux
    port map (
            O => \N__5758\,
            I => \N__5738\
        );

    \I__985\ : CascadeMux
    port map (
            O => \N__5757\,
            I => \N__5734\
        );

    \I__984\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5730\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5751\,
            I => \N__5725\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5746\,
            I => \N__5725\
        );

    \I__981\ : InMux
    port map (
            O => \N__5745\,
            I => \N__5720\
        );

    \I__980\ : InMux
    port map (
            O => \N__5744\,
            I => \N__5720\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__5741\,
            I => \N__5715\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5738\,
            I => \N__5715\
        );

    \I__977\ : InMux
    port map (
            O => \N__5737\,
            I => \N__5712\
        );

    \I__976\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5709\
        );

    \I__975\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5706\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__5730\,
            I => \N__5701\
        );

    \I__973\ : Span4Mux_h
    port map (
            O => \N__5725\,
            I => \N__5701\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5720\,
            I => \N__5698\
        );

    \I__971\ : Span4Mux_h
    port map (
            O => \N__5715\,
            I => \N__5695\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5712\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__5709\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5706\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__5701\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__966\ : Odrv4
    port map (
            O => \N__5698\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__965\ : Odrv4
    port map (
            O => \N__5695\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__964\ : InMux
    port map (
            O => \N__5682\,
            I => \N__5678\
        );

    \I__963\ : CascadeMux
    port map (
            O => \N__5681\,
            I => \N__5672\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5678\,
            I => \N__5669\
        );

    \I__961\ : InMux
    port map (
            O => \N__5677\,
            I => \N__5662\
        );

    \I__960\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5662\
        );

    \I__959\ : InMux
    port map (
            O => \N__5675\,
            I => \N__5662\
        );

    \I__958\ : InMux
    port map (
            O => \N__5672\,
            I => \N__5659\
        );

    \I__957\ : Odrv4
    port map (
            O => \N__5669\,
            I => \U712_CHIP_RAM.N_359\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__5662\,
            I => \U712_CHIP_RAM.N_359\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5659\,
            I => \U712_CHIP_RAM.N_359\
        );

    \I__954\ : IoInMux
    port map (
            O => \N__5652\,
            I => \N__5649\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5649\,
            I => \N__5646\
        );

    \I__952\ : IoSpan4Mux
    port map (
            O => \N__5646\,
            I => \N__5643\
        );

    \I__951\ : Span4Mux_s3_v
    port map (
            O => \N__5643\,
            I => \N__5639\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__5642\,
            I => \N__5636\
        );

    \I__949\ : Sp12to4
    port map (
            O => \N__5639\,
            I => \N__5633\
        );

    \I__948\ : InMux
    port map (
            O => \N__5636\,
            I => \N__5630\
        );

    \I__947\ : Odrv12
    port map (
            O => \N__5633\,
            I => \DBDIR_c\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__5630\,
            I => \DBDIR_c\
        );

    \I__945\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5622\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5622\,
            I => \N__5619\
        );

    \I__943\ : Sp12to4
    port map (
            O => \N__5619\,
            I => \N__5616\
        );

    \I__942\ : Span12Mux_v
    port map (
            O => \N__5616\,
            I => \N__5613\
        );

    \I__941\ : Span12Mux_h
    port map (
            O => \N__5613\,
            I => \N__5610\
        );

    \I__940\ : Odrv12
    port map (
            O => \N__5610\,
            I => \A_c_6\
        );

    \I__939\ : InMux
    port map (
            O => \N__5607\,
            I => \N__5604\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5604\,
            I => \N__5601\
        );

    \I__937\ : Span4Mux_v
    port map (
            O => \N__5601\,
            I => \N__5598\
        );

    \I__936\ : Sp12to4
    port map (
            O => \N__5598\,
            I => \N__5595\
        );

    \I__935\ : Odrv12
    port map (
            O => \N__5595\,
            I => \A_c_13\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__5592\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\
        );

    \I__933\ : InMux
    port map (
            O => \N__5589\,
            I => \N__5586\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__5586\,
            I => \N__5583\
        );

    \I__931\ : Span4Mux_h
    port map (
            O => \N__5583\,
            I => \N__5580\
        );

    \I__930\ : Odrv4
    port map (
            O => \N__5580\,
            I => \U712_CHIP_RAM.N_257\
        );

    \I__929\ : InMux
    port map (
            O => \N__5577\,
            I => \N__5572\
        );

    \I__928\ : InMux
    port map (
            O => \N__5576\,
            I => \N__5569\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__5575\,
            I => \N__5566\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5572\,
            I => \N__5560\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__5569\,
            I => \N__5560\
        );

    \I__924\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5554\
        );

    \I__923\ : InMux
    port map (
            O => \N__5565\,
            I => \N__5554\
        );

    \I__922\ : Span4Mux_v
    port map (
            O => \N__5560\,
            I => \N__5551\
        );

    \I__921\ : InMux
    port map (
            O => \N__5559\,
            I => \N__5548\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__5554\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__919\ : Odrv4
    port map (
            O => \N__5551\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5548\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__917\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5538\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5538\,
            I => \U712_CHIP_RAM.N_205\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__5535\,
            I => \U712_CHIP_RAM.N_205_cascade_\
        );

    \I__914\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5523\
        );

    \I__913\ : InMux
    port map (
            O => \N__5531\,
            I => \N__5523\
        );

    \I__912\ : InMux
    port map (
            O => \N__5530\,
            I => \N__5520\
        );

    \I__911\ : InMux
    port map (
            O => \N__5529\,
            I => \N__5517\
        );

    \I__910\ : InMux
    port map (
            O => \N__5528\,
            I => \N__5514\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5523\,
            I => \N__5511\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__5520\,
            I => \U712_CHIP_RAM.N_216\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5517\,
            I => \U712_CHIP_RAM.N_216\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5514\,
            I => \U712_CHIP_RAM.N_216\
        );

    \I__905\ : Odrv4
    port map (
            O => \N__5511\,
            I => \U712_CHIP_RAM.N_216\
        );

    \I__904\ : InMux
    port map (
            O => \N__5502\,
            I => \N__5499\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5499\,
            I => \U712_CHIP_RAM.N_291\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__5496\,
            I => \U712_CHIP_RAM.N_291_cascade_\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__5493\,
            I => \N__5490\
        );

    \I__900\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5487\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__5487\,
            I => \N__5484\
        );

    \I__898\ : Odrv4
    port map (
            O => \N__5484\,
            I => \U712_CHIP_RAM.N_204\
        );

    \I__897\ : InMux
    port map (
            O => \N__5481\,
            I => \N__5478\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5478\,
            I => \N__5475\
        );

    \I__895\ : Span4Mux_h
    port map (
            O => \N__5475\,
            I => \N__5472\
        );

    \I__894\ : Odrv4
    port map (
            O => \N__5472\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__893\ : IoInMux
    port map (
            O => \N__5469\,
            I => \N__5466\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5466\,
            I => \N__5462\
        );

    \I__891\ : InMux
    port map (
            O => \N__5465\,
            I => \N__5459\
        );

    \I__890\ : Span4Mux_s3_v
    port map (
            O => \N__5462\,
            I => \N__5455\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__5459\,
            I => \N__5452\
        );

    \I__888\ : InMux
    port map (
            O => \N__5458\,
            I => \N__5449\
        );

    \I__887\ : Span4Mux_h
    port map (
            O => \N__5455\,
            I => \N__5445\
        );

    \I__886\ : Span4Mux_h
    port map (
            O => \N__5452\,
            I => \N__5440\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5449\,
            I => \N__5440\
        );

    \I__884\ : InMux
    port map (
            O => \N__5448\,
            I => \N__5437\
        );

    \I__883\ : Sp12to4
    port map (
            O => \N__5445\,
            I => \N__5433\
        );

    \I__882\ : Sp12to4
    port map (
            O => \N__5440\,
            I => \N__5428\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5437\,
            I => \N__5428\
        );

    \I__880\ : InMux
    port map (
            O => \N__5436\,
            I => \N__5425\
        );

    \I__879\ : Odrv12
    port map (
            O => \N__5433\,
            I => \DBENn_c\
        );

    \I__878\ : Odrv12
    port map (
            O => \N__5428\,
            I => \DBENn_c\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5425\,
            I => \DBENn_c\
        );

    \I__876\ : InMux
    port map (
            O => \N__5418\,
            I => \N__5415\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5415\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__5412\,
            I => \N__5409\
        );

    \I__873\ : InMux
    port map (
            O => \N__5409\,
            I => \N__5404\
        );

    \I__872\ : InMux
    port map (
            O => \N__5408\,
            I => \N__5401\
        );

    \I__871\ : InMux
    port map (
            O => \N__5407\,
            I => \N__5398\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5404\,
            I => \U712_BYTE_ENABLE.N_319\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5401\,
            I => \U712_BYTE_ENABLE.N_319\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5398\,
            I => \U712_BYTE_ENABLE.N_319\
        );

    \I__867\ : InMux
    port map (
            O => \N__5391\,
            I => \N__5388\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5388\,
            I => \U712_BYTE_ENABLE.N_322\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__5385\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_cascade_\
        );

    \I__864\ : InMux
    port map (
            O => \N__5382\,
            I => \N__5378\
        );

    \I__863\ : InMux
    port map (
            O => \N__5381\,
            I => \N__5375\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__5378\,
            I => \N__5372\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5375\,
            I => \N__5368\
        );

    \I__860\ : Span4Mux_v
    port map (
            O => \N__5372\,
            I => \N__5365\
        );

    \I__859\ : InMux
    port map (
            O => \N__5371\,
            I => \N__5362\
        );

    \I__858\ : Span12Mux_h
    port map (
            O => \N__5368\,
            I => \N__5359\
        );

    \I__857\ : Sp12to4
    port map (
            O => \N__5365\,
            I => \N__5354\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__5362\,
            I => \N__5354\
        );

    \I__855\ : Span12Mux_h
    port map (
            O => \N__5359\,
            I => \N__5351\
        );

    \I__854\ : Span12Mux_h
    port map (
            O => \N__5354\,
            I => \N__5348\
        );

    \I__853\ : Span12Mux_v
    port map (
            O => \N__5351\,
            I => \N__5345\
        );

    \I__852\ : Span12Mux_v
    port map (
            O => \N__5348\,
            I => \N__5342\
        );

    \I__851\ : Odrv12
    port map (
            O => \N__5345\,
            I => \CASLn_c\
        );

    \I__850\ : Odrv12
    port map (
            O => \N__5342\,
            I => \CASLn_c\
        );

    \I__849\ : IoInMux
    port map (
            O => \N__5337\,
            I => \N__5334\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__5334\,
            I => \N__5331\
        );

    \I__847\ : IoSpan4Mux
    port map (
            O => \N__5331\,
            I => \N__5328\
        );

    \I__846\ : Span4Mux_s0_h
    port map (
            O => \N__5328\,
            I => \N__5325\
        );

    \I__845\ : Span4Mux_h
    port map (
            O => \N__5325\,
            I => \N__5322\
        );

    \I__844\ : Sp12to4
    port map (
            O => \N__5322\,
            I => \N__5319\
        );

    \I__843\ : Span12Mux_v
    port map (
            O => \N__5319\,
            I => \N__5316\
        );

    \I__842\ : Span12Mux_h
    port map (
            O => \N__5316\,
            I => \N__5313\
        );

    \I__841\ : Odrv12
    port map (
            O => \N__5313\,
            I => \N_42_i\
        );

    \I__840\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5307\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5307\,
            I => \N__5303\
        );

    \I__838\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5300\
        );

    \I__837\ : Span4Mux_v
    port map (
            O => \N__5303\,
            I => \N__5296\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__5300\,
            I => \N__5293\
        );

    \I__835\ : InMux
    port map (
            O => \N__5299\,
            I => \N__5290\
        );

    \I__834\ : Span4Mux_v
    port map (
            O => \N__5296\,
            I => \N__5285\
        );

    \I__833\ : Span4Mux_v
    port map (
            O => \N__5293\,
            I => \N__5285\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5290\,
            I => \N__5282\
        );

    \I__831\ : Odrv4
    port map (
            O => \N__5285\,
            I => \REG_CYCLEm\
        );

    \I__830\ : Odrv4
    port map (
            O => \N__5282\,
            I => \REG_CYCLEm\
        );

    \I__829\ : IoInMux
    port map (
            O => \N__5277\,
            I => \N__5274\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5274\,
            I => \N__5271\
        );

    \I__827\ : IoSpan4Mux
    port map (
            O => \N__5271\,
            I => \N__5268\
        );

    \I__826\ : IoSpan4Mux
    port map (
            O => \N__5268\,
            I => \N__5265\
        );

    \I__825\ : Span4Mux_s3_v
    port map (
            O => \N__5265\,
            I => \N__5262\
        );

    \I__824\ : Sp12to4
    port map (
            O => \N__5262\,
            I => \N__5259\
        );

    \I__823\ : Span12Mux_s11_v
    port map (
            O => \N__5259\,
            I => \N__5256\
        );

    \I__822\ : Odrv12
    port map (
            O => \N__5256\,
            I => \DRDENn_c\
        );

    \I__821\ : InMux
    port map (
            O => \N__5253\,
            I => \N__5250\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5250\,
            I => \N__5247\
        );

    \I__819\ : Span4Mux_h
    port map (
            O => \N__5247\,
            I => \N__5244\
        );

    \I__818\ : Sp12to4
    port map (
            O => \N__5244\,
            I => \N__5241\
        );

    \I__817\ : Span12Mux_v
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__816\ : Odrv12
    port map (
            O => \N__5238\,
            I => \A_c_8\
        );

    \I__815\ : InMux
    port map (
            O => \N__5235\,
            I => \N__5232\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__5232\,
            I => \N__5229\
        );

    \I__813\ : Span4Mux_v
    port map (
            O => \N__5229\,
            I => \N__5226\
        );

    \I__812\ : Span4Mux_v
    port map (
            O => \N__5226\,
            I => \N__5223\
        );

    \I__811\ : Sp12to4
    port map (
            O => \N__5223\,
            I => \N__5220\
        );

    \I__810\ : Odrv12
    port map (
            O => \N__5220\,
            I => \A_c_15\
        );

    \I__809\ : IoInMux
    port map (
            O => \N__5217\,
            I => \N__5214\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5214\,
            I => \N__5211\
        );

    \I__807\ : IoSpan4Mux
    port map (
            O => \N__5211\,
            I => \N__5208\
        );

    \I__806\ : Sp12to4
    port map (
            O => \N__5208\,
            I => \N__5205\
        );

    \I__805\ : Span12Mux_s7_h
    port map (
            O => \N__5205\,
            I => \N__5202\
        );

    \I__804\ : Span12Mux_h
    port map (
            O => \N__5202\,
            I => \N__5199\
        );

    \I__803\ : Odrv12
    port map (
            O => \N__5199\,
            I => \CLK_EN_c\
        );

    \I__802\ : InMux
    port map (
            O => \N__5196\,
            I => \N__5193\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__800\ : Span4Mux_v
    port map (
            O => \N__5190\,
            I => \N__5187\
        );

    \I__799\ : Odrv4
    port map (
            O => \N__5187\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__798\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5181\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5181\,
            I => \N__5178\
        );

    \I__796\ : Odrv4
    port map (
            O => \N__5178\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0\
        );

    \I__795\ : CEMux
    port map (
            O => \N__5175\,
            I => \N__5172\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__5172\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__5169\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_\
        );

    \I__792\ : InMux
    port map (
            O => \N__5166\,
            I => \N__5161\
        );

    \I__791\ : InMux
    port map (
            O => \N__5165\,
            I => \N__5158\
        );

    \I__790\ : InMux
    port map (
            O => \N__5164\,
            I => \N__5155\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5161\,
            I => \U712_CHIP_RAM.N_393\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5158\,
            I => \U712_CHIP_RAM.N_393\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5155\,
            I => \U712_CHIP_RAM.N_393\
        );

    \I__786\ : InMux
    port map (
            O => \N__5148\,
            I => \N__5145\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5145\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0\
        );

    \I__784\ : InMux
    port map (
            O => \N__5142\,
            I => \N__5139\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5139\,
            I => \U712_CHIP_RAM.REFRESH_SYNCZ0Z_1\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__5136\,
            I => \U712_CHIP_RAM.N_227_cascade_\
        );

    \I__781\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5130\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5130\,
            I => \N__5127\
        );

    \I__779\ : Odrv4
    port map (
            O => \N__5127\,
            I => \U712_CHIP_RAM.N_226\
        );

    \I__778\ : InMux
    port map (
            O => \N__5124\,
            I => \N__5121\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5121\,
            I => \U712_CHIP_RAM.N_245\
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__5118\,
            I => \U712_CHIP_RAM.N_181_cascade_\
        );

    \I__775\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5112\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5112\,
            I => \N__5109\
        );

    \I__773\ : Span4Mux_h
    port map (
            O => \N__5109\,
            I => \N__5106\
        );

    \I__772\ : Odrv4
    port map (
            O => \N__5106\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_a4_0_a3_0\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__5103\,
            I => \U712_CHIP_RAM.N_216_cascade_\
        );

    \I__770\ : InMux
    port map (
            O => \N__5100\,
            I => \N__5097\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5097\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_0\
        );

    \I__768\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5091\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__5091\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__5088\,
            I => \N__5081\
        );

    \I__765\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5070\
        );

    \I__764\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5070\
        );

    \I__763\ : InMux
    port map (
            O => \N__5085\,
            I => \N__5070\
        );

    \I__762\ : InMux
    port map (
            O => \N__5084\,
            I => \N__5070\
        );

    \I__761\ : InMux
    port map (
            O => \N__5081\,
            I => \N__5067\
        );

    \I__760\ : InMux
    port map (
            O => \N__5080\,
            I => \N__5062\
        );

    \I__759\ : InMux
    port map (
            O => \N__5079\,
            I => \N__5062\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5070\,
            I => \N__5059\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__5067\,
            I => \U712_CHIP_RAM.N_181\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__5062\,
            I => \U712_CHIP_RAM.N_181\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__5059\,
            I => \U712_CHIP_RAM.N_181\
        );

    \I__754\ : CEMux
    port map (
            O => \N__5052\,
            I => \N__5048\
        );

    \I__753\ : CEMux
    port map (
            O => \N__5051\,
            I => \N__5045\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__5048\,
            I => \N__5040\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__5045\,
            I => \N__5040\
        );

    \I__750\ : Span4Mux_v
    port map (
            O => \N__5040\,
            I => \N__5037\
        );

    \I__749\ : Span4Mux_h
    port map (
            O => \N__5037\,
            I => \N__5034\
        );

    \I__748\ : Odrv4
    port map (
            O => \N__5034\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__5031\,
            I => \U712_CHIP_RAM.N_204_cascade_\
        );

    \I__746\ : InMux
    port map (
            O => \N__5028\,
            I => \N__5025\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__5025\,
            I => \N__5022\
        );

    \I__744\ : Odrv4
    port map (
            O => \N__5022\,
            I => \U712_CHIP_RAM.N_279_1\
        );

    \I__743\ : CascadeMux
    port map (
            O => \N__5019\,
            I => \U712_CHIP_RAM.N_279_1_cascade_\
        );

    \I__742\ : InMux
    port map (
            O => \N__5016\,
            I => \N__5012\
        );

    \I__741\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5009\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5012\,
            I => \U712_CHIP_RAM.N_398\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5009\,
            I => \U712_CHIP_RAM.N_398\
        );

    \I__738\ : CascadeMux
    port map (
            O => \N__5004\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_1_cascade_\
        );

    \I__737\ : IoInMux
    port map (
            O => \N__5001\,
            I => \N__4998\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__4998\,
            I => \N__4995\
        );

    \I__735\ : Span12Mux_s5_v
    port map (
            O => \N__4995\,
            I => \N__4992\
        );

    \I__734\ : Odrv12
    port map (
            O => \N__4992\,
            I => \VBENn_c\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__4989\,
            I => \U712_CHIP_RAM.N_209_cascade_\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__4986\,
            I => \U712_CHIP_RAM.N_359_cascade_\
        );

    \I__731\ : CascadeMux
    port map (
            O => \N__4983\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0_cascade_\
        );

    \I__730\ : CascadeMux
    port map (
            O => \N__4980\,
            I => \U712_CHIP_RAM.N_290_cascade_\
        );

    \I__729\ : InMux
    port map (
            O => \N__4977\,
            I => \N__4972\
        );

    \I__728\ : InMux
    port map (
            O => \N__4976\,
            I => \N__4969\
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__4975\,
            I => \N__4966\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4972\,
            I => \N__4963\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4969\,
            I => \N__4960\
        );

    \I__724\ : InMux
    port map (
            O => \N__4966\,
            I => \N__4957\
        );

    \I__723\ : Span4Mux_v
    port map (
            O => \N__4963\,
            I => \N__4952\
        );

    \I__722\ : Span4Mux_v
    port map (
            O => \N__4960\,
            I => \N__4952\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4957\,
            I => \N__4949\
        );

    \I__720\ : Sp12to4
    port map (
            O => \N__4952\,
            I => \N__4946\
        );

    \I__719\ : Span12Mux_v
    port map (
            O => \N__4949\,
            I => \N__4943\
        );

    \I__718\ : Span12Mux_h
    port map (
            O => \N__4946\,
            I => \N__4940\
        );

    \I__717\ : Span12Mux_h
    port map (
            O => \N__4943\,
            I => \N__4935\
        );

    \I__716\ : Span12Mux_v
    port map (
            O => \N__4940\,
            I => \N__4935\
        );

    \I__715\ : Odrv12
    port map (
            O => \N__4935\,
            I => \CASUn_c\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__4932\,
            I => \U712_BYTE_ENABLE.N_319_cascade_\
        );

    \I__713\ : IoInMux
    port map (
            O => \N__4929\,
            I => \N__4926\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4926\,
            I => \N__4923\
        );

    \I__711\ : IoSpan4Mux
    port map (
            O => \N__4923\,
            I => \N__4920\
        );

    \I__710\ : Sp12to4
    port map (
            O => \N__4920\,
            I => \N__4917\
        );

    \I__709\ : Span12Mux_s9_h
    port map (
            O => \N__4917\,
            I => \N__4914\
        );

    \I__708\ : Span12Mux_h
    port map (
            O => \N__4914\,
            I => \N__4911\
        );

    \I__707\ : Odrv12
    port map (
            O => \N__4911\,
            I => \N_43_i\
        );

    \I__706\ : InMux
    port map (
            O => \N__4908\,
            I => \N__4905\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__4905\,
            I => \N__4901\
        );

    \I__704\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4898\
        );

    \I__703\ : Span4Mux_v
    port map (
            O => \N__4901\,
            I => \N__4895\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__4898\,
            I => \N__4892\
        );

    \I__701\ : Span4Mux_v
    port map (
            O => \N__4895\,
            I => \N__4889\
        );

    \I__700\ : Span12Mux_h
    port map (
            O => \N__4892\,
            I => \N__4886\
        );

    \I__699\ : Span4Mux_v
    port map (
            O => \N__4889\,
            I => \N__4883\
        );

    \I__698\ : Span12Mux_v
    port map (
            O => \N__4886\,
            I => \N__4880\
        );

    \I__697\ : Sp12to4
    port map (
            O => \N__4883\,
            I => \N__4877\
        );

    \I__696\ : Odrv12
    port map (
            O => \N__4880\,
            I => \SIZ_c_1\
        );

    \I__695\ : Odrv12
    port map (
            O => \N__4877\,
            I => \SIZ_c_1\
        );

    \I__694\ : InMux
    port map (
            O => \N__4872\,
            I => \N__4869\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4869\,
            I => \N__4865\
        );

    \I__692\ : InMux
    port map (
            O => \N__4868\,
            I => \N__4862\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__4865\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4862\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0\
        );

    \I__689\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4854\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__4854\,
            I => \U712_BYTE_ENABLE.N_321\
        );

    \I__687\ : InMux
    port map (
            O => \N__4851\,
            I => \N__4848\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4848\,
            I => \N__4844\
        );

    \I__685\ : InMux
    port map (
            O => \N__4847\,
            I => \N__4841\
        );

    \I__684\ : Span4Mux_v
    port map (
            O => \N__4844\,
            I => \N__4836\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4841\,
            I => \N__4836\
        );

    \I__682\ : Span4Mux_h
    port map (
            O => \N__4836\,
            I => \N__4831\
        );

    \I__681\ : InMux
    port map (
            O => \N__4835\,
            I => \N__4826\
        );

    \I__680\ : InMux
    port map (
            O => \N__4834\,
            I => \N__4826\
        );

    \I__679\ : Span4Mux_v
    port map (
            O => \N__4831\,
            I => \N__4823\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__4826\,
            I => \N__4820\
        );

    \I__677\ : Span4Mux_v
    port map (
            O => \N__4823\,
            I => \N__4817\
        );

    \I__676\ : Sp12to4
    port map (
            O => \N__4820\,
            I => \N__4814\
        );

    \I__675\ : Sp12to4
    port map (
            O => \N__4817\,
            I => \N__4809\
        );

    \I__674\ : Span12Mux_v
    port map (
            O => \N__4814\,
            I => \N__4809\
        );

    \I__673\ : Odrv12
    port map (
            O => \N__4809\,
            I => \A_c_1\
        );

    \I__672\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4803\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4803\,
            I => \U712_BYTE_ENABLE.un1_CLMBEn_i_0Z0Z_0\
        );

    \I__670\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4797\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__4797\,
            I => \N__4794\
        );

    \I__668\ : Span4Mux_v
    port map (
            O => \N__4794\,
            I => \N__4791\
        );

    \I__667\ : Span4Mux_h
    port map (
            O => \N__4791\,
            I => \N__4788\
        );

    \I__666\ : Span4Mux_v
    port map (
            O => \N__4788\,
            I => \N__4785\
        );

    \I__665\ : Odrv4
    port map (
            O => \N__4785\,
            I => \TACK_EN_i_ess\
        );

    \I__664\ : InMux
    port map (
            O => \N__4782\,
            I => \N__4777\
        );

    \I__663\ : InMux
    port map (
            O => \N__4781\,
            I => \N__4774\
        );

    \I__662\ : InMux
    port map (
            O => \N__4780\,
            I => \N__4771\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4777\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4774\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__4771\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__4764\,
            I => \N__4760\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__4763\,
            I => \N__4757\
        );

    \I__656\ : InMux
    port map (
            O => \N__4760\,
            I => \N__4754\
        );

    \I__655\ : InMux
    port map (
            O => \N__4757\,
            I => \N__4751\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4754\,
            I => \N__4748\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4751\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__652\ : Odrv4
    port map (
            O => \N__4748\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__651\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4738\
        );

    \I__650\ : InMux
    port map (
            O => \N__4742\,
            I => \N__4735\
        );

    \I__649\ : InMux
    port map (
            O => \N__4741\,
            I => \N__4732\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4738\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__4735\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__4732\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__4725\,
            I => \U712_CYCLE_TERM.N_233_i_0_en_cascade_\
        );

    \I__644\ : CEMux
    port map (
            O => \N__4722\,
            I => \N__4719\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4719\,
            I => \U712_CYCLE_TERM.N_233_i_0_en_0\
        );

    \I__642\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4713\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__4713\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\
        );

    \I__640\ : InMux
    port map (
            O => \N__4710\,
            I => \N__4707\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4707\,
            I => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\
        );

    \I__638\ : CascadeMux
    port map (
            O => \N__4704\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_i_2_cascade_\
        );

    \I__637\ : InMux
    port map (
            O => \N__4701\,
            I => \N__4697\
        );

    \I__636\ : InMux
    port map (
            O => \N__4700\,
            I => \N__4694\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4697\,
            I => \N__4691\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__4694\,
            I => \CPU_TACKm\
        );

    \I__633\ : Odrv4
    port map (
            O => \N__4691\,
            I => \CPU_TACKm\
        );

    \I__632\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4682\
        );

    \I__631\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4679\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4682\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__4679\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__628\ : InMux
    port map (
            O => \N__4674\,
            I => \N__4670\
        );

    \I__627\ : InMux
    port map (
            O => \N__4673\,
            I => \N__4667\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__4670\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4667\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__624\ : CascadeMux
    port map (
            O => \N__4662\,
            I => \N__4658\
        );

    \I__623\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4655\
        );

    \I__622\ : InMux
    port map (
            O => \N__4658\,
            I => \N__4652\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__4655\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__4652\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__619\ : InMux
    port map (
            O => \N__4647\,
            I => \N__4643\
        );

    \I__618\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4640\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__4643\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4640\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__615\ : InMux
    port map (
            O => \N__4635\,
            I => \N__4632\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__4632\,
            I => \U712_CHIP_RAM.N_218\
        );

    \I__613\ : CascadeMux
    port map (
            O => \N__4629\,
            I => \U712_CHIP_RAM.N_208_cascade_\
        );

    \I__612\ : CascadeMux
    port map (
            O => \N__4626\,
            I => \U712_CHIP_RAM.N_245_cascade_\
        );

    \I__611\ : InMux
    port map (
            O => \N__4623\,
            I => \N__4620\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4620\,
            I => \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a3_0_2\
        );

    \I__609\ : InMux
    port map (
            O => \N__4617\,
            I => \N__4614\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__4614\,
            I => \N__4611\
        );

    \I__607\ : Span4Mux_v
    port map (
            O => \N__4611\,
            I => \N__4608\
        );

    \I__606\ : Sp12to4
    port map (
            O => \N__4608\,
            I => \N__4605\
        );

    \I__605\ : Odrv12
    port map (
            O => \N__4605\,
            I => \A_c_4\
        );

    \I__604\ : InMux
    port map (
            O => \N__4602\,
            I => \N__4599\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__4599\,
            I => \N__4596\
        );

    \I__602\ : Sp12to4
    port map (
            O => \N__4596\,
            I => \N__4593\
        );

    \I__601\ : Span12Mux_v
    port map (
            O => \N__4593\,
            I => \N__4590\
        );

    \I__600\ : Odrv12
    port map (
            O => \N__4590\,
            I => \A_c_11\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__4587\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\
        );

    \I__598\ : InMux
    port map (
            O => \N__4584\,
            I => \N__4581\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4581\,
            I => \U712_BYTE_ENABLE.N_327\
        );

    \I__596\ : InMux
    port map (
            O => \N__4578\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__595\ : InMux
    port map (
            O => \N__4575\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__594\ : InMux
    port map (
            O => \N__4572\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__593\ : InMux
    port map (
            O => \N__4569\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__592\ : InMux
    port map (
            O => \N__4566\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__4563\,
            I => \U712_CHIP_RAM.N_282_cascade_\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__4560\,
            I => \U712_CHIP_RAM.N_265_cascade_\
        );

    \I__589\ : InMux
    port map (
            O => \N__4557\,
            I => \N__4553\
        );

    \I__588\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4550\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4553\,
            I => \REG_TACK\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4550\,
            I => \REG_TACK\
        );

    \I__585\ : CascadeMux
    port map (
            O => \N__4545\,
            I => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\
        );

    \I__584\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4539\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__4539\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_2\
        );

    \I__582\ : IoInMux
    port map (
            O => \N__4536\,
            I => \N__4533\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__4533\,
            I => \N__4530\
        );

    \I__580\ : Span4Mux_s1_h
    port map (
            O => \N__4530\,
            I => \N__4527\
        );

    \I__579\ : Sp12to4
    port map (
            O => \N__4527\,
            I => \N__4524\
        );

    \I__578\ : Span12Mux_v
    port map (
            O => \N__4524\,
            I => \N__4520\
        );

    \I__577\ : InMux
    port map (
            O => \N__4523\,
            I => \N__4517\
        );

    \I__576\ : Odrv12
    port map (
            O => \N__4520\,
            I => \TACK_OUTn\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4517\,
            I => \TACK_OUTn\
        );

    \I__574\ : InMux
    port map (
            O => \N__4512\,
            I => \N__4508\
        );

    \I__573\ : InMux
    port map (
            O => \N__4511\,
            I => \N__4505\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4508\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4505\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__570\ : InMux
    port map (
            O => \N__4500\,
            I => \N__4496\
        );

    \I__569\ : InMux
    port map (
            O => \N__4499\,
            I => \N__4493\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4496\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4493\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__566\ : InMux
    port map (
            O => \N__4488\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__565\ : InMux
    port map (
            O => \N__4485\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__4482\,
            I => \N__4479\
        );

    \I__563\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4474\
        );

    \I__562\ : InMux
    port map (
            O => \N__4478\,
            I => \N__4469\
        );

    \I__561\ : InMux
    port map (
            O => \N__4477\,
            I => \N__4469\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4474\,
            I => \N__4460\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4469\,
            I => \N__4460\
        );

    \I__558\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4451\
        );

    \I__557\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4451\
        );

    \I__556\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4451\
        );

    \I__555\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4451\
        );

    \I__554\ : Odrv4
    port map (
            O => \N__4460\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__4451\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__552\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4438\
        );

    \I__551\ : InMux
    port map (
            O => \N__4445\,
            I => \N__4438\
        );

    \I__550\ : InMux
    port map (
            O => \N__4444\,
            I => \N__4435\
        );

    \I__549\ : InMux
    port map (
            O => \N__4443\,
            I => \N__4432\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4438\,
            I => \N__4429\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4435\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__4432\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__4429\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__544\ : InMux
    port map (
            O => \N__4422\,
            I => \N__4419\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4419\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_i_0_0_3\
        );

    \I__542\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4410\
        );

    \I__541\ : InMux
    port map (
            O => \N__4415\,
            I => \N__4406\
        );

    \I__540\ : InMux
    port map (
            O => \N__4414\,
            I => \N__4403\
        );

    \I__539\ : InMux
    port map (
            O => \N__4413\,
            I => \N__4400\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4410\,
            I => \N__4397\
        );

    \I__537\ : InMux
    port map (
            O => \N__4409\,
            I => \N__4394\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4406\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4403\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__4400\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__533\ : Odrv4
    port map (
            O => \N__4397\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__4394\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__4383\,
            I => \N__4377\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__4382\,
            I => \N__4371\
        );

    \I__529\ : InMux
    port map (
            O => \N__4381\,
            I => \N__4367\
        );

    \I__528\ : InMux
    port map (
            O => \N__4380\,
            I => \N__4364\
        );

    \I__527\ : InMux
    port map (
            O => \N__4377\,
            I => \N__4361\
        );

    \I__526\ : InMux
    port map (
            O => \N__4376\,
            I => \N__4356\
        );

    \I__525\ : InMux
    port map (
            O => \N__4375\,
            I => \N__4356\
        );

    \I__524\ : InMux
    port map (
            O => \N__4374\,
            I => \N__4349\
        );

    \I__523\ : InMux
    port map (
            O => \N__4371\,
            I => \N__4349\
        );

    \I__522\ : InMux
    port map (
            O => \N__4370\,
            I => \N__4349\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4367\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__4364\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4361\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4356\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4349\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__516\ : IoInMux
    port map (
            O => \N__4338\,
            I => \N__4335\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__514\ : IoSpan4Mux
    port map (
            O => \N__4332\,
            I => \N__4329\
        );

    \I__513\ : Sp12to4
    port map (
            O => \N__4329\,
            I => \N__4326\
        );

    \I__512\ : Span12Mux_s7_v
    port map (
            O => \N__4326\,
            I => \N__4323\
        );

    \I__511\ : Odrv12
    port map (
            O => \N__4323\,
            I => \N_40_i\
        );

    \I__510\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4317\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4317\,
            I => \U712_REG_SM.N_261\
        );

    \I__508\ : CascadeMux
    port map (
            O => \N__4314\,
            I => \N__4307\
        );

    \I__507\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4304\
        );

    \I__506\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4301\
        );

    \I__505\ : InMux
    port map (
            O => \N__4311\,
            I => \N__4298\
        );

    \I__504\ : InMux
    port map (
            O => \N__4310\,
            I => \N__4293\
        );

    \I__503\ : InMux
    port map (
            O => \N__4307\,
            I => \N__4293\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4304\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__4301\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4298\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4293\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__4284\,
            I => \N__4280\
        );

    \I__497\ : InMux
    port map (
            O => \N__4283\,
            I => \N__4275\
        );

    \I__496\ : InMux
    port map (
            O => \N__4280\,
            I => \N__4272\
        );

    \I__495\ : InMux
    port map (
            O => \N__4279\,
            I => \N__4267\
        );

    \I__494\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4267\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__4275\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__4272\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4267\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__490\ : InMux
    port map (
            O => \N__4260\,
            I => \N__4257\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4257\,
            I => \N__4249\
        );

    \I__488\ : InMux
    port map (
            O => \N__4256\,
            I => \N__4246\
        );

    \I__487\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4243\
        );

    \I__486\ : InMux
    port map (
            O => \N__4254\,
            I => \N__4240\
        );

    \I__485\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4237\
        );

    \I__484\ : InMux
    port map (
            O => \N__4252\,
            I => \N__4234\
        );

    \I__483\ : Odrv4
    port map (
            O => \N__4249\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4246\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4243\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__4240\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4237\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4234\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__477\ : IoInMux
    port map (
            O => \N__4221\,
            I => \N__4218\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4218\,
            I => \N__4215\
        );

    \I__475\ : Span12Mux_s10_h
    port map (
            O => \N__4215\,
            I => \N__4212\
        );

    \I__474\ : Span12Mux_h
    port map (
            O => \N__4212\,
            I => \N__4209\
        );

    \I__473\ : Span12Mux_v
    port map (
            O => \N__4209\,
            I => \N__4206\
        );

    \I__472\ : Odrv12
    port map (
            O => \N__4206\,
            I => \N_41_i\
        );

    \I__471\ : InMux
    port map (
            O => \N__4203\,
            I => \N__4200\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4200\,
            I => \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_0\
        );

    \I__469\ : CascadeMux
    port map (
            O => \N__4197\,
            I => \N__4194\
        );

    \I__468\ : InMux
    port map (
            O => \N__4194\,
            I => \N__4191\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4191\,
            I => \U712_REG_SM.DS_EN_RNOZ0Z_0\
        );

    \I__466\ : InMux
    port map (
            O => \N__4188\,
            I => \N__4185\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4185\,
            I => \N__4182\
        );

    \I__464\ : Odrv4
    port map (
            O => \N__4182\,
            I => \U712_REG_SM.N_314\
        );

    \I__463\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4173\
        );

    \I__462\ : InMux
    port map (
            O => \N__4178\,
            I => \N__4170\
        );

    \I__461\ : InMux
    port map (
            O => \N__4177\,
            I => \N__4167\
        );

    \I__460\ : InMux
    port map (
            O => \N__4176\,
            I => \N__4164\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__4173\,
            I => \U712_REG_SM.N_225\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__4170\,
            I => \U712_REG_SM.N_225\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4167\,
            I => \U712_REG_SM.N_225\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__4164\,
            I => \U712_REG_SM.N_225\
        );

    \I__455\ : CascadeMux
    port map (
            O => \N__4155\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_1_1_3_cascade_\
        );

    \I__454\ : CascadeMux
    port map (
            O => \N__4152\,
            I => \N__4149\
        );

    \I__453\ : InMux
    port map (
            O => \N__4149\,
            I => \N__4146\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4146\,
            I => \U712_REG_SM.N_259\
        );

    \I__451\ : CascadeMux
    port map (
            O => \N__4143\,
            I => \U712_REG_SM.N_259_cascade_\
        );

    \I__450\ : InMux
    port map (
            O => \N__4140\,
            I => \N__4137\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__4137\,
            I => \N__4133\
        );

    \I__448\ : InMux
    port map (
            O => \N__4136\,
            I => \N__4130\
        );

    \I__447\ : Odrv4
    port map (
            O => \N__4133\,
            I => \U712_REG_SM.N_236\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__4130\,
            I => \U712_REG_SM.N_236\
        );

    \I__445\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4115\
        );

    \I__444\ : InMux
    port map (
            O => \N__4124\,
            I => \N__4115\
        );

    \I__443\ : InMux
    port map (
            O => \N__4123\,
            I => \N__4110\
        );

    \I__442\ : InMux
    port map (
            O => \N__4122\,
            I => \N__4110\
        );

    \I__441\ : InMux
    port map (
            O => \N__4121\,
            I => \N__4105\
        );

    \I__440\ : InMux
    port map (
            O => \N__4120\,
            I => \N__4105\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4115\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__4110\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__4105\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__436\ : IoInMux
    port map (
            O => \N__4098\,
            I => \N__4095\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__4095\,
            I => \N__4092\
        );

    \I__434\ : Span12Mux_s7_v
    port map (
            O => \N__4092\,
            I => \N__4088\
        );

    \I__433\ : InMux
    port map (
            O => \N__4091\,
            I => \N__4084\
        );

    \I__432\ : Span12Mux_v
    port map (
            O => \N__4088\,
            I => \N__4081\
        );

    \I__431\ : InMux
    port map (
            O => \N__4087\,
            I => \N__4078\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__4084\,
            I => \N__4075\
        );

    \I__429\ : Odrv12
    port map (
            O => \N__4081\,
            I => \REGENn_c\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__4078\,
            I => \REGENn_c\
        );

    \I__427\ : Odrv12
    port map (
            O => \N__4075\,
            I => \REGENn_c\
        );

    \I__426\ : InMux
    port map (
            O => \N__4068\,
            I => \N__4065\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__4065\,
            I => \U712_REG_SM.N_307\
        );

    \I__424\ : CascadeMux
    port map (
            O => \N__4062\,
            I => \N__4059\
        );

    \I__423\ : InMux
    port map (
            O => \N__4059\,
            I => \N__4055\
        );

    \I__422\ : InMux
    port map (
            O => \N__4058\,
            I => \N__4052\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__4055\,
            I => \U712_REG_SM.N_219\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__4052\,
            I => \U712_REG_SM.N_219\
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__4047\,
            I => \N__4044\
        );

    \I__418\ : InMux
    port map (
            O => \N__4044\,
            I => \N__4041\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__4041\,
            I => \U712_REG_SM.REG_TACK_RNOZ0Z_0\
        );

    \I__416\ : CascadeMux
    port map (
            O => \N__4038\,
            I => \N__4034\
        );

    \I__415\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4031\
        );

    \I__414\ : InMux
    port map (
            O => \N__4034\,
            I => \N__4028\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__4031\,
            I => \U712_REG_SM.N_235\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__4028\,
            I => \U712_REG_SM.N_235\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__4023\,
            I => \U712_CHIP_RAM.un5_DMA_CYCLE_START_0_cascade_\
        );

    \I__410\ : CascadeMux
    port map (
            O => \N__4020\,
            I => \U712_REG_SM.N_219_cascade_\
        );

    \I__409\ : InMux
    port map (
            O => \N__4017\,
            I => \N__4014\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__4014\,
            I => \U712_REG_SM.N_304\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__4011\,
            I => \U712_REG_SM.N_304_cascade_\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__4008\,
            I => \N__4005\
        );

    \I__405\ : InMux
    port map (
            O => \N__4005\,
            I => \N__4002\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4002\,
            I => \N__3999\
        );

    \I__403\ : Odrv4
    port map (
            O => \N__3999\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_0_i_0_1\
        );

    \I__402\ : InMux
    port map (
            O => \N__3996\,
            I => \N__3993\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__3993\,
            I => \N__3989\
        );

    \I__400\ : IoInMux
    port map (
            O => \N__3992\,
            I => \N__3986\
        );

    \I__399\ : Span4Mux_v
    port map (
            O => \N__3989\,
            I => \N__3983\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3986\,
            I => \N__3980\
        );

    \I__397\ : Sp12to4
    port map (
            O => \N__3983\,
            I => \N__3977\
        );

    \I__396\ : IoSpan4Mux
    port map (
            O => \N__3980\,
            I => \N__3974\
        );

    \I__395\ : Span12Mux_h
    port map (
            O => \N__3977\,
            I => \N__3971\
        );

    \I__394\ : IoSpan4Mux
    port map (
            O => \N__3974\,
            I => \N__3968\
        );

    \I__393\ : Span12Mux_v
    port map (
            O => \N__3971\,
            I => \N__3965\
        );

    \I__392\ : IoSpan4Mux
    port map (
            O => \N__3968\,
            I => \N__3962\
        );

    \I__391\ : Odrv12
    port map (
            O => \N__3965\,
            I => \C3_c\
        );

    \I__390\ : Odrv4
    port map (
            O => \N__3962\,
            I => \C3_c\
        );

    \I__389\ : InMux
    port map (
            O => \N__3957\,
            I => \N__3954\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3954\,
            I => \N__3950\
        );

    \I__387\ : IoInMux
    port map (
            O => \N__3953\,
            I => \N__3947\
        );

    \I__386\ : Span4Mux_v
    port map (
            O => \N__3950\,
            I => \N__3944\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__3947\,
            I => \N__3941\
        );

    \I__384\ : Sp12to4
    port map (
            O => \N__3944\,
            I => \N__3938\
        );

    \I__383\ : Span4Mux_s3_h
    port map (
            O => \N__3941\,
            I => \N__3935\
        );

    \I__382\ : Span12Mux_h
    port map (
            O => \N__3938\,
            I => \N__3930\
        );

    \I__381\ : Sp12to4
    port map (
            O => \N__3935\,
            I => \N__3930\
        );

    \I__380\ : Span12Mux_v
    port map (
            O => \N__3930\,
            I => \N__3927\
        );

    \I__379\ : Odrv12
    port map (
            O => \N__3927\,
            I => \C1_c\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__3924\,
            I => \N__3921\
        );

    \I__377\ : InMux
    port map (
            O => \N__3921\,
            I => \N__3918\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__3918\,
            I => \N__3915\
        );

    \I__375\ : Span4Mux_h
    port map (
            O => \N__3915\,
            I => \N__3912\
        );

    \I__374\ : Span4Mux_v
    port map (
            O => \N__3912\,
            I => \N__3909\
        );

    \I__373\ : Span4Mux_v
    port map (
            O => \N__3909\,
            I => \N__3906\
        );

    \I__372\ : Span4Mux_v
    port map (
            O => \N__3906\,
            I => \N__3903\
        );

    \I__371\ : Odrv4
    port map (
            O => \N__3903\,
            I => \REGSPACEn_c\
        );

    \I__370\ : InMux
    port map (
            O => \N__3900\,
            I => \N__3896\
        );

    \I__369\ : InMux
    port map (
            O => \N__3899\,
            I => \N__3893\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3896\,
            I => \N__3890\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__3893\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__366\ : Odrv4
    port map (
            O => \N__3890\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__365\ : IoInMux
    port map (
            O => \N__3885\,
            I => \N__3882\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3882\,
            I => \N__3879\
        );

    \I__363\ : IoSpan4Mux
    port map (
            O => \N__3879\,
            I => \N__3876\
        );

    \I__362\ : IoSpan4Mux
    port map (
            O => \N__3876\,
            I => \N__3873\
        );

    \I__361\ : Span4Mux_s3_h
    port map (
            O => \N__3873\,
            I => \N__3870\
        );

    \I__360\ : Odrv4
    port map (
            O => \N__3870\,
            I => \N_991_i\
        );

    \I__359\ : IoInMux
    port map (
            O => \N__3867\,
            I => \N__3864\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3864\,
            I => \N__3861\
        );

    \I__357\ : IoSpan4Mux
    port map (
            O => \N__3861\,
            I => \N__3858\
        );

    \I__356\ : Span4Mux_s2_v
    port map (
            O => \N__3858\,
            I => \N__3855\
        );

    \I__355\ : Span4Mux_v
    port map (
            O => \N__3855\,
            I => \N__3852\
        );

    \I__354\ : Odrv4
    port map (
            O => \N__3852\,
            I => \CLK80_PLL_i_i\
        );

    \I__353\ : IoInMux
    port map (
            O => \N__3849\,
            I => \N__3846\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__3846\,
            I => \N__3843\
        );

    \I__351\ : Span4Mux_s3_v
    port map (
            O => \N__3843\,
            I => \N__3840\
        );

    \I__350\ : Span4Mux_h
    port map (
            O => \N__3840\,
            I => \N__3837\
        );

    \I__349\ : Span4Mux_h
    port map (
            O => \N__3837\,
            I => \N__3834\
        );

    \I__348\ : Sp12to4
    port map (
            O => \N__3834\,
            I => \N__3831\
        );

    \I__347\ : Span12Mux_s8_v
    port map (
            O => \N__3831\,
            I => \N__3828\
        );

    \I__346\ : Span12Mux_h
    port map (
            O => \N__3828\,
            I => \N__3824\
        );

    \I__345\ : InMux
    port map (
            O => \N__3827\,
            I => \N__3821\
        );

    \I__344\ : Odrv12
    port map (
            O => \N__3824\,
            I => \ASn_c\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3821\,
            I => \ASn_c\
        );

    \I__342\ : CascadeMux
    port map (
            O => \N__3816\,
            I => \U712_REG_SM.N_238_cascade_\
        );

    \I__341\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3809\
        );

    \I__340\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3806\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__3809\,
            I => \U712_REG_SM.N_238\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__3806\,
            I => \U712_REG_SM.N_238\
        );

    \I__337\ : InMux
    port map (
            O => \N__3801\,
            I => \N__3797\
        );

    \I__336\ : InMux
    port map (
            O => \N__3800\,
            I => \N__3794\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__3797\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__3794\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__333\ : CascadeMux
    port map (
            O => \N__3789\,
            I => \N__3785\
        );

    \I__332\ : InMux
    port map (
            O => \N__3788\,
            I => \N__3780\
        );

    \I__331\ : InMux
    port map (
            O => \N__3785\,
            I => \N__3780\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__3780\,
            I => \U712_REG_SM.ASn_0_sqmuxa_1\
        );

    \I__329\ : IoInMux
    port map (
            O => \N__3777\,
            I => \N__3774\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__3774\,
            I => \N__3771\
        );

    \I__327\ : IoSpan4Mux
    port map (
            O => \N__3771\,
            I => \N__3768\
        );

    \I__326\ : Span4Mux_s2_v
    port map (
            O => \N__3768\,
            I => \N__3765\
        );

    \I__325\ : Sp12to4
    port map (
            O => \N__3765\,
            I => \N__3762\
        );

    \I__324\ : Span12Mux_v
    port map (
            O => \N__3762\,
            I => \N__3759\
        );

    \I__323\ : Odrv12
    port map (
            O => \N__3759\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__8863\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__8865\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__8866\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__8867\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__8868\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__8864\
        );

    \IN_MUX_bfv_7_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_9_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8568\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3953\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3992\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4800\,
            lcout => \N_991_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9105\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101111110000"
        )
    port map (
            in0 => \N__3812\,
            in1 => \N__3801\,
            in2 => \N__3789\,
            in3 => \N__4087\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9092\,
            ce => 'H',
            sr => \N__9997\
        );

    \U712_REG_SM.ASn_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__3827\,
            in1 => \N__3788\,
            in2 => \_gnd_net_\,
            in3 => \N__4140\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9092\,
            ce => 'H',
            sr => \N__9997\
        );

    \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4176\,
            in2 => \_gnd_net_\,
            in3 => \N__3900\,
            lcout => \U712_REG_SM.N_238\,
            ltout => \U712_REG_SM.N_238_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111110111"
        )
    port map (
            in0 => \N__8709\,
            in1 => \N__3800\,
            in2 => \N__3816\,
            in3 => \N__4254\,
            lcout => \U712_REG_SM.STATE_COUNT_srsts_i_0_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100010001"
        )
    port map (
            in0 => \N__8708\,
            in1 => \N__4017\,
            in2 => \N__4038\,
            in3 => \N__3813\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9096\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4413\,
            in2 => \_gnd_net_\,
            in3 => \N__4058\,
            lcout => \U712_REG_SM.ASn_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__4278\,
            in1 => \N__4370\,
            in2 => \N__4314\,
            in3 => \N__4120\,
            lcout => \U712_REG_SM.N_225\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__4124\,
            in1 => \N__4253\,
            in2 => \N__4383\,
            in3 => \N__8880\,
            lcout => \U712_REG_SM.N_236\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__4121\,
            in1 => \N__4279\,
            in2 => \N__4382\,
            in3 => \N__4310\,
            lcout => \U712_REG_SM.N_219\,
            ltout => \U712_REG_SM.N_219_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIEMV42_4_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8707\,
            in2 => \N__4020\,
            in3 => \N__4414\,
            lcout => \U712_REG_SM.N_304\,
            ltout => \U712_REG_SM.N_304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__8706\,
            in1 => \N__4444\,
            in2 => \N__4011\,
            in3 => \N__4178\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9098\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__4125\,
            in1 => \N__4374\,
            in2 => \N__4008\,
            in3 => \N__8881\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9098\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3996\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9099\,
            ce => 'H',
            sr => \N__9990\
        );

    \U712_REG_SM.C1_SYNC_1_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4313\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9099\,
            ce => 'H',
            sr => \N__9990\
        );

    \U712_REG_SM.C1_SYNC_0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3957\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9099\,
            ce => 'H',
            sr => \N__9990\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001101"
        )
    port map (
            in0 => \N__5879\,
            in1 => \N__3899\,
            in2 => \N__3924\,
            in3 => \N__5299\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9099\,
            ce => 'H',
            sr => \N__9990\
        );

    \U712_REG_SM.C3_SYNC_1_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4381\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9099\,
            ce => 'H',
            sr => \N__9990\
        );

    \DBR_SYNC_0_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8923\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9101\,
            ce => 'H',
            sr => \N__9982\
        );

    \U712_REG_SM.REG_CYCLE_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8705\,
            in1 => \N__8911\,
            in2 => \_gnd_net_\,
            in3 => \N__4091\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10136\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6429\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9085\,
            ce => 'H',
            sr => \N__9996\
        );

    \U712_REG_SM.REG_TACK_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__4037\,
            in1 => \N__4068\,
            in2 => \N__4047\,
            in3 => \N__4557\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9085\,
            ce => 'H',
            sr => \N__9996\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4478\,
            in1 => \N__4256\,
            in2 => \_gnd_net_\,
            in3 => \N__4177\,
            lcout => \U712_REG_SM.N_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__6654\,
            in1 => \N__4409\,
            in2 => \N__4062\,
            in3 => \N__4446\,
            lcout => \U712_REG_SM.REG_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4445\,
            in1 => \N__4252\,
            in2 => \_gnd_net_\,
            in3 => \N__4477\,
            lcout => \U712_REG_SM.N_235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4499\,
            in2 => \_gnd_net_\,
            in3 => \N__4511\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un5_DMA_CYCLE_START_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__5737\,
            in1 => \N__4542\,
            in2 => \N__4023\,
            in3 => \N__6755\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9093\,
            ce => 'H',
            sr => \N__9987\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000100010"
        )
    port map (
            in0 => \N__8702\,
            in1 => \N__6201\,
            in2 => \N__5757\,
            in3 => \N__5811\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_a4_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4977\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5382\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9093\,
            ce => 'H',
            sr => \N__9987\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__6202\,
            in1 => \N__6880\,
            in2 => \_gnd_net_\,
            in3 => \N__5481\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9093\,
            ce => 'H',
            sr => \N__9987\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOO5O1_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001001000000"
        )
    port map (
            in0 => \N__7025\,
            in1 => \N__6200\,
            in2 => \N__6911\,
            in3 => \N__7177\,
            lcout => \U712_CHIP_RAM.N_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__4422\,
            in1 => \N__4179\,
            in2 => \N__4152\,
            in3 => \N__4468\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI07K21_1_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4376\,
            in1 => \N__4123\,
            in2 => \N__6450\,
            in3 => \N__6461\,
            lcout => OPEN,
            ltout => \U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_1_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI35EO1_1_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4283\,
            in2 => \N__4155\,
            in3 => \N__4311\,
            lcout => \U712_REG_SM.N_259\,
            ltout => \U712_REG_SM.N_259_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000011000000"
        )
    port map (
            in0 => \N__4467\,
            in1 => \N__8700\,
            in2 => \N__4143\,
            in3 => \N__4136\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_3_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111101110"
        )
    port map (
            in0 => \N__4122\,
            in1 => \N__4465\,
            in2 => \_gnd_net_\,
            in3 => \N__4375\,
            lcout => \U712_REG_SM.N_261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6650\,
            in1 => \N__6702\,
            in2 => \_gnd_net_\,
            in3 => \N__5733\,
            lcout => \U712_CHIP_RAM.N_257\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__4255\,
            in1 => \N__4415\,
            in2 => \N__4482\,
            in3 => \N__8882\,
            lcout => \U712_REG_SM.N_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__4466\,
            in1 => \N__8701\,
            in2 => \_gnd_net_\,
            in3 => \N__4443\,
            lcout => \U712_REG_SM.STATE_COUNT_srsts_i_i_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__6649\,
            in1 => \N__4416\,
            in2 => \_gnd_net_\,
            in3 => \N__4380\,
            lcout => \U712_REG_SM.DS_EN_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_40_i_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__4847\,
            in1 => \N__4872\,
            in2 => \N__5412\,
            in3 => \N__4584\,
            lcout => \N_40_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_2_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111111"
        )
    port map (
            in0 => \N__4320\,
            in1 => \N__4312\,
            in2 => \N__4284\,
            in3 => \N__4260\,
            lcout => \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001100"
        )
    port map (
            in0 => \N__5756\,
            in1 => \N__6239\,
            in2 => \N__6141\,
            in3 => \N__5810\,
            lcout => \U712_CHIP_RAM.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_41_i_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110011"
        )
    port map (
            in0 => \N__5465\,
            in1 => \N__4806\,
            in2 => \N__4975\,
            in3 => \N__6764\,
            lcout => \N_41_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001101"
        )
    port map (
            in0 => \N__4203\,
            in1 => \N__8474\,
            in2 => \N__4197\,
            in3 => \N__4188\,
            lcout => \DS_ENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9100\,
            ce => 'H',
            sr => \N__9959\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4701\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4556\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111110001000"
        )
    port map (
            in0 => \N__8817\,
            in1 => \N__6391\,
            in2 => \N__4545\,
            in3 => \N__4742\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9082\,
            ce => 'H',
            sr => \N__9994\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010001010000"
        )
    port map (
            in0 => \N__6390\,
            in1 => \N__4716\,
            in2 => \N__4763\,
            in3 => \N__4781\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9082\,
            ce => 'H',
            sr => \N__9994\
        );

    \U712_CHIP_RAM.CAS_SYNC_2_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4500\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9086\,
            ce => 'H',
            sr => \N__9988\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111000100"
        )
    port map (
            in0 => \N__6395\,
            in1 => \N__4523\,
            in2 => \N__8826\,
            in3 => \N__6425\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9086\,
            ce => 'H',
            sr => \N__9988\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4512\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9086\,
            ce => 'H',
            sr => \N__9988\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6125\,
            in2 => \_gnd_net_\,
            in3 => \N__6238\,
            lcout => \U712_CHIP_RAM.N_243\,
            ltout => OPEN,
            carryin => \bfn_7_9_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5084\,
            in1 => \N__6920\,
            in2 => \_gnd_net_\,
            in3 => \N__4488\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__9089\,
            ce => \N__5052\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7038\,
            in2 => \_gnd_net_\,
            in3 => \N__4485\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5085\,
            in1 => \N__7216\,
            in2 => \_gnd_net_\,
            in3 => \N__4578\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__9089\,
            ce => \N__5052\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5079\,
            in1 => \N__4661\,
            in2 => \_gnd_net_\,
            in3 => \N__4575\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__9089\,
            ce => \N__5052\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5086\,
            in1 => \N__4674\,
            in2 => \_gnd_net_\,
            in3 => \N__4572\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__9089\,
            ce => \N__5052\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5080\,
            in1 => \N__4686\,
            in2 => \_gnd_net_\,
            in3 => \N__4569\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__9089\,
            ce => \N__5052\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5087\,
            in1 => \N__4647\,
            in2 => \_gnd_net_\,
            in3 => \N__4566\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9089\,
            ce => \N__5052\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5166\,
            in1 => \N__7920\,
            in2 => \N__7251\,
            in3 => \N__7113\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_282_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__7114\,
            in1 => \N__4623\,
            in2 => \N__4563\,
            in3 => \N__6116\,
            lcout => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__7290\,
            in1 => \N__6910\,
            in2 => \N__7252\,
            in3 => \N__5577\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_265_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111001"
        )
    port map (
            in0 => \N__7049\,
            in1 => \N__7237\,
            in2 => \N__4560\,
            in3 => \N__6795\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__4700\,
            in1 => \N__4710\,
            in2 => \N__4704\,
            in3 => \N__5530\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9094\,
            ce => 'H',
            sr => \N__9969\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4685\,
            in1 => \N__4673\,
            in2 => \N__4662\,
            in3 => \N__4646\,
            lcout => \U712_CHIP_RAM.N_208\,
            ltout => \U712_CHIP_RAM.N_208_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4635\,
            in2 => \N__4629\,
            in3 => \N__6082\,
            lcout => \U712_CHIP_RAM.N_398\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIP7DI_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5576\,
            in2 => \_gnd_net_\,
            in3 => \N__7230\,
            lcout => \U712_CHIP_RAM.N_245\,
            ltout => \U712_CHIP_RAM.N_245_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6929\,
            in1 => \N__7048\,
            in2 => \N__4626\,
            in3 => \N__7913\,
            lcout => \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4617\,
            in1 => \N__4602\,
            in2 => \_gnd_net_\,
            in3 => \N__8206\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__7914\,
            in1 => \N__8207\,
            in2 => \N__4587\,
            in3 => \N__9330\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__4851\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4868\,
            lcout => \U712_BYTE_ENABLE.N_322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__5458\,
            in1 => \N__5381\,
            in2 => \_gnd_net_\,
            in3 => \N__6757\,
            lcout => \U712_BYTE_ENABLE.N_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__7925\,
            in1 => \N__8413\,
            in2 => \_gnd_net_\,
            in3 => \N__4904\,
            lcout => \U712_BYTE_ENABLE.N_319\,
            ltout => \U712_BYTE_ENABLE.N_319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_43_i_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__4976\,
            in1 => \N__5418\,
            in2 => \N__4932\,
            in3 => \N__4857\,
            lcout => \N_43_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__4908\,
            in1 => \N__8453\,
            in2 => \_gnd_net_\,
            in3 => \N__7926\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_1_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4835\,
            in1 => \N__8455\,
            in2 => \_gnd_net_\,
            in3 => \N__7930\,
            lcout => \U712_BYTE_ENABLE.N_321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_0_0_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__8454\,
            in1 => \N__4834\,
            in2 => \N__7932\,
            in3 => \N__5408\,
            lcout => \U712_BYTE_ENABLE.un1_CLMBEn_i_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__8703\,
            in1 => \N__4743\,
            in2 => \_gnd_net_\,
            in3 => \N__4782\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9079\,
            ce => \N__4722\,
            sr => \N__9995\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__8699\,
            in1 => \N__4780\,
            in2 => \N__4764\,
            in3 => \N__4741\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_233_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4725\,
            in3 => \N__10020\,
            lcout => \U712_CYCLE_TERM.N_233_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__6418\,
            in1 => \_gnd_net_\,
            in2 => \N__6372\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a3_0_a3_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5310\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7919\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7180\,
            in2 => \_gnd_net_\,
            in3 => \N__7008\,
            lcout => \U712_CHIP_RAM.N_209\,
            ltout => \U712_CHIP_RAM.N_209_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__6240\,
            in1 => \N__7275\,
            in2 => \N__4989\,
            in3 => \N__7115\,
            lcout => \U712_CHIP_RAM.N_359\,
            ltout => \U712_CHIP_RAM.N_359_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__5761\,
            in1 => \_gnd_net_\,
            in2 => \N__4986\,
            in3 => \N__5921\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010110011111100"
        )
    port map (
            in0 => \N__6128\,
            in1 => \N__5436\,
            in2 => \N__4983\,
            in3 => \N__9345\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9083\,
            ce => 'H',
            sr => \N__9979\
        );

    \U712_CHIP_RAM.REFRESH_RNILCLN6_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__5760\,
            in1 => \N__5809\,
            in2 => \N__5681\,
            in3 => \N__5028\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111111"
        )
    port map (
            in0 => \N__6241\,
            in1 => \N__7021\,
            in2 => \_gnd_net_\,
            in3 => \N__6163\,
            lcout => \U712_CHIP_RAM.N_226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7239\,
            in1 => \N__5541\,
            in2 => \N__6129\,
            in3 => \N__5529\,
            lcout => \U712_CHIP_RAM.N_290\,
            ltout => \U712_CHIP_RAM.N_290_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__5962\,
            in1 => \N__8681\,
            in2 => \N__4980\,
            in3 => \N__5016\,
            lcout => \U712_CHIP_RAM.N_181\,
            ltout => \U712_CHIP_RAM.N_181_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__5964\,
            in1 => \N__5196\,
            in2 => \N__5118\,
            in3 => \N__5115\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9087\,
            ce => \N__5051\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6220\,
            in2 => \_gnd_net_\,
            in3 => \N__7097\,
            lcout => \U712_CHIP_RAM.N_216\,
            ltout => \U712_CHIP_RAM.N_216_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001100"
        )
    port map (
            in0 => \N__7238\,
            in1 => \N__5148\,
            in2 => \N__5103\,
            in3 => \N__5100\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_2_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5559\,
            in2 => \_gnd_net_\,
            in3 => \N__5164\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__5094\,
            in1 => \N__8680\,
            in2 => \N__5088\,
            in3 => \N__5941\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9087\,
            ce => \N__5051\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_SYNC_RNI2HJQ_1_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__5142\,
            in1 => \N__6335\,
            in2 => \_gnd_net_\,
            in3 => \N__6440\,
            lcout => \U712_CHIP_RAM.N_204\,
            ltout => \U712_CHIP_RAM.N_204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIRS4M1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8675\,
            in2 => \N__5031\,
            in3 => \N__5827\,
            lcout => \U712_CHIP_RAM.N_279_1\,
            ltout => \U712_CHIP_RAM.N_279_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIGKJ14_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5793\,
            in1 => \N__5758\,
            in2 => \N__5019\,
            in3 => \N__5165\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIAQERA_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__5531\,
            in1 => \N__5015\,
            in2 => \N__5004\,
            in3 => \N__8676\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI2B8VE_3_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__7179\,
            in1 => \N__5532\,
            in2 => \N__5169\,
            in3 => \N__6837\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__6990\,
            in1 => \_gnd_net_\,
            in2 => \N__6912\,
            in3 => \N__6077\,
            lcout => \U712_CHIP_RAM.N_393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7178\,
            in1 => \N__6991\,
            in2 => \N__6117\,
            in3 => \N__6884\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_SYNC_1_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6336\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.REFRESH_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9090\,
            ce => 'H',
            sr => \N__9960\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110001010"
        )
    port map (
            in0 => \N__7043\,
            in1 => \N__7286\,
            in2 => \N__6255\,
            in3 => \N__7244\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__7243\,
            in1 => \N__6245\,
            in2 => \N__6933\,
            in3 => \N__7042\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIJC372_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__7039\,
            in1 => \N__6925\,
            in2 => \N__6253\,
            in3 => \N__7285\,
            lcout => \U712_CHIP_RAM.N_227\,
            ltout => \U712_CHIP_RAM.N_227_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111011"
        )
    port map (
            in0 => \N__6783\,
            in1 => \N__6121\,
            in2 => \N__5136\,
            in3 => \N__5133\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9095\,
            ce => \N__6284\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010100"
        )
    port map (
            in0 => \N__7041\,
            in1 => \N__6120\,
            in2 => \N__6254\,
            in3 => \N__5124\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6LG83_0_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6119\,
            in1 => \N__7112\,
            in2 => \N__7253\,
            in3 => \N__7040\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6924\,
            in2 => \_gnd_net_\,
            in3 => \N__6118\,
            lcout => \U712_CHIP_RAM.N_303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a3_0_0_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5448\,
            in2 => \_gnd_net_\,
            in3 => \N__6756\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0\,
            ltout => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_42_i_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__5407\,
            in1 => \N__5391\,
            in2 => \N__5385\,
            in3 => \N__5371\,
            lcout => \N_42_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_0_a3_0_a3_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6765\,
            in2 => \_gnd_net_\,
            in3 => \N__5306\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5253\,
            in1 => \N__5235\,
            in2 => \_gnd_net_\,
            in3 => \N__8203\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6127\,
            in1 => \N__7246\,
            in2 => \N__7050\,
            in3 => \N__7128\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9076\,
            ce => \N__5175\,
            sr => \N__9989\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6566\,
            in2 => \_gnd_net_\,
            in3 => \N__6126\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10019\,
            in2 => \_gnd_net_\,
            in3 => \N__5184\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5625\,
            in1 => \N__5607\,
            in2 => \_gnd_net_\,
            in3 => \N__8204\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8205\,
            in1 => \N__7888\,
            in2 => \N__5592\,
            in3 => \N__9387\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111110000"
        )
    port map (
            in0 => \N__5589\,
            in1 => \_gnd_net_\,
            in2 => \N__5575\,
            in3 => \N__5943\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9080\,
            ce => 'H',
            sr => \N__9970\
        );

    \U712_CHIP_RAM.DMA_CYCLE_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__6723\,
            in1 => \N__5677\,
            in2 => \N__5766\,
            in3 => \N__5502\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9080\,
            ce => 'H',
            sr => \N__9970\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICREN6_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__5676\,
            in1 => \N__5762\,
            in2 => \_gnd_net_\,
            in3 => \N__5978\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIMTA11_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000100010"
        )
    port map (
            in0 => \N__5565\,
            in1 => \N__7009\,
            in2 => \_gnd_net_\,
            in3 => \N__6931\,
            lcout => \U712_CHIP_RAM.N_205\,
            ltout => \U712_CHIP_RAM.N_205_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_0_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__7245\,
            in1 => \N__6107\,
            in2 => \N__5535\,
            in3 => \N__5528\,
            lcout => \U712_CHIP_RAM.N_291\,
            ltout => \U712_CHIP_RAM.N_291_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__5979\,
            in1 => \N__5675\,
            in2 => \N__5496\,
            in3 => \N__10018\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI06U42_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5792\,
            in1 => \N__5828\,
            in2 => \N__5493\,
            in3 => \N__5744\,
            lcout => \U712_CHIP_RAM.N_395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6913\,
            in2 => \_gnd_net_\,
            in3 => \N__6081\,
            lcout => \U712_CHIP_RAM.N_342\,
            ltout => \U712_CHIP_RAM.N_342_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7217\,
            in1 => \N__7031\,
            in2 => \N__6006\,
            in3 => \N__7129\,
            lcout => \U712_CHIP_RAM.N_352\,
            ltout => \U712_CHIP_RAM.N_352_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_1_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10358\,
            in1 => \N__6003\,
            in2 => \N__5982\,
            in3 => \N__5977\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_293_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_0_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5963\,
            in1 => \N__5745\,
            in2 => \N__5946\,
            in3 => \N__8952\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__5894\,
            in1 => \N__5942\,
            in2 => \N__5925\,
            in3 => \N__5922\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9084\,
            ce => 'H',
            sr => \N__9961\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010001"
        )
    port map (
            in0 => \N__5883\,
            in1 => \N__5850\,
            in2 => \N__7902\,
            in3 => \N__5829\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9088\,
            ce => 'H',
            sr => \N__9953\
        );

    \U712_CHIP_RAM.REFRESH_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111111011"
        )
    port map (
            in0 => \N__7704\,
            in1 => \N__7761\,
            in2 => \N__8538\,
            in3 => \N__7422\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9088\,
            ce => 'H',
            sr => \N__9953\
        );

    \U712_CHIP_RAM.DBDIR_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111010011110000"
        )
    port map (
            in0 => \N__6701\,
            in1 => \N__5759\,
            in2 => \N__5642\,
            in3 => \N__5682\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9088\,
            ce => 'H',
            sr => \N__9953\
        );

    \DBR_SYNC_1_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6468\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9088\,
            ce => 'H',
            sr => \N__9953\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6368\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9088\,
            ce => 'H',
            sr => \N__9953\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8825\,
            in2 => \_gnd_net_\,
            in3 => \N__6399\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9088\,
            ce => 'H',
            sr => \N__9953\
        );

    \U712_CHIP_RAM.REFRESH_SYNC_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9264\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6354\,
            lcout => \U712_CHIP_RAM.REFRESH_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9088\,
            ce => 'H',
            sr => \N__9953\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6327\,
            in1 => \N__6147\,
            in2 => \N__6321\,
            in3 => \N__6781\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9091\,
            ce => \N__6285\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__6782\,
            in1 => \N__6309\,
            in2 => \N__6174\,
            in3 => \N__6012\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9091\,
            ce => \N__6285\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__6297\,
            in1 => \N__6291\,
            in2 => \_gnd_net_\,
            in3 => \N__6780\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9091\,
            ce => \N__6285\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110001"
        )
    port map (
            in0 => \N__6252\,
            in1 => \N__6932\,
            in2 => \N__6139\,
            in3 => \N__6170\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110010000"
        )
    port map (
            in0 => \N__7250\,
            in1 => \N__7044\,
            in2 => \N__6140\,
            in3 => \N__6018\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR4F93_1_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__8674\,
            in1 => \N__6794\,
            in2 => \_gnd_net_\,
            in3 => \N__7131\,
            lcout => \U712_CHIP_RAM.N_241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__6754\,
            in1 => \N__6688\,
            in2 => \_gnd_net_\,
            in3 => \N__6639\,
            lcout => \N_256\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__7915\,
            in1 => \N__6588\,
            in2 => \N__8237\,
            in3 => \N__9408\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__7983\,
            in1 => \N__6555\,
            in2 => \N__7931\,
            in3 => \N__9234\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9075\,
            ce => \N__8988\,
            sr => \N__9980\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__9221\,
            in1 => \N__9678\,
            in2 => \N__9189\,
            in3 => \N__6513\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9077\,
            ce => \N__8983\,
            sr => \N__9971\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7299\,
            in1 => \N__6474\,
            in2 => \_gnd_net_\,
            in3 => \N__7332\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9077\,
            ce => \N__8983\,
            sr => \N__9971\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__7845\,
            in1 => \N__7497\,
            in2 => \N__8219\,
            in3 => \N__9357\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101000000"
        )
    port map (
            in0 => \N__7881\,
            in1 => \N__9419\,
            in2 => \N__8220\,
            in3 => \N__9162\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7844\,
            in1 => \N__7326\,
            in2 => \_gnd_net_\,
            in3 => \N__9396\,
            lcout => \U712_CHIP_RAM.N_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100110001"
        )
    port map (
            in0 => \N__8047\,
            in1 => \N__8080\,
            in2 => \N__8307\,
            in3 => \N__8187\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8300\,
            in2 => \_gnd_net_\,
            in3 => \N__8046\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8191\,
            in2 => \N__7308\,
            in3 => \N__7305\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100111011"
        )
    port map (
            in0 => \N__9420\,
            in1 => \N__8193\,
            in2 => \N__9178\,
            in3 => \N__7880\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__7030\,
            in1 => \N__7284\,
            in2 => \N__7254\,
            in3 => \N__7130\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9081\,
            ce => \N__7062\,
            sr => \N__9954\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJOND1_1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__8662\,
            in1 => \N__7029\,
            in2 => \_gnd_net_\,
            in3 => \N__6930\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6825\,
            in1 => \N__6810\,
            in2 => \_gnd_net_\,
            in3 => \N__8192\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__8164\,
            in1 => \N__8304\,
            in2 => \_gnd_net_\,
            in3 => \N__8028\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7530\,
            in1 => \N__7512\,
            in2 => \_gnd_net_\,
            in3 => \N__8163\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8165\,
            in1 => \N__7488\,
            in2 => \_gnd_net_\,
            in3 => \N__7473\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8162\,
            in1 => \N__7455\,
            in2 => \_gnd_net_\,
            in3 => \N__7434\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8071\,
            in1 => \N__8140\,
            in2 => \N__8034\,
            in3 => \N__8282\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100111111"
        )
    port map (
            in0 => \N__7751\,
            in1 => \N__7718\,
            in2 => \N__7683\,
            in3 => \N__7733\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__9528\,
            in1 => \N__7982\,
            in2 => \N__7924\,
            in3 => \N__7416\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9070\,
            ce => \N__8984\,
            sr => \N__9972\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__9218\,
            in1 => \N__9789\,
            in2 => \N__9192\,
            in3 => \N__7374\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9070\,
            ce => \N__8984\,
            sr => \N__9972\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__9217\,
            in1 => \N__9642\,
            in2 => \N__9191\,
            in3 => \N__7539\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9070\,
            ce => \N__8984\,
            sr => \N__9972\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10017\,
            in2 => \_gnd_net_\,
            in3 => \N__7650\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7889\,
            in2 => \_gnd_net_\,
            in3 => \N__8221\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__9219\,
            in1 => \N__9732\,
            in2 => \N__9188\,
            in3 => \N__7644\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9078\,
            ce => \N__8993\,
            sr => \N__9955\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__9177\,
            in1 => \N__9220\,
            in2 => \N__9846\,
            in3 => \N__7563\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9078\,
            ce => \N__8993\,
            sr => \N__9955\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7551\,
            in1 => \N__7767\,
            in2 => \_gnd_net_\,
            in3 => \N__7599\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9078\,
            ce => \N__8993\,
            sr => \N__9955\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__7857\,
            in1 => \N__7569\,
            in2 => \N__8239\,
            in3 => \N__9366\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__8231\,
            in1 => \N__7557\,
            in2 => \N__7923\,
            in3 => \N__9318\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111010101"
        )
    port map (
            in0 => \N__7969\,
            in1 => \N__7956\,
            in2 => \N__7921\,
            in3 => \N__10152\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__7856\,
            in1 => \N__7545\,
            in2 => \N__8238\,
            in3 => \N__9375\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__7970\,
            in1 => \N__7955\,
            in2 => \N__7922\,
            in3 => \N__10151\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8555\,
            in2 => \_gnd_net_\,
            in3 => \N__7664\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7752\,
            in2 => \_gnd_net_\,
            in3 => \N__7737\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__8862\,
            ce => 'H',
            sr => \N__8517\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7734\,
            in2 => \_gnd_net_\,
            in3 => \N__7722\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__8862\,
            ce => 'H',
            sr => \N__8517\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7719\,
            in2 => \_gnd_net_\,
            in3 => \N__7707\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__8862\,
            ce => 'H',
            sr => \N__8517\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7700\,
            in2 => \_gnd_net_\,
            in3 => \N__7686\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__8862\,
            ce => 'H',
            sr => \N__8517\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7682\,
            in2 => \_gnd_net_\,
            in3 => \N__7668\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__8862\,
            ce => 'H',
            sr => \N__8517\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7665\,
            in2 => \_gnd_net_\,
            in3 => \N__7653\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__8862\,
            ce => 'H',
            sr => \N__8517\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8556\,
            in2 => \_gnd_net_\,
            in3 => \N__8544\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__8862\,
            ce => 'H',
            sr => \N__8517\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8531\,
            in2 => \_gnd_net_\,
            in3 => \N__8541\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8862\,
            ce => 'H',
            sr => \N__8517\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__8489\,
            in1 => \N__8463\,
            in2 => \_gnd_net_\,
            in3 => \N__8423\,
            lcout => \un1_LDSn_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__8490\,
            in1 => \N__8462\,
            in2 => \_gnd_net_\,
            in3 => \N__8424\,
            lcout => \un1_UDSn_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RASn_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8305\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9066\,
            ce => 'H',
            sr => \N__9986\
        );

    \U712_CHIP_RAM.CRCSn_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8090\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9067\,
            ce => 'H',
            sr => \N__9978\
        );

    \U712_CHIP_RAM.WEn_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8048\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9068\,
            ce => 'H',
            sr => \N__9968\
        );

    \U712_CHIP_RAM.CASn_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8250\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9068\,
            ce => 'H',
            sr => \N__9968\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8306\,
            in1 => \N__8246\,
            in2 => \N__8091\,
            in3 => \N__8055\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9069\,
            ce => \N__8989\,
            sr => \N__9958\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9629\,
            in1 => \N__10359\,
            in2 => \_gnd_net_\,
            in3 => \N__9260\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10132\,
            ce => \N__10086\,
            sr => \N__9952\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__9222\,
            in1 => \N__9777\,
            in2 => \N__9190\,
            in3 => \N__9126\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9071\,
            ce => \N__8994\,
            sr => \N__9949\
        );

    \U712_CHIP_RAM.DMA_A20_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__10346\,
            in1 => \N__8937\,
            in2 => \N__9628\,
            in3 => \N__8951\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__9947\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS10_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8924\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10140\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10\,
            ltout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8931\,
            in3 => \N__10015\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101010"
        )
    port map (
            in0 => \N__10016\,
            in1 => \_gnd_net_\,
            in2 => \N__8928\,
            in3 => \N__8883\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_RNI8MQ3_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8821\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8704\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10338\,
            in1 => \N__9576\,
            in2 => \_gnd_net_\,
            in3 => \N__9829\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__9306\,
            sr => \N__9962\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10411\,
            in1 => \N__10347\,
            in2 => \_gnd_net_\,
            in3 => \N__9828\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__9305\,
            sr => \N__9956\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10412\,
            in1 => \N__10342\,
            in2 => \_gnd_net_\,
            in3 => \N__10198\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__9291\,
            sr => \N__9950\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9472\,
            in1 => \N__10340\,
            in2 => \_gnd_net_\,
            in3 => \N__9515\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__9291\,
            sr => \N__9950\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9556\,
            in1 => \_gnd_net_\,
            in2 => \N__10357\,
            in3 => \N__9618\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__9291\,
            sr => \N__9950\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9768\,
            in1 => \N__10341\,
            in2 => \_gnd_net_\,
            in3 => \N__9516\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__9291\,
            sr => \N__9950\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__9473\,
            in1 => \_gnd_net_\,
            in2 => \N__9666\,
            in3 => \N__10339\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__9290\,
            sr => \N__9948\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9720\,
            in1 => \N__10303\,
            in2 => \_gnd_net_\,
            in3 => \N__9764\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__9292\,
            sr => \N__9946\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10304\,
            in1 => \N__9721\,
            in2 => \_gnd_net_\,
            in3 => \N__10188\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__9292\,
            sr => \N__9946\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10299\,
            in1 => \N__9575\,
            in2 => \_gnd_net_\,
            in3 => \N__9831\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10133\,
            ce => \N__10090\,
            sr => \N__9973\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10298\,
            in1 => \N__10413\,
            in2 => \_gnd_net_\,
            in3 => \N__9830\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10133\,
            ce => \N__10090\,
            sr => \N__9973\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10296\,
            in1 => \N__9723\,
            in2 => \_gnd_net_\,
            in3 => \N__9763\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10130\,
            ce => \N__10092\,
            sr => \N__9963\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9762\,
            in1 => \N__10295\,
            in2 => \_gnd_net_\,
            in3 => \N__9514\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10130\,
            ce => \N__10092\,
            sr => \N__9963\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10200\,
            in1 => \N__10353\,
            in2 => \_gnd_net_\,
            in3 => \N__9722\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10129\,
            ce => \N__10091\,
            sr => \N__9957\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9465\,
            in1 => \N__10294\,
            in2 => \_gnd_net_\,
            in3 => \N__9662\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10128\,
            ce => \N__10064\,
            sr => \N__9951\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10297\,
            in1 => \N__9630\,
            in2 => \_gnd_net_\,
            in3 => \N__9574\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10135\,
            ce => \N__10098\,
            sr => \N__9981\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10352\,
            in1 => \N__9508\,
            in2 => \_gnd_net_\,
            in3 => \N__9477\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10134\,
            ce => \N__10093\,
            sr => \N__9974\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10404\,
            in1 => \N__10351\,
            in2 => \_gnd_net_\,
            in3 => \N__10199\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10131\,
            ce => \N__10097\,
            sr => \N__9964\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 3 2024 18:22:34

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    A : in std_logic_vector(20 downto 0);
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    DRDDIR : out std_logic;
    DBDIR : in std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RAMENn : out std_logic;
    TSn : in std_logic;
    RASn : out std_logic;
    CLMBEn : out std_logic;
    RESETn : in std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    TACKn : out std_logic;
    CLKEN : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__7716\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_OUT_i_i\ : std_logic;
signal \N_620_i\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_5\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_15\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_4\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \CLK40_OUT_i_i\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_REG_SM.STATE_COUNT5\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \CLK40_OUT_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_45_0_0_en_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \U712_CYCLE_TERM.N_45_0_0_en_0\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \A_c_14\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1_0_cascade_\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \CLLBEn_c\ : std_logic;
signal \U712_REG_SM.N_160\ : std_logic;
signal \U712_CHIP_RAM.A_m_14\ : std_logic;
signal \A_c_7\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.A_m_10\ : std_logic;
signal \A_c_3\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_80_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_3_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_83\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_i_1\ : std_logic;
signal \U712_CHIP_RAM.N_110\ : std_logic;
signal \U712_CHIP_RAM.N_110_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_58\ : std_logic;
signal \U712_CHIP_RAM.N_58_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_118\ : std_logic;
signal \U712_CHIP_RAM.N_118_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_0_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_o2_0_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_40_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD14\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_10_u_0_1_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.N_40\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_1\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_6_tz\ : std_logic;
signal \U712_REG_SM.N_148_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_157_0\ : std_logic;
signal \U712_REG_SM.N_157_0_cascade_\ : std_logic;
signal \U712_REG_SM.REG_TACK_7_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_5\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_3_0_1\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_0\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_1\ : std_logic;
signal \U712_REG_SM.N_146_0_cascade_\ : std_logic;
signal \U712_REG_SM.DS_EN_0_sqmuxa_1\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA21_0_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_i_1\ : std_logic;
signal \U712_CHIP_RAM.N_116_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_117\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_67_i_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_26\ : std_logic;
signal \U712_CHIP_RAM.N_116\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_1_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_2_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.N_100\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_2\ : std_logic;
signal \U712_CHIP_RAM.N_87\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a5_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_a5_0_0_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_21_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_10_u_0_2_0\ : std_logic;
signal \U712_CHIP_RAM.N_13\ : std_logic;
signal \U712_CHIP_RAM.N_13_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_0_a2_0\ : std_logic;
signal \N_23_i\ : std_logic;
signal \CUMBEn_c\ : std_logic;
signal \U712_REG_SM.N_148_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_155_0_cascade_\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_145_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_145_0_cascade_\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \N_22_i\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA21_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_a5_0_1_3\ : std_logic;
signal \U712_CHIP_RAM.N_82\ : std_logic;
signal \U712_CHIP_RAM.N_105\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_ac0_1_out\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_ac0_1_out_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_ac0_3_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_ac0_3_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_36\ : std_logic;
signal \U712_CHIP_RAM.N_44\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_c6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_c4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_c6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER19_i_0_1_0\ : std_logic;
signal \U712_REG_SM.N_152_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_RNIVQBP4Z0Z_6\ : std_logic;
signal \U712_REG_SM.DS_EN_7_0\ : std_logic;
signal \U712_REG_SM.N_149_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_a3_0_0_3\ : std_logic;
signal \U712_REG_SM.N_156_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_155_0\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U712_REG_SM.LDS_OUT_2_0_0\ : std_logic;
signal \U712_REG_SM.LDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_LDSn_i\ : std_logic;
signal \U712_REG_SM.UDS_OUTZ0\ : std_logic;
signal \U712_REG_SM.DS_ENZ0\ : std_logic;
signal \U712_REG_SM_un1_UDSn_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \U712_REG_SM.N_182\ : std_logic;
signal \U712_REG_SM.N_146_0\ : std_logic;
signal \ASn_c\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \U712_REG_SM.N_177_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \DRDDIR_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \CLKEN_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    CLKEN <= \CLKEN_wire\;
    BANK1 <= \BANK1_wire\;
    CMA <= \CMA_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \TSn_wire\ <= TSn;
    UDSn <= \UDSn_wire\;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    LDSn <= \LDSn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_OUT_i\,
            REFERENCECLK => \N__2729\,
            RESETB => \N__6861\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_OUT\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7716\,
            DIN => \N__7715\,
            DOUT => \N__7714\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7716\,
            PADOUT => \N__7715\,
            PADIN => \N__7714\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6872\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7707\,
            DIN => \N__7706\,
            DOUT => \N__7705\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7707\,
            PADOUT => \N__7706\,
            PADIN => \N__7705\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7698\,
            DIN => \N__7697\,
            DOUT => \N__7696\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7698\,
            PADOUT => \N__7697\,
            PADIN => \N__7696\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6176\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7689\,
            DIN => \N__7688\,
            DOUT => \N__7687\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7689\,
            PADOUT => \N__7688\,
            PADIN => \N__7687\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6674\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7680\,
            DIN => \N__7679\,
            DOUT => \N__7678\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7680\,
            PADOUT => \N__7679\,
            PADIN => \N__7678\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKEN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7671\,
            DIN => \N__7670\,
            DOUT => \N__7669\,
            PACKAGEPIN => \CLKEN_wire\
        );

    \CLKEN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7671\,
            PADOUT => \N__7670\,
            PADIN => \N__7669\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6871\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7662\,
            DIN => \N__7661\,
            DOUT => \N__7660\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7662\,
            PADOUT => \N__7661\,
            PADIN => \N__7660\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7653\,
            DIN => \N__7652\,
            DOUT => \N__7651\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7653\,
            PADOUT => \N__7652\,
            PADIN => \N__7651\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7644\,
            DIN => \N__7643\,
            DOUT => \N__7642\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7644\,
            PADOUT => \N__7643\,
            PADIN => \N__7642\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7635\,
            DIN => \N__7634\,
            DOUT => \N__7633\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7635\,
            PADOUT => \N__7634\,
            PADIN => \N__7633\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3023\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7626\,
            DIN => \N__7625\,
            DOUT => \N__7624\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7626\,
            PADOUT => \N__7625\,
            PADIN => \N__7624\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3423\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7617\,
            DIN => \N__7616\,
            DOUT => \N__7615\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7617\,
            PADOUT => \N__7616\,
            PADIN => \N__7615\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRDENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7608\,
            DIN => \N__7607\,
            DOUT => \N__7606\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7608\,
            PADOUT => \N__7607\,
            PADIN => \N__7606\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4139\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7599\,
            DIN => \N__7598\,
            DOUT => \N__7597\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7599\,
            PADOUT => \N__7598\,
            PADIN => \N__7597\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7590\,
            DIN => \N__7589\,
            DOUT => \N__7588\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7590\,
            PADOUT => \N__7589\,
            PADIN => \N__7588\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3308\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7581\,
            DIN => \N__7580\,
            DOUT => \N__7579\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7581\,
            PADOUT => \N__7580\,
            PADIN => \N__7579\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7572\,
            DIN => \N__7571\,
            DOUT => \N__7570\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7572\,
            PADOUT => \N__7571\,
            PADIN => \N__7570\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7563\,
            DIN => \N__7562\,
            DOUT => \N__7561\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7563\,
            PADOUT => \N__7562\,
            PADIN => \N__7561\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2798\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7554\,
            DIN => \N__7553\,
            DOUT => \N__7552\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7554\,
            PADOUT => \N__7553\,
            PADIN => \N__7552\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7545\,
            DIN => \N__7544\,
            DOUT => \N__7543\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7545\,
            PADOUT => \N__7544\,
            PADIN => \N__7543\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6392\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7536\,
            DIN => \N__7535\,
            DOUT => \N__7534\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7536\,
            PADOUT => \N__7535\,
            PADIN => \N__7534\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7527\,
            DIN => \N__7526\,
            DOUT => \N__7525\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7527\,
            PADOUT => \N__7526\,
            PADIN => \N__7525\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7518\,
            DIN => \N__7517\,
            DOUT => \N__7516\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7518\,
            PADOUT => \N__7517\,
            PADIN => \N__7516\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3737\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7509\,
            DIN => \N__7508\,
            DOUT => \N__7507\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7509\,
            PADOUT => \N__7508\,
            PADIN => \N__7507\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7500\,
            DIN => \N__7499\,
            DOUT => \N__7498\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7500\,
            PADOUT => \N__7499\,
            PADIN => \N__7498\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6452\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7491\,
            DIN => \N__7490\,
            DOUT => \N__7489\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7491\,
            PADOUT => \N__7490\,
            PADIN => \N__7489\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7482\,
            DIN => \N__7481\,
            DOUT => \N__7480\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7482\,
            PADOUT => \N__7481\,
            PADIN => \N__7480\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7473\,
            DIN => \N__7472\,
            DOUT => \N__7471\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7473\,
            PADOUT => \N__7472\,
            PADIN => \N__7471\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7464\,
            DIN => \N__7463\,
            DOUT => \N__7462\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7464\,
            PADOUT => \N__7463\,
            PADIN => \N__7462\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7455\,
            DIN => \N__7454\,
            DOUT => \N__7453\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7455\,
            PADOUT => \N__7454\,
            PADIN => \N__7453\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7446\,
            DIN => \N__7445\,
            DOUT => \N__7444\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7446\,
            PADOUT => \N__7445\,
            PADIN => \N__7444\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3068\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7437\,
            DIN => \N__7436\,
            DOUT => \N__7435\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7437\,
            PADOUT => \N__7436\,
            PADIN => \N__7435\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7428\,
            DIN => \N__7427\,
            DOUT => \N__7426\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7428\,
            PADOUT => \N__7427\,
            PADIN => \N__7426\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7419\,
            DIN => \N__7418\,
            DOUT => \N__7417\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7419\,
            PADOUT => \N__7418\,
            PADIN => \N__7417\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7410\,
            DIN => \N__7409\,
            DOUT => \N__7408\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7410\,
            PADOUT => \N__7409\,
            PADIN => \N__7408\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2906\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7401\,
            DIN => \N__7400\,
            DOUT => \N__7399\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7401\,
            PADOUT => \N__7400\,
            PADIN => \N__7399\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6509\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7392\,
            DIN => \N__7391\,
            DOUT => \N__7390\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7392\,
            PADOUT => \N__7391\,
            PADIN => \N__7390\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7383\,
            DIN => \N__7382\,
            DOUT => \N__7381\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7383\,
            PADOUT => \N__7382\,
            PADIN => \N__7381\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6248\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7374\,
            DIN => \N__7373\,
            DOUT => \N__7372\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7374\,
            PADOUT => \N__7373\,
            PADIN => \N__7372\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7365\,
            DIN => \N__7364\,
            DOUT => \N__7363\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7365\,
            PADOUT => \N__7364\,
            PADIN => \N__7363\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7356\,
            DIN => \N__7355\,
            DOUT => \N__7354\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7356\,
            PADOUT => \N__7355\,
            PADIN => \N__7354\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2867\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7347\,
            DIN => \N__7346\,
            DOUT => \N__7345\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7347\,
            PADOUT => \N__7346\,
            PADIN => \N__7345\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6074\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7338\,
            DIN => \N__7337\,
            DOUT => \N__7336\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7338\,
            PADOUT => \N__7337\,
            PADIN => \N__7336\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2747\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7329\,
            DIN => \N__7328\,
            DOUT => \N__7327\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7329\,
            PADOUT => \N__7328\,
            PADIN => \N__7327\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7320\,
            DIN => \N__7319\,
            DOUT => \N__7318\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7320\,
            PADOUT => \N__7319\,
            PADIN => \N__7318\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7311\,
            DIN => \N__7310\,
            DOUT => \N__7309\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7311\,
            PADOUT => \N__7310\,
            PADIN => \N__7309\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4598\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7302\,
            DIN => \N__7301\,
            DOUT => \N__7300\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7302\,
            PADOUT => \N__7301\,
            PADIN => \N__7300\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7293\,
            DIN => \N__7292\,
            DOUT => \N__7291\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7293\,
            PADOUT => \N__7292\,
            PADIN => \N__7291\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2978\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7284\,
            DIN => \N__7283\,
            DOUT => \N__7282\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7284\,
            PADOUT => \N__7283\,
            PADIN => \N__7282\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6813\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7275\,
            DIN => \N__7274\,
            DOUT => \N__7273\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7275\,
            PADOUT => \N__7274\,
            PADIN => \N__7273\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3782\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7266\,
            DIN => \N__7265\,
            DOUT => \N__7264\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7266\,
            PADOUT => \N__7265\,
            PADIN => \N__7264\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4106\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7257\,
            DIN => \N__7256\,
            DOUT => \N__7255\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7257\,
            PADOUT => \N__7256\,
            PADIN => \N__7255\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6073\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7248\,
            DIN => \N__7247\,
            DOUT => \N__7246\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7248\,
            PADOUT => \N__7247\,
            PADIN => \N__7246\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7239\,
            DIN => \N__7238\,
            DOUT => \N__7237\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7239\,
            PADOUT => \N__7238\,
            PADIN => \N__7237\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7230\,
            DIN => \N__7229\,
            DOUT => \N__7228\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7230\,
            PADOUT => \N__7229\,
            PADIN => \N__7228\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4769\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7221\,
            DIN => \N__7220\,
            DOUT => \N__7219\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7221\,
            PADOUT => \N__7220\,
            PADIN => \N__7219\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4745\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7212\,
            DIN => \N__7211\,
            DOUT => \N__7210\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7212\,
            PADOUT => \N__7211\,
            PADIN => \N__7210\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4436\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7203\,
            DIN => \N__7202\,
            DOUT => \N__7201\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7203\,
            PADOUT => \N__7202\,
            PADIN => \N__7201\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7194\,
            DIN => \N__7193\,
            DOUT => \N__7192\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7194\,
            PADOUT => \N__7193\,
            PADIN => \N__7192\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7185\,
            DIN => \N__7184\,
            DOUT => \N__7183\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7185\,
            PADOUT => \N__7184\,
            PADIN => \N__7183\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7176\,
            DIN => \N__7175\,
            DOUT => \N__7174\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7176\,
            PADOUT => \N__7175\,
            PADIN => \N__7174\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3692\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7167\,
            DIN => \N__7166\,
            DOUT => \N__7165\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7167\,
            PADOUT => \N__7166\,
            PADIN => \N__7165\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7158\,
            DIN => \N__7157\,
            DOUT => \N__7156\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7158\,
            PADOUT => \N__7157\,
            PADIN => \N__7156\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4460\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7149\,
            DIN => \N__7148\,
            DOUT => \N__7147\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7149\,
            PADOUT => \N__7148\,
            PADIN => \N__7147\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2852\,
            DIN0 => OPEN,
            DOUT0 => \N__2894\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7140\,
            DIN => \N__7139\,
            DOUT => \N__7138\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7140\,
            PADOUT => \N__7139\,
            PADIN => \N__7138\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2927\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1701\ : InMux
    port map (
            O => \N__7121\,
            I => \N__7110\
        );

    \I__1700\ : InMux
    port map (
            O => \N__7120\,
            I => \N__7107\
        );

    \I__1699\ : InMux
    port map (
            O => \N__7119\,
            I => \N__7104\
        );

    \I__1698\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7099\
        );

    \I__1697\ : InMux
    port map (
            O => \N__7117\,
            I => \N__7099\
        );

    \I__1696\ : InMux
    port map (
            O => \N__7116\,
            I => \N__7092\
        );

    \I__1695\ : InMux
    port map (
            O => \N__7115\,
            I => \N__7092\
        );

    \I__1694\ : InMux
    port map (
            O => \N__7114\,
            I => \N__7092\
        );

    \I__1693\ : InMux
    port map (
            O => \N__7113\,
            I => \N__7089\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__7110\,
            I => \N__7074\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__7107\,
            I => \N__7063\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__7104\,
            I => \N__7060\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__7099\,
            I => \N__7056\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__7092\,
            I => \N__7052\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__7089\,
            I => \N__7047\
        );

    \I__1686\ : SRMux
    port map (
            O => \N__7088\,
            I => \N__6977\
        );

    \I__1685\ : SRMux
    port map (
            O => \N__7087\,
            I => \N__6977\
        );

    \I__1684\ : SRMux
    port map (
            O => \N__7086\,
            I => \N__6977\
        );

    \I__1683\ : SRMux
    port map (
            O => \N__7085\,
            I => \N__6977\
        );

    \I__1682\ : SRMux
    port map (
            O => \N__7084\,
            I => \N__6977\
        );

    \I__1681\ : SRMux
    port map (
            O => \N__7083\,
            I => \N__6977\
        );

    \I__1680\ : SRMux
    port map (
            O => \N__7082\,
            I => \N__6977\
        );

    \I__1679\ : SRMux
    port map (
            O => \N__7081\,
            I => \N__6977\
        );

    \I__1678\ : SRMux
    port map (
            O => \N__7080\,
            I => \N__6977\
        );

    \I__1677\ : SRMux
    port map (
            O => \N__7079\,
            I => \N__6977\
        );

    \I__1676\ : SRMux
    port map (
            O => \N__7078\,
            I => \N__6977\
        );

    \I__1675\ : SRMux
    port map (
            O => \N__7077\,
            I => \N__6977\
        );

    \I__1674\ : Glb2LocalMux
    port map (
            O => \N__7074\,
            I => \N__6977\
        );

    \I__1673\ : SRMux
    port map (
            O => \N__7073\,
            I => \N__6977\
        );

    \I__1672\ : SRMux
    port map (
            O => \N__7072\,
            I => \N__6977\
        );

    \I__1671\ : SRMux
    port map (
            O => \N__7071\,
            I => \N__6977\
        );

    \I__1670\ : SRMux
    port map (
            O => \N__7070\,
            I => \N__6977\
        );

    \I__1669\ : SRMux
    port map (
            O => \N__7069\,
            I => \N__6977\
        );

    \I__1668\ : SRMux
    port map (
            O => \N__7068\,
            I => \N__6977\
        );

    \I__1667\ : SRMux
    port map (
            O => \N__7067\,
            I => \N__6977\
        );

    \I__1666\ : SRMux
    port map (
            O => \N__7066\,
            I => \N__6977\
        );

    \I__1665\ : Glb2LocalMux
    port map (
            O => \N__7063\,
            I => \N__6977\
        );

    \I__1664\ : Glb2LocalMux
    port map (
            O => \N__7060\,
            I => \N__6977\
        );

    \I__1663\ : SRMux
    port map (
            O => \N__7059\,
            I => \N__6977\
        );

    \I__1662\ : Glb2LocalMux
    port map (
            O => \N__7056\,
            I => \N__6977\
        );

    \I__1661\ : SRMux
    port map (
            O => \N__7055\,
            I => \N__6977\
        );

    \I__1660\ : Glb2LocalMux
    port map (
            O => \N__7052\,
            I => \N__6977\
        );

    \I__1659\ : SRMux
    port map (
            O => \N__7051\,
            I => \N__6977\
        );

    \I__1658\ : SRMux
    port map (
            O => \N__7050\,
            I => \N__6977\
        );

    \I__1657\ : Glb2LocalMux
    port map (
            O => \N__7047\,
            I => \N__6977\
        );

    \I__1656\ : SRMux
    port map (
            O => \N__7046\,
            I => \N__6977\
        );

    \I__1655\ : SRMux
    port map (
            O => \N__7045\,
            I => \N__6977\
        );

    \I__1654\ : SRMux
    port map (
            O => \N__7044\,
            I => \N__6977\
        );

    \I__1653\ : GlobalMux
    port map (
            O => \N__6977\,
            I => \N__6974\
        );

    \I__1652\ : gio2CtrlBuf
    port map (
            O => \N__6974\,
            I => \RESETn_c_i_g\
        );

    \I__1651\ : InMux
    port map (
            O => \N__6971\,
            I => \N__6963\
        );

    \I__1650\ : InMux
    port map (
            O => \N__6970\,
            I => \N__6960\
        );

    \I__1649\ : InMux
    port map (
            O => \N__6969\,
            I => \N__6951\
        );

    \I__1648\ : InMux
    port map (
            O => \N__6968\,
            I => \N__6951\
        );

    \I__1647\ : InMux
    port map (
            O => \N__6967\,
            I => \N__6951\
        );

    \I__1646\ : InMux
    port map (
            O => \N__6966\,
            I => \N__6948\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__6963\,
            I => \N__6942\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__6960\,
            I => \N__6942\
        );

    \I__1643\ : InMux
    port map (
            O => \N__6959\,
            I => \N__6939\
        );

    \I__1642\ : InMux
    port map (
            O => \N__6958\,
            I => \N__6936\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__6951\,
            I => \N__6933\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__6948\,
            I => \N__6930\
        );

    \I__1639\ : InMux
    port map (
            O => \N__6947\,
            I => \N__6927\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__6942\,
            I => \N__6924\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__6939\,
            I => \N__6921\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__6936\,
            I => \N__6918\
        );

    \I__1635\ : Span4Mux_v
    port map (
            O => \N__6933\,
            I => \N__6913\
        );

    \I__1634\ : Span4Mux_v
    port map (
            O => \N__6930\,
            I => \N__6913\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__6927\,
            I => \N__6910\
        );

    \I__1632\ : Span4Mux_h
    port map (
            O => \N__6924\,
            I => \N__6903\
        );

    \I__1631\ : Span4Mux_v
    port map (
            O => \N__6921\,
            I => \N__6903\
        );

    \I__1630\ : Span4Mux_v
    port map (
            O => \N__6918\,
            I => \N__6903\
        );

    \I__1629\ : Sp12to4
    port map (
            O => \N__6913\,
            I => \N__6900\
        );

    \I__1628\ : Span12Mux_v
    port map (
            O => \N__6910\,
            I => \N__6895\
        );

    \I__1627\ : Sp12to4
    port map (
            O => \N__6903\,
            I => \N__6895\
        );

    \I__1626\ : Span12Mux_h
    port map (
            O => \N__6900\,
            I => \N__6892\
        );

    \I__1625\ : Span12Mux_h
    port map (
            O => \N__6895\,
            I => \N__6889\
        );

    \I__1624\ : Odrv12
    port map (
            O => \N__6892\,
            I => \RESETn_c\
        );

    \I__1623\ : Odrv12
    port map (
            O => \N__6889\,
            I => \RESETn_c\
        );

    \I__1622\ : IoInMux
    port map (
            O => \N__6884\,
            I => \N__6881\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__6881\,
            I => \N__6878\
        );

    \I__1620\ : Span12Mux_s7_v
    port map (
            O => \N__6878\,
            I => \N__6875\
        );

    \I__1619\ : Odrv12
    port map (
            O => \N__6875\,
            I => \RESETn_c_i\
        );

    \I__1618\ : IoInMux
    port map (
            O => \N__6872\,
            I => \N__6868\
        );

    \I__1617\ : IoInMux
    port map (
            O => \N__6871\,
            I => \N__6865\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__6868\,
            I => \N__6862\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__6865\,
            I => \N__6858\
        );

    \I__1614\ : Span4Mux_s3_v
    port map (
            O => \N__6862\,
            I => \N__6855\
        );

    \I__1613\ : IoInMux
    port map (
            O => \N__6861\,
            I => \N__6852\
        );

    \I__1612\ : IoSpan4Mux
    port map (
            O => \N__6858\,
            I => \N__6849\
        );

    \I__1611\ : Span4Mux_v
    port map (
            O => \N__6855\,
            I => \N__6846\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__6852\,
            I => \N__6843\
        );

    \I__1609\ : Sp12to4
    port map (
            O => \N__6849\,
            I => \N__6840\
        );

    \I__1608\ : Span4Mux_h
    port map (
            O => \N__6846\,
            I => \N__6837\
        );

    \I__1607\ : Span4Mux_s3_v
    port map (
            O => \N__6843\,
            I => \N__6834\
        );

    \I__1606\ : Span12Mux_s7_h
    port map (
            O => \N__6840\,
            I => \N__6831\
        );

    \I__1605\ : Span4Mux_h
    port map (
            O => \N__6837\,
            I => \N__6826\
        );

    \I__1604\ : Span4Mux_v
    port map (
            O => \N__6834\,
            I => \N__6826\
        );

    \I__1603\ : Odrv12
    port map (
            O => \N__6831\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1602\ : Odrv4
    port map (
            O => \N__6826\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__6821\,
            I => \N__6817\
        );

    \I__1600\ : InMux
    port map (
            O => \N__6820\,
            I => \N__6814\
        );

    \I__1599\ : InMux
    port map (
            O => \N__6817\,
            I => \N__6810\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__6814\,
            I => \N__6806\
        );

    \I__1597\ : IoInMux
    port map (
            O => \N__6813\,
            I => \N__6803\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__6810\,
            I => \N__6800\
        );

    \I__1595\ : InMux
    port map (
            O => \N__6809\,
            I => \N__6797\
        );

    \I__1594\ : Span4Mux_v
    port map (
            O => \N__6806\,
            I => \N__6794\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__6803\,
            I => \N__6791\
        );

    \I__1592\ : Span4Mux_h
    port map (
            O => \N__6800\,
            I => \N__6786\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__6797\,
            I => \N__6786\
        );

    \I__1590\ : Span4Mux_h
    port map (
            O => \N__6794\,
            I => \N__6783\
        );

    \I__1589\ : Span12Mux_s9_v
    port map (
            O => \N__6791\,
            I => \N__6780\
        );

    \I__1588\ : Span4Mux_v
    port map (
            O => \N__6786\,
            I => \N__6777\
        );

    \I__1587\ : Span4Mux_v
    port map (
            O => \N__6783\,
            I => \N__6774\
        );

    \I__1586\ : Span12Mux_v
    port map (
            O => \N__6780\,
            I => \N__6770\
        );

    \I__1585\ : Span4Mux_h
    port map (
            O => \N__6777\,
            I => \N__6767\
        );

    \I__1584\ : Sp12to4
    port map (
            O => \N__6774\,
            I => \N__6764\
        );

    \I__1583\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6761\
        );

    \I__1582\ : Span12Mux_h
    port map (
            O => \N__6770\,
            I => \N__6758\
        );

    \I__1581\ : Sp12to4
    port map (
            O => \N__6767\,
            I => \N__6755\
        );

    \I__1580\ : Span12Mux_v
    port map (
            O => \N__6764\,
            I => \N__6750\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__6761\,
            I => \N__6750\
        );

    \I__1578\ : Span12Mux_h
    port map (
            O => \N__6758\,
            I => \N__6747\
        );

    \I__1577\ : Span12Mux_v
    port map (
            O => \N__6755\,
            I => \N__6742\
        );

    \I__1576\ : Span12Mux_h
    port map (
            O => \N__6750\,
            I => \N__6742\
        );

    \I__1575\ : Odrv12
    port map (
            O => \N__6747\,
            I => \DRDENn_c\
        );

    \I__1574\ : Odrv12
    port map (
            O => \N__6742\,
            I => \DRDENn_c\
        );

    \I__1573\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6733\
        );

    \I__1572\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6730\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__6733\,
            I => \N__6727\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__6730\,
            I => \N__6724\
        );

    \I__1569\ : Span4Mux_v
    port map (
            O => \N__6727\,
            I => \N__6719\
        );

    \I__1568\ : Span4Mux_v
    port map (
            O => \N__6724\,
            I => \N__6715\
        );

    \I__1567\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6712\
        );

    \I__1566\ : InMux
    port map (
            O => \N__6722\,
            I => \N__6709\
        );

    \I__1565\ : Span4Mux_v
    port map (
            O => \N__6719\,
            I => \N__6706\
        );

    \I__1564\ : InMux
    port map (
            O => \N__6718\,
            I => \N__6703\
        );

    \I__1563\ : Sp12to4
    port map (
            O => \N__6715\,
            I => \N__6696\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__6712\,
            I => \N__6696\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__6709\,
            I => \N__6696\
        );

    \I__1560\ : Sp12to4
    port map (
            O => \N__6706\,
            I => \N__6693\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__6703\,
            I => \N__6690\
        );

    \I__1558\ : Span12Mux_h
    port map (
            O => \N__6696\,
            I => \N__6687\
        );

    \I__1557\ : Span12Mux_h
    port map (
            O => \N__6693\,
            I => \N__6682\
        );

    \I__1556\ : Span12Mux_v
    port map (
            O => \N__6690\,
            I => \N__6682\
        );

    \I__1555\ : Span12Mux_v
    port map (
            O => \N__6687\,
            I => \N__6677\
        );

    \I__1554\ : Span12Mux_h
    port map (
            O => \N__6682\,
            I => \N__6677\
        );

    \I__1553\ : Odrv12
    port map (
            O => \N__6677\,
            I => \RnW_c\
        );

    \I__1552\ : IoInMux
    port map (
            O => \N__6674\,
            I => \N__6671\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__6671\,
            I => \N__6668\
        );

    \I__1550\ : IoSpan4Mux
    port map (
            O => \N__6668\,
            I => \N__6665\
        );

    \I__1549\ : Sp12to4
    port map (
            O => \N__6665\,
            I => \N__6662\
        );

    \I__1548\ : Span12Mux_s9_h
    port map (
            O => \N__6662\,
            I => \N__6659\
        );

    \I__1547\ : Odrv12
    port map (
            O => \N__6659\,
            I => \DRDDIR_c\
        );

    \I__1546\ : InMux
    port map (
            O => \N__6656\,
            I => \N__6650\
        );

    \I__1545\ : InMux
    port map (
            O => \N__6655\,
            I => \N__6643\
        );

    \I__1544\ : InMux
    port map (
            O => \N__6654\,
            I => \N__6643\
        );

    \I__1543\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6643\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__6650\,
            I => \N__6640\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__6643\,
            I => \U712_REG_SM.N_155_0\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__6640\,
            I => \U712_REG_SM.N_155_0\
        );

    \I__1539\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6626\
        );

    \I__1538\ : InMux
    port map (
            O => \N__6634\,
            I => \N__6626\
        );

    \I__1537\ : InMux
    port map (
            O => \N__6633\,
            I => \N__6621\
        );

    \I__1536\ : InMux
    port map (
            O => \N__6632\,
            I => \N__6621\
        );

    \I__1535\ : InMux
    port map (
            O => \N__6631\,
            I => \N__6618\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__6626\,
            I => \N__6615\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__6621\,
            I => \N__6610\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__6618\,
            I => \N__6610\
        );

    \I__1531\ : Span4Mux_v
    port map (
            O => \N__6615\,
            I => \N__6604\
        );

    \I__1530\ : Span4Mux_v
    port map (
            O => \N__6610\,
            I => \N__6604\
        );

    \I__1529\ : InMux
    port map (
            O => \N__6609\,
            I => \N__6601\
        );

    \I__1528\ : Span4Mux_h
    port map (
            O => \N__6604\,
            I => \N__6598\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__6601\,
            I => \N__6595\
        );

    \I__1526\ : Sp12to4
    port map (
            O => \N__6598\,
            I => \N__6590\
        );

    \I__1525\ : Span12Mux_v
    port map (
            O => \N__6595\,
            I => \N__6590\
        );

    \I__1524\ : Odrv12
    port map (
            O => \N__6590\,
            I => \A_c_0\
        );

    \I__1523\ : CascadeMux
    port map (
            O => \N__6587\,
            I => \N__6583\
        );

    \I__1522\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6576\
        );

    \I__1521\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6576\
        );

    \I__1520\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6573\
        );

    \I__1519\ : InMux
    port map (
            O => \N__6581\,
            I => \N__6570\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__6576\,
            I => \N__6563\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__6573\,
            I => \N__6563\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__6570\,
            I => \N__6563\
        );

    \I__1515\ : Span4Mux_v
    port map (
            O => \N__6563\,
            I => \N__6560\
        );

    \I__1514\ : Sp12to4
    port map (
            O => \N__6560\,
            I => \N__6556\
        );

    \I__1513\ : InMux
    port map (
            O => \N__6559\,
            I => \N__6553\
        );

    \I__1512\ : Span12Mux_h
    port map (
            O => \N__6556\,
            I => \N__6550\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__6553\,
            I => \N__6547\
        );

    \I__1510\ : Span12Mux_v
    port map (
            O => \N__6550\,
            I => \N__6544\
        );

    \I__1509\ : Span12Mux_v
    port map (
            O => \N__6547\,
            I => \N__6541\
        );

    \I__1508\ : Odrv12
    port map (
            O => \N__6544\,
            I => \SIZ_c_0\
        );

    \I__1507\ : Odrv12
    port map (
            O => \N__6541\,
            I => \SIZ_c_0\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__6536\,
            I => \N__6532\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__6535\,
            I => \N__6529\
        );

    \I__1504\ : InMux
    port map (
            O => \N__6532\,
            I => \N__6524\
        );

    \I__1503\ : InMux
    port map (
            O => \N__6529\,
            I => \N__6524\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__6524\,
            I => \U712_REG_SM.LDS_OUT_2_0_0\
        );

    \I__1501\ : InMux
    port map (
            O => \N__6521\,
            I => \N__6517\
        );

    \I__1500\ : InMux
    port map (
            O => \N__6520\,
            I => \N__6514\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__6517\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__6514\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__1497\ : IoInMux
    port map (
            O => \N__6509\,
            I => \N__6506\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__6506\,
            I => \N__6503\
        );

    \I__1495\ : IoSpan4Mux
    port map (
            O => \N__6503\,
            I => \N__6500\
        );

    \I__1494\ : Span4Mux_s2_v
    port map (
            O => \N__6500\,
            I => \N__6497\
        );

    \I__1493\ : Sp12to4
    port map (
            O => \N__6497\,
            I => \N__6494\
        );

    \I__1492\ : Span12Mux_h
    port map (
            O => \N__6494\,
            I => \N__6491\
        );

    \I__1491\ : Odrv12
    port map (
            O => \N__6491\,
            I => \U712_REG_SM_un1_LDSn_i\
        );

    \I__1490\ : InMux
    port map (
            O => \N__6488\,
            I => \N__6485\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__6485\,
            I => \N__6481\
        );

    \I__1488\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6478\
        );

    \I__1487\ : Odrv4
    port map (
            O => \N__6481\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__6478\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__1485\ : InMux
    port map (
            O => \N__6473\,
            I => \N__6470\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__6470\,
            I => \N__6465\
        );

    \I__1483\ : InMux
    port map (
            O => \N__6469\,
            I => \N__6462\
        );

    \I__1482\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6459\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__6465\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__6462\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__6459\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1478\ : IoInMux
    port map (
            O => \N__6452\,
            I => \N__6449\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__6449\,
            I => \N__6446\
        );

    \I__1476\ : Span12Mux_s2_v
    port map (
            O => \N__6446\,
            I => \N__6443\
        );

    \I__1475\ : Span12Mux_h
    port map (
            O => \N__6443\,
            I => \N__6440\
        );

    \I__1474\ : Odrv12
    port map (
            O => \N__6440\,
            I => \U712_REG_SM_un1_UDSn_i\
        );

    \I__1473\ : InMux
    port map (
            O => \N__6437\,
            I => \N__6433\
        );

    \I__1472\ : InMux
    port map (
            O => \N__6436\,
            I => \N__6430\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__6433\,
            I => \N__6427\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__6430\,
            I => \N__6424\
        );

    \I__1469\ : Span4Mux_h
    port map (
            O => \N__6427\,
            I => \N__6421\
        );

    \I__1468\ : Span4Mux_h
    port map (
            O => \N__6424\,
            I => \N__6415\
        );

    \I__1467\ : Span4Mux_v
    port map (
            O => \N__6421\,
            I => \N__6415\
        );

    \I__1466\ : InMux
    port map (
            O => \N__6420\,
            I => \N__6410\
        );

    \I__1465\ : Span4Mux_v
    port map (
            O => \N__6415\,
            I => \N__6407\
        );

    \I__1464\ : InMux
    port map (
            O => \N__6414\,
            I => \N__6404\
        );

    \I__1463\ : InMux
    port map (
            O => \N__6413\,
            I => \N__6401\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__6410\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1461\ : Odrv4
    port map (
            O => \N__6407\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__6404\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__6401\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1458\ : IoInMux
    port map (
            O => \N__6392\,
            I => \N__6389\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__6389\,
            I => \N__6386\
        );

    \I__1456\ : Span12Mux_s7_v
    port map (
            O => \N__6386\,
            I => \N__6383\
        );

    \I__1455\ : Odrv12
    port map (
            O => \N__6383\,
            I => \CRCSn_c\
        );

    \I__1454\ : InMux
    port map (
            O => \N__6380\,
            I => \N__6371\
        );

    \I__1453\ : InMux
    port map (
            O => \N__6379\,
            I => \N__6366\
        );

    \I__1452\ : InMux
    port map (
            O => \N__6378\,
            I => \N__6366\
        );

    \I__1451\ : InMux
    port map (
            O => \N__6377\,
            I => \N__6359\
        );

    \I__1450\ : InMux
    port map (
            O => \N__6376\,
            I => \N__6355\
        );

    \I__1449\ : InMux
    port map (
            O => \N__6375\,
            I => \N__6350\
        );

    \I__1448\ : InMux
    port map (
            O => \N__6374\,
            I => \N__6350\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__6371\,
            I => \N__6347\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__6366\,
            I => \N__6344\
        );

    \I__1445\ : CascadeMux
    port map (
            O => \N__6365\,
            I => \N__6341\
        );

    \I__1444\ : InMux
    port map (
            O => \N__6364\,
            I => \N__6338\
        );

    \I__1443\ : InMux
    port map (
            O => \N__6363\,
            I => \N__6335\
        );

    \I__1442\ : InMux
    port map (
            O => \N__6362\,
            I => \N__6332\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__6359\,
            I => \N__6329\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__6358\,
            I => \N__6324\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__6355\,
            I => \N__6319\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__6350\,
            I => \N__6319\
        );

    \I__1437\ : Span4Mux_h
    port map (
            O => \N__6347\,
            I => \N__6313\
        );

    \I__1436\ : Span4Mux_h
    port map (
            O => \N__6344\,
            I => \N__6313\
        );

    \I__1435\ : InMux
    port map (
            O => \N__6341\,
            I => \N__6310\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__6338\,
            I => \N__6307\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__6335\,
            I => \N__6300\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__6332\,
            I => \N__6300\
        );

    \I__1431\ : Span4Mux_v
    port map (
            O => \N__6329\,
            I => \N__6300\
        );

    \I__1430\ : InMux
    port map (
            O => \N__6328\,
            I => \N__6297\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__6327\,
            I => \N__6293\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6324\,
            I => \N__6289\
        );

    \I__1427\ : Span4Mux_h
    port map (
            O => \N__6319\,
            I => \N__6286\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6318\,
            I => \N__6283\
        );

    \I__1425\ : Span4Mux_v
    port map (
            O => \N__6313\,
            I => \N__6280\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__6310\,
            I => \N__6271\
        );

    \I__1423\ : Span4Mux_h
    port map (
            O => \N__6307\,
            I => \N__6271\
        );

    \I__1422\ : Span4Mux_h
    port map (
            O => \N__6300\,
            I => \N__6271\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__6297\,
            I => \N__6271\
        );

    \I__1420\ : InMux
    port map (
            O => \N__6296\,
            I => \N__6268\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6263\
        );

    \I__1418\ : InMux
    port map (
            O => \N__6292\,
            I => \N__6263\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__6289\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1416\ : Odrv4
    port map (
            O => \N__6286\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__6283\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__6280\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__6271\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6268\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6263\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1410\ : IoInMux
    port map (
            O => \N__6248\,
            I => \N__6245\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__6245\,
            I => \N__6242\
        );

    \I__1408\ : Span4Mux_s2_v
    port map (
            O => \N__6242\,
            I => \N__6239\
        );

    \I__1407\ : Span4Mux_v
    port map (
            O => \N__6239\,
            I => \N__6236\
        );

    \I__1406\ : Span4Mux_v
    port map (
            O => \N__6236\,
            I => \N__6233\
        );

    \I__1405\ : Sp12to4
    port map (
            O => \N__6233\,
            I => \N__6230\
        );

    \I__1404\ : Odrv12
    port map (
            O => \N__6230\,
            I => \RASn_c\
        );

    \I__1403\ : InMux
    port map (
            O => \N__6227\,
            I => \N__6221\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6226\,
            I => \N__6218\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6213\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6224\,
            I => \N__6210\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__6221\,
            I => \N__6205\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6218\,
            I => \N__6205\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__6217\,
            I => \N__6201\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6216\,
            I => \N__6198\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__6213\,
            I => \N__6191\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6210\,
            I => \N__6191\
        );

    \I__1393\ : Span4Mux_h
    port map (
            O => \N__6205\,
            I => \N__6191\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6188\
        );

    \I__1391\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6185\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6198\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1389\ : Odrv4
    port map (
            O => \N__6191\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__6188\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__6185\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1386\ : IoInMux
    port map (
            O => \N__6176\,
            I => \N__6173\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__6173\,
            I => \N__6170\
        );

    \I__1384\ : Span12Mux_s5_v
    port map (
            O => \N__6170\,
            I => \N__6167\
        );

    \I__1383\ : Span12Mux_h
    port map (
            O => \N__6167\,
            I => \N__6164\
        );

    \I__1382\ : Odrv12
    port map (
            O => \N__6164\,
            I => \CASn_c\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__6161\,
            I => \N__6157\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6160\,
            I => \N__6153\
        );

    \I__1379\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6146\
        );

    \I__1378\ : InMux
    port map (
            O => \N__6156\,
            I => \N__6146\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__6153\,
            I => \N__6143\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6152\,
            I => \N__6140\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6151\,
            I => \N__6137\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__6146\,
            I => \N__6130\
        );

    \I__1373\ : Span4Mux_h
    port map (
            O => \N__6143\,
            I => \N__6130\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__6140\,
            I => \N__6130\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__6137\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__1370\ : Odrv4
    port map (
            O => \N__6130\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6125\,
            I => \N__6122\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__6122\,
            I => \N__6118\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6121\,
            I => \N__6115\
        );

    \I__1366\ : Span4Mux_h
    port map (
            O => \N__6118\,
            I => \N__6108\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__6115\,
            I => \N__6108\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6114\,
            I => \N__6105\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6113\,
            I => \N__6102\
        );

    \I__1362\ : Odrv4
    port map (
            O => \N__6108\,
            I => \U712_REG_SM.N_182\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6105\,
            I => \U712_REG_SM.N_182\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__6102\,
            I => \U712_REG_SM.N_182\
        );

    \I__1359\ : InMux
    port map (
            O => \N__6095\,
            I => \N__6092\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__6092\,
            I => \N__6087\
        );

    \I__1357\ : InMux
    port map (
            O => \N__6091\,
            I => \N__6084\
        );

    \I__1356\ : InMux
    port map (
            O => \N__6090\,
            I => \N__6081\
        );

    \I__1355\ : Odrv12
    port map (
            O => \N__6087\,
            I => \U712_REG_SM.N_146_0\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6084\,
            I => \U712_REG_SM.N_146_0\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__6081\,
            I => \U712_REG_SM.N_146_0\
        );

    \I__1352\ : IoInMux
    port map (
            O => \N__6074\,
            I => \N__6070\
        );

    \I__1351\ : IoInMux
    port map (
            O => \N__6073\,
            I => \N__6067\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6070\,
            I => \N__6064\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6067\,
            I => \N__6061\
        );

    \I__1348\ : Span4Mux_s1_v
    port map (
            O => \N__6064\,
            I => \N__6058\
        );

    \I__1347\ : Span4Mux_s1_v
    port map (
            O => \N__6061\,
            I => \N__6055\
        );

    \I__1346\ : Sp12to4
    port map (
            O => \N__6058\,
            I => \N__6052\
        );

    \I__1345\ : Sp12to4
    port map (
            O => \N__6055\,
            I => \N__6049\
        );

    \I__1344\ : Span12Mux_h
    port map (
            O => \N__6052\,
            I => \N__6044\
        );

    \I__1343\ : Span12Mux_h
    port map (
            O => \N__6049\,
            I => \N__6044\
        );

    \I__1342\ : Span12Mux_v
    port map (
            O => \N__6044\,
            I => \N__6041\
        );

    \I__1341\ : Odrv12
    port map (
            O => \N__6041\,
            I => \ASn_c\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6035\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__6035\,
            I => \N__6008\
        );

    \I__1338\ : ClkMux
    port map (
            O => \N__6034\,
            I => \N__5933\
        );

    \I__1337\ : ClkMux
    port map (
            O => \N__6033\,
            I => \N__5933\
        );

    \I__1336\ : ClkMux
    port map (
            O => \N__6032\,
            I => \N__5933\
        );

    \I__1335\ : ClkMux
    port map (
            O => \N__6031\,
            I => \N__5933\
        );

    \I__1334\ : ClkMux
    port map (
            O => \N__6030\,
            I => \N__5933\
        );

    \I__1333\ : ClkMux
    port map (
            O => \N__6029\,
            I => \N__5933\
        );

    \I__1332\ : ClkMux
    port map (
            O => \N__6028\,
            I => \N__5933\
        );

    \I__1331\ : ClkMux
    port map (
            O => \N__6027\,
            I => \N__5933\
        );

    \I__1330\ : ClkMux
    port map (
            O => \N__6026\,
            I => \N__5933\
        );

    \I__1329\ : ClkMux
    port map (
            O => \N__6025\,
            I => \N__5933\
        );

    \I__1328\ : ClkMux
    port map (
            O => \N__6024\,
            I => \N__5933\
        );

    \I__1327\ : ClkMux
    port map (
            O => \N__6023\,
            I => \N__5933\
        );

    \I__1326\ : ClkMux
    port map (
            O => \N__6022\,
            I => \N__5933\
        );

    \I__1325\ : ClkMux
    port map (
            O => \N__6021\,
            I => \N__5933\
        );

    \I__1324\ : ClkMux
    port map (
            O => \N__6020\,
            I => \N__5933\
        );

    \I__1323\ : ClkMux
    port map (
            O => \N__6019\,
            I => \N__5933\
        );

    \I__1322\ : ClkMux
    port map (
            O => \N__6018\,
            I => \N__5933\
        );

    \I__1321\ : ClkMux
    port map (
            O => \N__6017\,
            I => \N__5933\
        );

    \I__1320\ : ClkMux
    port map (
            O => \N__6016\,
            I => \N__5933\
        );

    \I__1319\ : ClkMux
    port map (
            O => \N__6015\,
            I => \N__5933\
        );

    \I__1318\ : ClkMux
    port map (
            O => \N__6014\,
            I => \N__5933\
        );

    \I__1317\ : ClkMux
    port map (
            O => \N__6013\,
            I => \N__5933\
        );

    \I__1316\ : ClkMux
    port map (
            O => \N__6012\,
            I => \N__5933\
        );

    \I__1315\ : ClkMux
    port map (
            O => \N__6011\,
            I => \N__5933\
        );

    \I__1314\ : Glb2LocalMux
    port map (
            O => \N__6008\,
            I => \N__5933\
        );

    \I__1313\ : ClkMux
    port map (
            O => \N__6007\,
            I => \N__5933\
        );

    \I__1312\ : ClkMux
    port map (
            O => \N__6006\,
            I => \N__5933\
        );

    \I__1311\ : ClkMux
    port map (
            O => \N__6005\,
            I => \N__5933\
        );

    \I__1310\ : ClkMux
    port map (
            O => \N__6004\,
            I => \N__5933\
        );

    \I__1309\ : ClkMux
    port map (
            O => \N__6003\,
            I => \N__5933\
        );

    \I__1308\ : ClkMux
    port map (
            O => \N__6002\,
            I => \N__5933\
        );

    \I__1307\ : ClkMux
    port map (
            O => \N__6001\,
            I => \N__5933\
        );

    \I__1306\ : ClkMux
    port map (
            O => \N__6000\,
            I => \N__5933\
        );

    \I__1305\ : GlobalMux
    port map (
            O => \N__5933\,
            I => \CLK80_OUT\
        );

    \I__1304\ : CEMux
    port map (
            O => \N__5930\,
            I => \N__5927\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__5927\,
            I => \U712_REG_SM.N_177_0\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__5924\,
            I => \N__5921\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5921\,
            I => \N__5918\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__5918\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_c6\
        );

    \I__1299\ : InMux
    port map (
            O => \N__5915\,
            I => \N__5908\
        );

    \I__1298\ : InMux
    port map (
            O => \N__5914\,
            I => \N__5908\
        );

    \I__1297\ : InMux
    port map (
            O => \N__5913\,
            I => \N__5905\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__5908\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__5905\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5900\,
            I => \N__5896\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5899\,
            I => \N__5893\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__5896\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5893\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__5888\,
            I => \N__5880\
        );

    \I__1289\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5877\
        );

    \I__1288\ : InMux
    port map (
            O => \N__5886\,
            I => \N__5874\
        );

    \I__1287\ : InMux
    port map (
            O => \N__5885\,
            I => \N__5868\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5884\,
            I => \N__5861\
        );

    \I__1285\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5861\
        );

    \I__1284\ : InMux
    port map (
            O => \N__5880\,
            I => \N__5861\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__5877\,
            I => \N__5856\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__5874\,
            I => \N__5853\
        );

    \I__1281\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5843\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5872\,
            I => \N__5840\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5871\,
            I => \N__5837\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5868\,
            I => \N__5832\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5861\,
            I => \N__5832\
        );

    \I__1276\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5827\
        );

    \I__1275\ : InMux
    port map (
            O => \N__5859\,
            I => \N__5827\
        );

    \I__1274\ : Span4Mux_h
    port map (
            O => \N__5856\,
            I => \N__5822\
        );

    \I__1273\ : Span4Mux_h
    port map (
            O => \N__5853\,
            I => \N__5822\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5819\
        );

    \I__1271\ : InMux
    port map (
            O => \N__5851\,
            I => \N__5810\
        );

    \I__1270\ : InMux
    port map (
            O => \N__5850\,
            I => \N__5810\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5849\,
            I => \N__5810\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5848\,
            I => \N__5810\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5847\,
            I => \N__5805\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5846\,
            I => \N__5805\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__5843\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5840\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5837\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1262\ : Odrv4
    port map (
            O => \N__5832\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__5827\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__5822\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__5819\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__5810\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5805\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__5786\,
            I => \N__5775\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5785\,
            I => \N__5770\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5767\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5760\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5782\,
            I => \N__5760\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5781\,
            I => \N__5760\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5780\,
            I => \N__5755\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5779\,
            I => \N__5755\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5778\,
            I => \N__5746\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5775\,
            I => \N__5746\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5774\,
            I => \N__5746\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5746\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5770\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__5767\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5760\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5755\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__5746\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1239\ : CascadeMux
    port map (
            O => \N__5735\,
            I => \N__5731\
        );

    \I__1238\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5723\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5718\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5730\,
            I => \N__5718\
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__5729\,
            I => \N__5714\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__5728\,
            I => \N__5711\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__5727\,
            I => \N__5708\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__5726\,
            I => \N__5705\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__5723\,
            I => \N__5700\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5718\,
            I => \N__5696\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5717\,
            I => \N__5691\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5714\,
            I => \N__5691\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5711\,
            I => \N__5688\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5708\,
            I => \N__5685\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5680\
        );

    \I__1224\ : InMux
    port map (
            O => \N__5704\,
            I => \N__5680\
        );

    \I__1223\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5677\
        );

    \I__1222\ : Span4Mux_h
    port map (
            O => \N__5700\,
            I => \N__5674\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5699\,
            I => \N__5671\
        );

    \I__1220\ : Span4Mux_v
    port map (
            O => \N__5696\,
            I => \N__5666\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5691\,
            I => \N__5666\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5688\,
            I => \N__5659\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__5685\,
            I => \N__5659\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__5680\,
            I => \N__5659\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__5677\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__5674\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5671\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1212\ : Odrv4
    port map (
            O => \N__5666\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1211\ : Odrv12
    port map (
            O => \N__5659\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5648\,
            I => \N__5643\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__5647\,
            I => \N__5640\
        );

    \I__1208\ : CascadeMux
    port map (
            O => \N__5646\,
            I => \N__5634\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__5643\,
            I => \N__5631\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5640\,
            I => \N__5626\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__5639\,
            I => \N__5622\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5638\,
            I => \N__5614\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5611\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5608\
        );

    \I__1201\ : Span4Mux_v
    port map (
            O => \N__5631\,
            I => \N__5605\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5630\,
            I => \N__5602\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5629\,
            I => \N__5599\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5626\,
            I => \N__5596\
        );

    \I__1197\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5591\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5591\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5621\,
            I => \N__5586\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5620\,
            I => \N__5586\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5619\,
            I => \N__5579\
        );

    \I__1192\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5579\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5579\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__5614\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5611\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__5608\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__5605\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5602\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__5599\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1184\ : Odrv4
    port map (
            O => \N__5596\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5591\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__5586\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5579\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5555\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5555\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER19_i_0_1_0\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5552\,
            I => \N__5548\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5551\,
            I => \N__5545\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__5548\,
            I => \U712_REG_SM.N_152_0\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__5545\,
            I => \U712_REG_SM.N_152_0\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5537\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5537\,
            I => \N__5533\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5530\
        );

    \I__1171\ : Odrv4
    port map (
            O => \N__5533\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5530\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1169\ : CascadeMux
    port map (
            O => \N__5525\,
            I => \N__5522\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5518\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5521\,
            I => \N__5515\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5518\,
            I => \U712_REG_SM.STATE_COUNT_RNIVQBP4Z0Z_6\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5515\,
            I => \U712_REG_SM.STATE_COUNT_RNIVQBP4Z0Z_6\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5510\,
            I => \N__5507\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5507\,
            I => \U712_REG_SM.DS_EN_7_0\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5504\,
            I => \N__5500\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5503\,
            I => \N__5496\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5500\,
            I => \N__5493\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5499\,
            I => \N__5490\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5496\,
            I => \U712_REG_SM.N_149_0\
        );

    \I__1157\ : Odrv4
    port map (
            O => \N__5493\,
            I => \U712_REG_SM.N_149_0\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5490\,
            I => \U712_REG_SM.N_149_0\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__5483\,
            I => \N__5480\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5480\,
            I => \N__5477\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__5477\,
            I => \N__5474\
        );

    \I__1152\ : Span4Mux_v
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__5471\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_a3_0_0_3\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5462\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5467\,
            I => \N__5462\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__5462\,
            I => \U712_REG_SM.N_156_0\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5456\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5456\,
            I => \N__5451\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5448\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5454\,
            I => \N__5445\
        );

    \I__1143\ : Span4Mux_v
    port map (
            O => \N__5451\,
            I => \N__5440\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__5448\,
            I => \N__5440\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5445\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__5440\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5432\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__5432\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_a5_0_1_3\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__5429\,
            I => \N__5426\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5426\,
            I => \N__5419\
        );

    \I__1135\ : InMux
    port map (
            O => \N__5425\,
            I => \N__5419\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5424\,
            I => \N__5416\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__5419\,
            I => \U712_CHIP_RAM.N_82\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__5416\,
            I => \U712_CHIP_RAM.N_82\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5411\,
            I => \N__5406\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__5410\,
            I => \N__5403\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5409\,
            I => \N__5400\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5406\,
            I => \N__5397\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5394\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5400\,
            I => \U712_CHIP_RAM.N_105\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__5397\,
            I => \U712_CHIP_RAM.N_105\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5394\,
            I => \U712_CHIP_RAM.N_105\
        );

    \I__1123\ : InMux
    port map (
            O => \N__5387\,
            I => \N__5384\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__5384\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_ac0_1_out\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__5381\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_ac0_1_out_cascade_\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5378\,
            I => \N__5375\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__5375\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_ac0_3_0\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__5372\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_ac0_3_0_cascade_\
        );

    \I__1117\ : InMux
    port map (
            O => \N__5369\,
            I => \N__5364\
        );

    \I__1116\ : InMux
    port map (
            O => \N__5368\,
            I => \N__5357\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5367\,
            I => \N__5349\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__5364\,
            I => \N__5346\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5363\,
            I => \N__5341\
        );

    \I__1112\ : InMux
    port map (
            O => \N__5362\,
            I => \N__5341\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5361\,
            I => \N__5336\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5360\,
            I => \N__5336\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__5357\,
            I => \N__5333\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5356\,
            I => \N__5328\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5355\,
            I => \N__5328\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5354\,
            I => \N__5325\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5322\
        );

    \I__1104\ : InMux
    port map (
            O => \N__5352\,
            I => \N__5319\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5349\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__5346\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5341\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5336\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1099\ : Odrv4
    port map (
            O => \N__5333\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5328\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5325\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5322\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5319\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__5300\,
            I => \N__5296\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5299\,
            I => \N__5291\
        );

    \I__1092\ : InMux
    port map (
            O => \N__5296\,
            I => \N__5291\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5291\,
            I => \N__5287\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5290\,
            I => \N__5284\
        );

    \I__1089\ : Span4Mux_h
    port map (
            O => \N__5287\,
            I => \N__5276\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5284\,
            I => \N__5273\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5283\,
            I => \N__5270\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5282\,
            I => \N__5267\
        );

    \I__1085\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5262\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5280\,
            I => \N__5262\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5259\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__5276\,
            I => \U712_CHIP_RAM.N_36\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__5273\,
            I => \U712_CHIP_RAM.N_36\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__5270\,
            I => \U712_CHIP_RAM.N_36\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__5267\,
            I => \U712_CHIP_RAM.N_36\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__5262\,
            I => \U712_CHIP_RAM.N_36\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5259\,
            I => \U712_CHIP_RAM.N_36\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__1075\ : InMux
    port map (
            O => \N__5243\,
            I => \N__5237\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5242\,
            I => \N__5232\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5232\
        );

    \I__1072\ : InMux
    port map (
            O => \N__5240\,
            I => \N__5229\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__5237\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__5232\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5229\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__5222\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_c6_cascade_\
        );

    \I__1067\ : InMux
    port map (
            O => \N__5219\,
            I => \N__5212\
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__5218\,
            I => \N__5209\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__5217\,
            I => \N__5206\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__5216\,
            I => \N__5197\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5215\,
            I => \N__5194\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__5212\,
            I => \N__5191\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5186\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5206\,
            I => \N__5186\
        );

    \I__1059\ : InMux
    port map (
            O => \N__5205\,
            I => \N__5179\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5179\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5179\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5174\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5174\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5200\,
            I => \N__5169\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5197\,
            I => \N__5169\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5194\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1051\ : Odrv4
    port map (
            O => \N__5191\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__5186\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__5179\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5174\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5169\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5151\
        );

    \I__1045\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5146\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5154\,
            I => \N__5146\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5151\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_c4\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5146\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_c4\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__5141\,
            I => \N__5138\
        );

    \I__1040\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5133\
        );

    \I__1039\ : InMux
    port map (
            O => \N__5137\,
            I => \N__5130\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5136\,
            I => \N__5127\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__5133\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5130\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5127\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1034\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5116\
        );

    \I__1033\ : IoInMux
    port map (
            O => \N__5119\,
            I => \N__5113\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5116\,
            I => \N__5110\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__5113\,
            I => \N__5107\
        );

    \I__1030\ : Span4Mux_v
    port map (
            O => \N__5110\,
            I => \N__5104\
        );

    \I__1029\ : Span4Mux_s3_h
    port map (
            O => \N__5107\,
            I => \N__5101\
        );

    \I__1028\ : Sp12to4
    port map (
            O => \N__5104\,
            I => \N__5098\
        );

    \I__1027\ : Sp12to4
    port map (
            O => \N__5101\,
            I => \N__5095\
        );

    \I__1026\ : Span12Mux_h
    port map (
            O => \N__5098\,
            I => \N__5092\
        );

    \I__1025\ : Span12Mux_v
    port map (
            O => \N__5095\,
            I => \N__5089\
        );

    \I__1024\ : Odrv12
    port map (
            O => \N__5092\,
            I => \C1_c\
        );

    \I__1023\ : Odrv12
    port map (
            O => \N__5089\,
            I => \C1_c\
        );

    \I__1022\ : CascadeMux
    port map (
            O => \N__5084\,
            I => \N__5079\
        );

    \I__1021\ : InMux
    port map (
            O => \N__5083\,
            I => \N__5076\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5071\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5079\,
            I => \N__5071\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5076\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5071\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__1016\ : InMux
    port map (
            O => \N__5066\,
            I => \N__5060\
        );

    \I__1015\ : InMux
    port map (
            O => \N__5065\,
            I => \N__5055\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5064\,
            I => \N__5055\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5052\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5060\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__5055\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__5052\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5045\,
            I => \N__5042\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5042\,
            I => \U712_REG_SM.N_145_0\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5031\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5028\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5025\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5036\,
            I => \N__5022\
        );

    \I__1003\ : InMux
    port map (
            O => \N__5035\,
            I => \N__5017\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5034\,
            I => \N__5017\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__5031\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5028\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5025\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__5022\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5017\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__996\ : InMux
    port map (
            O => \N__5006\,
            I => \N__5003\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5003\,
            I => \N__4999\
        );

    \I__994\ : CascadeMux
    port map (
            O => \N__5002\,
            I => \N__4992\
        );

    \I__993\ : Span4Mux_h
    port map (
            O => \N__4999\,
            I => \N__4988\
        );

    \I__992\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4985\
        );

    \I__991\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4980\
        );

    \I__990\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4980\
        );

    \I__989\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4977\
        );

    \I__988\ : InMux
    port map (
            O => \N__4992\,
            I => \N__4972\
        );

    \I__987\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4972\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__4988\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__4985\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__4980\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4977\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4972\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__4961\,
            I => \U712_REG_SM.N_145_0_cascade_\
        );

    \I__980\ : CascadeMux
    port map (
            O => \N__4958\,
            I => \N__4955\
        );

    \I__979\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__4952\,
            I => \N__4947\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__4951\,
            I => \N__4941\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__4950\,
            I => \N__4938\
        );

    \I__975\ : Span4Mux_h
    port map (
            O => \N__4947\,
            I => \N__4933\
        );

    \I__974\ : InMux
    port map (
            O => \N__4946\,
            I => \N__4930\
        );

    \I__973\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4925\
        );

    \I__972\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4925\
        );

    \I__971\ : InMux
    port map (
            O => \N__4941\,
            I => \N__4922\
        );

    \I__970\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4915\
        );

    \I__969\ : InMux
    port map (
            O => \N__4937\,
            I => \N__4915\
        );

    \I__968\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4915\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__4933\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4930\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__4925\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__4922\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__4915\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__962\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4901\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4901\,
            I => \N__4898\
        );

    \I__960\ : Span4Mux_v
    port map (
            O => \N__4898\,
            I => \N__4895\
        );

    \I__959\ : Sp12to4
    port map (
            O => \N__4895\,
            I => \N__4892\
        );

    \I__958\ : Span12Mux_h
    port map (
            O => \N__4892\,
            I => \N__4889\
        );

    \I__957\ : Odrv12
    port map (
            O => \N__4889\,
            I => \C3_c\
        );

    \I__956\ : InMux
    port map (
            O => \N__4886\,
            I => \N__4879\
        );

    \I__955\ : InMux
    port map (
            O => \N__4885\,
            I => \N__4876\
        );

    \I__954\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4873\
        );

    \I__953\ : InMux
    port map (
            O => \N__4883\,
            I => \N__4868\
        );

    \I__952\ : InMux
    port map (
            O => \N__4882\,
            I => \N__4868\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4879\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__4876\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4873\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4868\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__947\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4853\
        );

    \I__946\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4853\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4853\,
            I => \N__4849\
        );

    \I__944\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4846\
        );

    \I__943\ : Span4Mux_v
    port map (
            O => \N__4849\,
            I => \N__4841\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4846\,
            I => \N__4841\
        );

    \I__941\ : Span4Mux_h
    port map (
            O => \N__4841\,
            I => \N__4837\
        );

    \I__940\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4834\
        );

    \I__939\ : Span4Mux_v
    port map (
            O => \N__4837\,
            I => \N__4831\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4834\,
            I => \N__4828\
        );

    \I__937\ : Sp12to4
    port map (
            O => \N__4831\,
            I => \N__4823\
        );

    \I__936\ : Span12Mux_v
    port map (
            O => \N__4828\,
            I => \N__4823\
        );

    \I__935\ : Odrv12
    port map (
            O => \N__4823\,
            I => \A_c_1\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__4820\,
            I => \N__4815\
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__4819\,
            I => \N__4812\
        );

    \I__932\ : CascadeMux
    port map (
            O => \N__4818\,
            I => \N__4808\
        );

    \I__931\ : InMux
    port map (
            O => \N__4815\,
            I => \N__4805\
        );

    \I__930\ : InMux
    port map (
            O => \N__4812\,
            I => \N__4800\
        );

    \I__929\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4800\
        );

    \I__928\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4797\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4805\,
            I => \N__4794\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4800\,
            I => \N__4789\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4797\,
            I => \N__4789\
        );

    \I__924\ : Span4Mux_h
    port map (
            O => \N__4794\,
            I => \N__4786\
        );

    \I__923\ : Span12Mux_v
    port map (
            O => \N__4789\,
            I => \N__4783\
        );

    \I__922\ : Sp12to4
    port map (
            O => \N__4786\,
            I => \N__4780\
        );

    \I__921\ : Span12Mux_h
    port map (
            O => \N__4783\,
            I => \N__4777\
        );

    \I__920\ : Span12Mux_v
    port map (
            O => \N__4780\,
            I => \N__4774\
        );

    \I__919\ : Odrv12
    port map (
            O => \N__4777\,
            I => \SIZ_c_1\
        );

    \I__918\ : Odrv12
    port map (
            O => \N__4774\,
            I => \SIZ_c_1\
        );

    \I__917\ : IoInMux
    port map (
            O => \N__4769\,
            I => \N__4766\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__915\ : IoSpan4Mux
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__914\ : IoSpan4Mux
    port map (
            O => \N__4760\,
            I => \N__4757\
        );

    \I__913\ : Sp12to4
    port map (
            O => \N__4757\,
            I => \N__4754\
        );

    \I__912\ : Span12Mux_s9_h
    port map (
            O => \N__4754\,
            I => \N__4751\
        );

    \I__911\ : Span12Mux_v
    port map (
            O => \N__4751\,
            I => \N__4748\
        );

    \I__910\ : Odrv12
    port map (
            O => \N__4748\,
            I => \N_22_i\
        );

    \I__909\ : IoInMux
    port map (
            O => \N__4745\,
            I => \N__4742\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4742\,
            I => \N__4739\
        );

    \I__907\ : Span4Mux_s1_h
    port map (
            O => \N__4739\,
            I => \N__4736\
        );

    \I__906\ : Span4Mux_h
    port map (
            O => \N__4736\,
            I => \N__4733\
        );

    \I__905\ : Sp12to4
    port map (
            O => \N__4733\,
            I => \N__4730\
        );

    \I__904\ : Span12Mux_s6_v
    port map (
            O => \N__4730\,
            I => \N__4727\
        );

    \I__903\ : Span12Mux_h
    port map (
            O => \N__4727\,
            I => \N__4724\
        );

    \I__902\ : Odrv12
    port map (
            O => \N__4724\,
            I => \WEn_c\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__4721\,
            I => \N__4715\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__4720\,
            I => \N__4711\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__4719\,
            I => \N__4704\
        );

    \I__898\ : InMux
    port map (
            O => \N__4718\,
            I => \N__4701\
        );

    \I__897\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4697\
        );

    \I__896\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4694\
        );

    \I__895\ : InMux
    port map (
            O => \N__4711\,
            I => \N__4689\
        );

    \I__894\ : InMux
    port map (
            O => \N__4710\,
            I => \N__4689\
        );

    \I__893\ : InMux
    port map (
            O => \N__4709\,
            I => \N__4686\
        );

    \I__892\ : InMux
    port map (
            O => \N__4708\,
            I => \N__4683\
        );

    \I__891\ : InMux
    port map (
            O => \N__4707\,
            I => \N__4678\
        );

    \I__890\ : InMux
    port map (
            O => \N__4704\,
            I => \N__4678\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4701\,
            I => \N__4673\
        );

    \I__888\ : InMux
    port map (
            O => \N__4700\,
            I => \N__4670\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__4697\,
            I => \N__4667\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__4694\,
            I => \N__4662\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4689\,
            I => \N__4662\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4686\,
            I => \N__4656\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__4683\,
            I => \N__4656\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4678\,
            I => \N__4653\
        );

    \I__881\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4650\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__4676\,
            I => \N__4647\
        );

    \I__879\ : Span4Mux_v
    port map (
            O => \N__4673\,
            I => \N__4642\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4670\,
            I => \N__4639\
        );

    \I__877\ : Span4Mux_v
    port map (
            O => \N__4667\,
            I => \N__4636\
        );

    \I__876\ : Span4Mux_h
    port map (
            O => \N__4662\,
            I => \N__4633\
        );

    \I__875\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4630\
        );

    \I__874\ : Span4Mux_h
    port map (
            O => \N__4656\,
            I => \N__4623\
        );

    \I__873\ : Span4Mux_h
    port map (
            O => \N__4653\,
            I => \N__4623\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4650\,
            I => \N__4623\
        );

    \I__871\ : InMux
    port map (
            O => \N__4647\,
            I => \N__4620\
        );

    \I__870\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4615\
        );

    \I__869\ : InMux
    port map (
            O => \N__4645\,
            I => \N__4615\
        );

    \I__868\ : Odrv4
    port map (
            O => \N__4642\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__867\ : Odrv4
    port map (
            O => \N__4639\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__866\ : Odrv4
    port map (
            O => \N__4636\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__4633\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4630\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__863\ : Odrv4
    port map (
            O => \N__4623\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4620\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4615\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__860\ : IoInMux
    port map (
            O => \N__4598\,
            I => \N__4595\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4595\,
            I => \N__4592\
        );

    \I__858\ : Span4Mux_s3_v
    port map (
            O => \N__4592\,
            I => \N__4589\
        );

    \I__857\ : Span4Mux_v
    port map (
            O => \N__4589\,
            I => \N__4586\
        );

    \I__856\ : Span4Mux_v
    port map (
            O => \N__4586\,
            I => \N__4583\
        );

    \I__855\ : Sp12to4
    port map (
            O => \N__4583\,
            I => \N__4580\
        );

    \I__854\ : Odrv12
    port map (
            O => \N__4580\,
            I => \CMA_c_10\
        );

    \I__853\ : CEMux
    port map (
            O => \N__4577\,
            I => \N__4573\
        );

    \I__852\ : CEMux
    port map (
            O => \N__4576\,
            I => \N__4567\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4573\,
            I => \N__4564\
        );

    \I__850\ : CEMux
    port map (
            O => \N__4572\,
            I => \N__4561\
        );

    \I__849\ : CEMux
    port map (
            O => \N__4571\,
            I => \N__4557\
        );

    \I__848\ : CEMux
    port map (
            O => \N__4570\,
            I => \N__4554\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4567\,
            I => \N__4548\
        );

    \I__846\ : Span4Mux_v
    port map (
            O => \N__4564\,
            I => \N__4543\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4561\,
            I => \N__4543\
        );

    \I__844\ : CEMux
    port map (
            O => \N__4560\,
            I => \N__4540\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4557\,
            I => \N__4537\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4554\,
            I => \N__4534\
        );

    \I__841\ : CEMux
    port map (
            O => \N__4553\,
            I => \N__4531\
        );

    \I__840\ : CEMux
    port map (
            O => \N__4552\,
            I => \N__4528\
        );

    \I__839\ : CEMux
    port map (
            O => \N__4551\,
            I => \N__4525\
        );

    \I__838\ : Span4Mux_v
    port map (
            O => \N__4548\,
            I => \N__4518\
        );

    \I__837\ : Span4Mux_h
    port map (
            O => \N__4543\,
            I => \N__4518\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4540\,
            I => \N__4518\
        );

    \I__835\ : Span4Mux_h
    port map (
            O => \N__4537\,
            I => \N__4511\
        );

    \I__834\ : Span4Mux_v
    port map (
            O => \N__4534\,
            I => \N__4511\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4531\,
            I => \N__4511\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4528\,
            I => \N__4508\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4525\,
            I => \N__4505\
        );

    \I__830\ : Span4Mux_h
    port map (
            O => \N__4518\,
            I => \N__4502\
        );

    \I__829\ : Sp12to4
    port map (
            O => \N__4511\,
            I => \N__4497\
        );

    \I__828\ : Sp12to4
    port map (
            O => \N__4508\,
            I => \N__4497\
        );

    \I__827\ : Span4Mux_v
    port map (
            O => \N__4505\,
            I => \N__4494\
        );

    \I__826\ : Odrv4
    port map (
            O => \N__4502\,
            I => \U712_CHIP_RAM.un1_CMA21_0_i_0\
        );

    \I__825\ : Odrv12
    port map (
            O => \N__4497\,
            I => \U712_CHIP_RAM.un1_CMA21_0_i_0\
        );

    \I__824\ : Odrv4
    port map (
            O => \N__4494\,
            I => \U712_CHIP_RAM.un1_CMA21_0_i_0\
        );

    \I__823\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4481\
        );

    \I__822\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4481\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4481\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_10_u_0_2_0\
        );

    \I__820\ : InMux
    port map (
            O => \N__4478\,
            I => \N__4472\
        );

    \I__819\ : InMux
    port map (
            O => \N__4477\,
            I => \N__4472\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4472\,
            I => \U712_CHIP_RAM.N_13\
        );

    \I__817\ : CascadeMux
    port map (
            O => \N__4469\,
            I => \U712_CHIP_RAM.N_13_cascade_\
        );

    \I__816\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4463\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4463\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_0_a2_0\
        );

    \I__814\ : IoInMux
    port map (
            O => \N__4460\,
            I => \N__4457\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__4457\,
            I => \N__4454\
        );

    \I__812\ : IoSpan4Mux
    port map (
            O => \N__4454\,
            I => \N__4451\
        );

    \I__811\ : Span4Mux_s1_h
    port map (
            O => \N__4451\,
            I => \N__4448\
        );

    \I__810\ : Sp12to4
    port map (
            O => \N__4448\,
            I => \N__4445\
        );

    \I__809\ : Span12Mux_h
    port map (
            O => \N__4445\,
            I => \N__4442\
        );

    \I__808\ : Span12Mux_v
    port map (
            O => \N__4442\,
            I => \N__4439\
        );

    \I__807\ : Odrv12
    port map (
            O => \N__4439\,
            I => \N_23_i\
        );

    \I__806\ : IoInMux
    port map (
            O => \N__4436\,
            I => \N__4433\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__4433\,
            I => \N__4430\
        );

    \I__804\ : Span4Mux_s2_h
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__803\ : Span4Mux_h
    port map (
            O => \N__4427\,
            I => \N__4424\
        );

    \I__802\ : Sp12to4
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__801\ : Span12Mux_s9_v
    port map (
            O => \N__4421\,
            I => \N__4418\
        );

    \I__800\ : Span12Mux_h
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__799\ : Odrv12
    port map (
            O => \N__4415\,
            I => \CUMBEn_c\
        );

    \I__798\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4408\
        );

    \I__797\ : InMux
    port map (
            O => \N__4411\,
            I => \N__4405\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4408\,
            I => \U712_REG_SM.N_148_0\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__4405\,
            I => \U712_REG_SM.N_148_0\
        );

    \I__794\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4396\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__4399\,
            I => \N__4393\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4396\,
            I => \N__4390\
        );

    \I__791\ : InMux
    port map (
            O => \N__4393\,
            I => \N__4387\
        );

    \I__790\ : Span4Mux_h
    port map (
            O => \N__4390\,
            I => \N__4384\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__4387\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__788\ : Odrv4
    port map (
            O => \N__4384\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__787\ : CascadeMux
    port map (
            O => \N__4379\,
            I => \U712_REG_SM.N_155_0_cascade_\
        );

    \I__786\ : InMux
    port map (
            O => \N__4376\,
            I => \N__4372\
        );

    \I__785\ : InMux
    port map (
            O => \N__4375\,
            I => \N__4368\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4372\,
            I => \N__4362\
        );

    \I__783\ : InMux
    port map (
            O => \N__4371\,
            I => \N__4359\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__4368\,
            I => \N__4356\
        );

    \I__781\ : InMux
    port map (
            O => \N__4367\,
            I => \N__4351\
        );

    \I__780\ : InMux
    port map (
            O => \N__4366\,
            I => \N__4351\
        );

    \I__779\ : InMux
    port map (
            O => \N__4365\,
            I => \N__4348\
        );

    \I__778\ : Odrv4
    port map (
            O => \N__4362\,
            I => \U712_CHIP_RAM.N_100\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__4359\,
            I => \U712_CHIP_RAM.N_100\
        );

    \I__776\ : Odrv4
    port map (
            O => \N__4356\,
            I => \U712_CHIP_RAM.N_100\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4351\,
            I => \U712_CHIP_RAM.N_100\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4348\,
            I => \U712_CHIP_RAM.N_100\
        );

    \I__773\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4334\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__4334\,
            I => \N__4328\
        );

    \I__771\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4325\
        );

    \I__770\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4320\
        );

    \I__769\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4320\
        );

    \I__768\ : Odrv4
    port map (
            O => \N__4328\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_2\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4325\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_2\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4320\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_2\
        );

    \I__765\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4310\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4310\,
            I => \U712_CHIP_RAM.N_87\
        );

    \I__763\ : InMux
    port map (
            O => \N__4307\,
            I => \N__4304\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4304\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a5_1\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__4301\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_a5_0_0_3_cascade_\
        );

    \I__760\ : CascadeMux
    port map (
            O => \N__4298\,
            I => \U712_CHIP_RAM.N_21_cascade_\
        );

    \I__759\ : InMux
    port map (
            O => \N__4295\,
            I => \N__4292\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4292\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_i_1\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__4289\,
            I => \U712_CHIP_RAM.N_116_cascade_\
        );

    \I__756\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4282\
        );

    \I__755\ : InMux
    port map (
            O => \N__4285\,
            I => \N__4279\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__4282\,
            I => \U712_CHIP_RAM.N_117\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4279\,
            I => \U712_CHIP_RAM.N_117\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__4274\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_67_i_i_0_cascade_\
        );

    \I__751\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4268\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__4268\,
            I => \U712_CHIP_RAM.N_26\
        );

    \I__749\ : InMux
    port map (
            O => \N__4265\,
            I => \N__4260\
        );

    \I__748\ : InMux
    port map (
            O => \N__4264\,
            I => \N__4257\
        );

    \I__747\ : InMux
    port map (
            O => \N__4263\,
            I => \N__4254\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4260\,
            I => \U712_CHIP_RAM.N_116\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4257\,
            I => \U712_CHIP_RAM.N_116\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__4254\,
            I => \U712_CHIP_RAM.N_116\
        );

    \I__743\ : CascadeMux
    port map (
            O => \N__4247\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_1_3_cascade_\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__741\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4238\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4238\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_2_3\
        );

    \I__739\ : InMux
    port map (
            O => \N__4235\,
            I => \N__4232\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4232\,
            I => \N__4229\
        );

    \I__737\ : Span4Mux_h
    port map (
            O => \N__4229\,
            I => \N__4225\
        );

    \I__736\ : InMux
    port map (
            O => \N__4228\,
            I => \N__4222\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__4225\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__4222\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__4217\,
            I => \N__4214\
        );

    \I__732\ : InMux
    port map (
            O => \N__4214\,
            I => \N__4210\
        );

    \I__731\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4205\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4210\,
            I => \N__4202\
        );

    \I__729\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4199\
        );

    \I__728\ : InMux
    port map (
            O => \N__4208\,
            I => \N__4196\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__4205\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__4202\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4199\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__4196\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__723\ : InMux
    port map (
            O => \N__4187\,
            I => \N__4183\
        );

    \I__722\ : InMux
    port map (
            O => \N__4186\,
            I => \N__4179\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4183\,
            I => \N__4176\
        );

    \I__720\ : InMux
    port map (
            O => \N__4182\,
            I => \N__4173\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__4179\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__718\ : Odrv4
    port map (
            O => \N__4176\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4173\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__4166\,
            I => \U712_REG_SM.N_146_0_cascade_\
        );

    \I__715\ : InMux
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__4160\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa_1\
        );

    \I__713\ : InMux
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__711\ : Span4Mux_h
    port map (
            O => \N__4151\,
            I => \N__4148\
        );

    \I__710\ : Sp12to4
    port map (
            O => \N__4148\,
            I => \N__4145\
        );

    \I__709\ : Span12Mux_v
    port map (
            O => \N__4145\,
            I => \N__4142\
        );

    \I__708\ : Odrv12
    port map (
            O => \N__4142\,
            I => \A_c_17\
        );

    \I__707\ : IoInMux
    port map (
            O => \N__4139\,
            I => \N__4136\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4136\,
            I => \N__4133\
        );

    \I__705\ : Span12Mux_s6_h
    port map (
            O => \N__4133\,
            I => \N__4130\
        );

    \I__704\ : Span12Mux_h
    port map (
            O => \N__4130\,
            I => \N__4127\
        );

    \I__703\ : Odrv12
    port map (
            O => \N__4127\,
            I => \CMA_c_8\
        );

    \I__702\ : InMux
    port map (
            O => \N__4124\,
            I => \N__4121\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__4121\,
            I => \N__4118\
        );

    \I__700\ : Span4Mux_h
    port map (
            O => \N__4118\,
            I => \N__4115\
        );

    \I__699\ : Sp12to4
    port map (
            O => \N__4115\,
            I => \N__4112\
        );

    \I__698\ : Span12Mux_v
    port map (
            O => \N__4112\,
            I => \N__4109\
        );

    \I__697\ : Odrv12
    port map (
            O => \N__4109\,
            I => \A_c_19\
        );

    \I__696\ : IoInMux
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4103\,
            I => \N__4100\
        );

    \I__694\ : IoSpan4Mux
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__693\ : Span4Mux_s2_h
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__692\ : Span4Mux_h
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__691\ : Sp12to4
    port map (
            O => \N__4091\,
            I => \N__4088\
        );

    \I__690\ : Span12Mux_h
    port map (
            O => \N__4088\,
            I => \N__4085\
        );

    \I__689\ : Odrv12
    port map (
            O => \N__4085\,
            I => \CMA_c_9\
        );

    \I__688\ : InMux
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__4079\,
            I => \U712_CHIP_RAM.un1_CMA21_0_i\
        );

    \I__686\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4073\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_10_u_0_1_0\
        );

    \I__684\ : InMux
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4067\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\
        );

    \I__682\ : InMux
    port map (
            O => \N__4064\,
            I => \N__4060\
        );

    \I__681\ : InMux
    port map (
            O => \N__4063\,
            I => \N__4057\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__4060\,
            I => \U712_CHIP_RAM.N_40\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__4057\,
            I => \U712_CHIP_RAM.N_40\
        );

    \I__678\ : InMux
    port map (
            O => \N__4052\,
            I => \N__4049\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4049\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_1\
        );

    \I__676\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4043\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__4043\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_6_tz\
        );

    \I__674\ : CascadeMux
    port map (
            O => \N__4040\,
            I => \U712_REG_SM.N_148_0_cascade_\
        );

    \I__673\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4034\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4034\,
            I => \U712_REG_SM.N_157_0\
        );

    \I__671\ : CascadeMux
    port map (
            O => \N__4031\,
            I => \U712_REG_SM.N_157_0_cascade_\
        );

    \I__670\ : InMux
    port map (
            O => \N__4028\,
            I => \N__4025\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__4025\,
            I => \U712_REG_SM.REG_TACK_7_0\
        );

    \I__668\ : InMux
    port map (
            O => \N__4022\,
            I => \N__4016\
        );

    \I__667\ : InMux
    port map (
            O => \N__4021\,
            I => \N__4016\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__4016\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__665\ : InMux
    port map (
            O => \N__4013\,
            I => \N__4006\
        );

    \I__664\ : InMux
    port map (
            O => \N__4012\,
            I => \N__4006\
        );

    \I__663\ : InMux
    port map (
            O => \N__4011\,
            I => \N__4003\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__4006\,
            I => \N__4000\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4003\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__4000\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__3995\,
            I => \N__3991\
        );

    \I__658\ : InMux
    port map (
            O => \N__3994\,
            I => \N__3986\
        );

    \I__657\ : InMux
    port map (
            O => \N__3991\,
            I => \N__3986\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3986\,
            I => \U712_REG_SM.un1_STATE_COUNT_3_0_1\
        );

    \I__655\ : CascadeMux
    port map (
            O => \N__3983\,
            I => \U712_CHIP_RAM.N_110_cascade_\
        );

    \I__654\ : InMux
    port map (
            O => \N__3980\,
            I => \N__3977\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3977\,
            I => \U712_CHIP_RAM.N_58\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__3974\,
            I => \U712_CHIP_RAM.N_58_cascade_\
        );

    \I__651\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3965\
        );

    \I__650\ : InMux
    port map (
            O => \N__3970\,
            I => \N__3965\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3965\,
            I => \U712_CHIP_RAM.N_118\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__3962\,
            I => \U712_CHIP_RAM.N_118_cascade_\
        );

    \I__647\ : InMux
    port map (
            O => \N__3959\,
            I => \N__3956\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3956\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_0_sqmuxa\
        );

    \I__645\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3950\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3950\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_o2_0_0\
        );

    \I__643\ : InMux
    port map (
            O => \N__3947\,
            I => \N__3943\
        );

    \I__642\ : InMux
    port map (
            O => \N__3946\,
            I => \N__3940\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3943\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3940\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__639\ : InMux
    port map (
            O => \N__3935\,
            I => \N__3927\
        );

    \I__638\ : InMux
    port map (
            O => \N__3934\,
            I => \N__3920\
        );

    \I__637\ : InMux
    port map (
            O => \N__3933\,
            I => \N__3920\
        );

    \I__636\ : InMux
    port map (
            O => \N__3932\,
            I => \N__3920\
        );

    \I__635\ : InMux
    port map (
            O => \N__3931\,
            I => \N__3915\
        );

    \I__634\ : InMux
    port map (
            O => \N__3930\,
            I => \N__3915\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3927\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3920\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3915\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__630\ : InMux
    port map (
            O => \N__3908\,
            I => \N__3905\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3905\,
            I => \N__3898\
        );

    \I__628\ : InMux
    port map (
            O => \N__3904\,
            I => \N__3893\
        );

    \I__627\ : InMux
    port map (
            O => \N__3903\,
            I => \N__3893\
        );

    \I__626\ : InMux
    port map (
            O => \N__3902\,
            I => \N__3888\
        );

    \I__625\ : InMux
    port map (
            O => \N__3901\,
            I => \N__3888\
        );

    \I__624\ : Odrv4
    port map (
            O => \N__3898\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3893\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3888\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__3881\,
            I => \U712_CHIP_RAM.N_40_cascade_\
        );

    \I__620\ : InMux
    port map (
            O => \N__3878\,
            I => \N__3870\
        );

    \I__619\ : InMux
    port map (
            O => \N__3877\,
            I => \N__3870\
        );

    \I__618\ : InMux
    port map (
            O => \N__3876\,
            I => \N__3867\
        );

    \I__617\ : InMux
    port map (
            O => \N__3875\,
            I => \N__3864\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__3870\,
            I => \U712_CHIP_RAM.SDRAM_CMD14\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3867\,
            I => \U712_CHIP_RAM.SDRAM_CMD14\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3864\,
            I => \U712_CHIP_RAM.SDRAM_CMD14\
        );

    \I__613\ : CascadeMux
    port map (
            O => \N__3857\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\
        );

    \I__612\ : CascadeMux
    port map (
            O => \N__3854\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_2_cascade_\
        );

    \I__611\ : InMux
    port map (
            O => \N__3851\,
            I => \N__3848\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3848\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_3_0_0\
        );

    \I__609\ : InMux
    port map (
            O => \N__3845\,
            I => \N__3839\
        );

    \I__608\ : InMux
    port map (
            O => \N__3844\,
            I => \N__3839\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3839\,
            I => \U712_CHIP_RAM.N_83\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__3836\,
            I => \N__3832\
        );

    \I__605\ : InMux
    port map (
            O => \N__3835\,
            I => \N__3828\
        );

    \I__604\ : InMux
    port map (
            O => \N__3832\,
            I => \N__3825\
        );

    \I__603\ : InMux
    port map (
            O => \N__3831\,
            I => \N__3822\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3828\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3825\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3822\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__3815\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1_cascade_\
        );

    \I__598\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3807\
        );

    \I__597\ : InMux
    port map (
            O => \N__3811\,
            I => \N__3804\
        );

    \I__596\ : InMux
    port map (
            O => \N__3810\,
            I => \N__3801\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3807\,
            I => \U712_CHIP_RAM.CPU_CYCLEZ0\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3804\,
            I => \U712_CHIP_RAM.CPU_CYCLEZ0\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3801\,
            I => \U712_CHIP_RAM.CPU_CYCLEZ0\
        );

    \I__592\ : InMux
    port map (
            O => \N__3794\,
            I => \N__3791\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3791\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_i_1\
        );

    \I__590\ : InMux
    port map (
            O => \N__3788\,
            I => \N__3785\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3785\,
            I => \U712_CHIP_RAM.N_110\
        );

    \I__588\ : IoInMux
    port map (
            O => \N__3782\,
            I => \N__3779\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__3779\,
            I => \N__3776\
        );

    \I__586\ : Span12Mux_s2_v
    port map (
            O => \N__3776\,
            I => \N__3773\
        );

    \I__585\ : Span12Mux_v
    port map (
            O => \N__3773\,
            I => \N__3770\
        );

    \I__584\ : Odrv12
    port map (
            O => \N__3770\,
            I => \CLLBEn_c\
        );

    \I__583\ : InMux
    port map (
            O => \N__3767\,
            I => \N__3764\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3764\,
            I => \U712_REG_SM.N_160\
        );

    \I__581\ : InMux
    port map (
            O => \N__3761\,
            I => \N__3758\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3758\,
            I => \U712_CHIP_RAM.A_m_14\
        );

    \I__579\ : InMux
    port map (
            O => \N__3755\,
            I => \N__3752\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3752\,
            I => \N__3749\
        );

    \I__577\ : Span4Mux_v
    port map (
            O => \N__3749\,
            I => \N__3746\
        );

    \I__576\ : Span4Mux_v
    port map (
            O => \N__3746\,
            I => \N__3743\
        );

    \I__575\ : Sp12to4
    port map (
            O => \N__3743\,
            I => \N__3740\
        );

    \I__574\ : Odrv12
    port map (
            O => \N__3740\,
            I => \A_c_7\
        );

    \I__573\ : IoInMux
    port map (
            O => \N__3737\,
            I => \N__3734\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3734\,
            I => \N__3731\
        );

    \I__571\ : IoSpan4Mux
    port map (
            O => \N__3731\,
            I => \N__3728\
        );

    \I__570\ : Sp12to4
    port map (
            O => \N__3728\,
            I => \N__3725\
        );

    \I__569\ : Span12Mux_s7_h
    port map (
            O => \N__3725\,
            I => \N__3722\
        );

    \I__568\ : Span12Mux_h
    port map (
            O => \N__3722\,
            I => \N__3719\
        );

    \I__567\ : Odrv12
    port map (
            O => \N__3719\,
            I => \CMA_c_5\
        );

    \I__566\ : InMux
    port map (
            O => \N__3716\,
            I => \N__3713\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3713\,
            I => \U712_CHIP_RAM.A_m_10\
        );

    \I__564\ : InMux
    port map (
            O => \N__3710\,
            I => \N__3707\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3707\,
            I => \N__3704\
        );

    \I__562\ : Sp12to4
    port map (
            O => \N__3704\,
            I => \N__3701\
        );

    \I__561\ : Span12Mux_v
    port map (
            O => \N__3701\,
            I => \N__3698\
        );

    \I__560\ : Span12Mux_h
    port map (
            O => \N__3698\,
            I => \N__3695\
        );

    \I__559\ : Odrv12
    port map (
            O => \N__3695\,
            I => \A_c_3\
        );

    \I__558\ : IoInMux
    port map (
            O => \N__3692\,
            I => \N__3689\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3689\,
            I => \N__3686\
        );

    \I__556\ : Span12Mux_s1_v
    port map (
            O => \N__3686\,
            I => \N__3683\
        );

    \I__555\ : Span12Mux_v
    port map (
            O => \N__3683\,
            I => \N__3680\
        );

    \I__554\ : Odrv12
    port map (
            O => \N__3680\,
            I => \CMA_c_1\
        );

    \I__553\ : SRMux
    port map (
            O => \N__3677\,
            I => \N__3674\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3674\,
            I => \N__3671\
        );

    \I__551\ : Odrv4
    port map (
            O => \N__3671\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__550\ : InMux
    port map (
            O => \N__3668\,
            I => \N__3665\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3665\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__3662\,
            I => \U712_CHIP_RAM.N_80_cascade_\
        );

    \I__547\ : InMux
    port map (
            O => \N__3659\,
            I => \N__3656\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3656\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__545\ : InMux
    port map (
            O => \N__3653\,
            I => \N__3650\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3650\,
            I => \N__3647\
        );

    \I__543\ : Span4Mux_v
    port map (
            O => \N__3647\,
            I => \N__3644\
        );

    \I__542\ : Sp12to4
    port map (
            O => \N__3644\,
            I => \N__3641\
        );

    \I__541\ : Span12Mux_h
    port map (
            O => \N__3641\,
            I => \N__3638\
        );

    \I__540\ : Span12Mux_v
    port map (
            O => \N__3638\,
            I => \N__3635\
        );

    \I__539\ : Odrv12
    port map (
            O => \N__3635\,
            I => \DBRn_c\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__3632\,
            I => \N__3629\
        );

    \I__537\ : InMux
    port map (
            O => \N__3629\,
            I => \N__3625\
        );

    \I__536\ : InMux
    port map (
            O => \N__3628\,
            I => \N__3622\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3625\,
            I => \CPU_TACKm\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3622\,
            I => \CPU_TACKm\
        );

    \I__533\ : CascadeMux
    port map (
            O => \N__3617\,
            I => \N__3614\
        );

    \I__532\ : InMux
    port map (
            O => \N__3614\,
            I => \N__3610\
        );

    \I__531\ : InMux
    port map (
            O => \N__3613\,
            I => \N__3607\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3610\,
            I => \REG_TACK\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3607\,
            I => \REG_TACK\
        );

    \I__528\ : InMux
    port map (
            O => \N__3602\,
            I => \N__3599\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3599\,
            I => \N__3595\
        );

    \I__526\ : InMux
    port map (
            O => \N__3598\,
            I => \N__3592\
        );

    \I__525\ : Span4Mux_h
    port map (
            O => \N__3595\,
            I => \N__3586\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3592\,
            I => \N__3586\
        );

    \I__523\ : InMux
    port map (
            O => \N__3591\,
            I => \N__3583\
        );

    \I__522\ : Span4Mux_v
    port map (
            O => \N__3586\,
            I => \N__3580\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3583\,
            I => \N__3577\
        );

    \I__520\ : Span4Mux_h
    port map (
            O => \N__3580\,
            I => \N__3574\
        );

    \I__519\ : Span12Mux_h
    port map (
            O => \N__3577\,
            I => \N__3571\
        );

    \I__518\ : Sp12to4
    port map (
            O => \N__3574\,
            I => \N__3568\
        );

    \I__517\ : Span12Mux_v
    port map (
            O => \N__3571\,
            I => \N__3565\
        );

    \I__516\ : Odrv12
    port map (
            O => \N__3568\,
            I => \TSn_c\
        );

    \I__515\ : Odrv12
    port map (
            O => \N__3565\,
            I => \TSn_c\
        );

    \I__514\ : InMux
    port map (
            O => \N__3560\,
            I => \N__3556\
        );

    \I__513\ : InMux
    port map (
            O => \N__3559\,
            I => \N__3553\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3556\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3553\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__510\ : InMux
    port map (
            O => \N__3548\,
            I => \N__3544\
        );

    \I__509\ : InMux
    port map (
            O => \N__3547\,
            I => \N__3541\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3544\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3541\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__506\ : InMux
    port map (
            O => \N__3536\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__505\ : InMux
    port map (
            O => \N__3533\,
            I => \N__3529\
        );

    \I__504\ : InMux
    port map (
            O => \N__3532\,
            I => \N__3526\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3529\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3526\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__501\ : InMux
    port map (
            O => \N__3521\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__3518\,
            I => \N__3514\
        );

    \I__499\ : InMux
    port map (
            O => \N__3517\,
            I => \N__3511\
        );

    \I__498\ : InMux
    port map (
            O => \N__3514\,
            I => \N__3508\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3511\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3508\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__495\ : InMux
    port map (
            O => \N__3503\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__494\ : InMux
    port map (
            O => \N__3500\,
            I => \N__3496\
        );

    \I__493\ : InMux
    port map (
            O => \N__3499\,
            I => \N__3493\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3496\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3493\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__490\ : InMux
    port map (
            O => \N__3488\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__489\ : InMux
    port map (
            O => \N__3485\,
            I => \N__3481\
        );

    \I__488\ : InMux
    port map (
            O => \N__3484\,
            I => \N__3478\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3481\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3478\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__485\ : InMux
    port map (
            O => \N__3473\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__484\ : InMux
    port map (
            O => \N__3470\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__3467\,
            I => \N__3463\
        );

    \I__482\ : InMux
    port map (
            O => \N__3466\,
            I => \N__3460\
        );

    \I__481\ : InMux
    port map (
            O => \N__3463\,
            I => \N__3457\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3460\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3457\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__478\ : ClkMux
    port map (
            O => \N__3452\,
            I => \N__3449\
        );

    \I__477\ : GlobalMux
    port map (
            O => \N__3449\,
            I => \N__3446\
        );

    \I__476\ : gio2CtrlBuf
    port map (
            O => \N__3446\,
            I => \C1_c_g\
        );

    \I__475\ : CascadeMux
    port map (
            O => \N__3443\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1_0_cascade_\
        );

    \I__474\ : CascadeMux
    port map (
            O => \N__3440\,
            I => \N__3436\
        );

    \I__473\ : InMux
    port map (
            O => \N__3439\,
            I => \N__3433\
        );

    \I__472\ : InMux
    port map (
            O => \N__3436\,
            I => \N__3430\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3433\,
            I => \N__3427\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3430\,
            I => \N__3424\
        );

    \I__469\ : Span12Mux_h
    port map (
            O => \N__3427\,
            I => \N__3420\
        );

    \I__468\ : Span4Mux_h
    port map (
            O => \N__3424\,
            I => \N__3417\
        );

    \I__467\ : IoInMux
    port map (
            O => \N__3423\,
            I => \N__3414\
        );

    \I__466\ : Span12Mux_v
    port map (
            O => \N__3420\,
            I => \N__3409\
        );

    \I__465\ : Sp12to4
    port map (
            O => \N__3417\,
            I => \N__3409\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3414\,
            I => \N__3406\
        );

    \I__463\ : Span12Mux_v
    port map (
            O => \N__3409\,
            I => \N__3403\
        );

    \I__462\ : IoSpan4Mux
    port map (
            O => \N__3406\,
            I => \N__3400\
        );

    \I__461\ : Odrv12
    port map (
            O => \N__3403\,
            I => \RAMENn_c\
        );

    \I__460\ : Odrv4
    port map (
            O => \N__3400\,
            I => \RAMENn_c\
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__3395\,
            I => \N__3392\
        );

    \I__458\ : InMux
    port map (
            O => \N__3392\,
            I => \N__3389\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3389\,
            I => \N__3385\
        );

    \I__456\ : InMux
    port map (
            O => \N__3388\,
            I => \N__3382\
        );

    \I__455\ : Odrv4
    port map (
            O => \N__3385\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__3382\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__3377\,
            I => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\
        );

    \I__452\ : CascadeMux
    port map (
            O => \N__3374\,
            I => \U712_CYCLE_TERM.N_45_0_0_en_cascade_\
        );

    \I__451\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3366\
        );

    \I__450\ : InMux
    port map (
            O => \N__3370\,
            I => \N__3361\
        );

    \I__449\ : InMux
    port map (
            O => \N__3369\,
            I => \N__3361\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3366\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3361\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__3356\,
            I => \N__3352\
        );

    \I__445\ : InMux
    port map (
            O => \N__3355\,
            I => \N__3349\
        );

    \I__444\ : InMux
    port map (
            O => \N__3352\,
            I => \N__3345\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__3349\,
            I => \N__3342\
        );

    \I__442\ : InMux
    port map (
            O => \N__3348\,
            I => \N__3339\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3345\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__440\ : Odrv4
    port map (
            O => \N__3342\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3339\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__438\ : InMux
    port map (
            O => \N__3332\,
            I => \N__3329\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__3329\,
            I => \N__3326\
        );

    \I__436\ : Span12Mux_s11_v
    port map (
            O => \N__3326\,
            I => \N__3323\
        );

    \I__435\ : Odrv12
    port map (
            O => \N__3323\,
            I => \TACK_EN_i_ess\
        );

    \I__434\ : CEMux
    port map (
            O => \N__3320\,
            I => \N__3317\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3317\,
            I => \N__3314\
        );

    \I__432\ : Span4Mux_v
    port map (
            O => \N__3314\,
            I => \N__3311\
        );

    \I__431\ : Odrv4
    port map (
            O => \N__3311\,
            I => \U712_CYCLE_TERM.N_45_0_0_en_0\
        );

    \I__430\ : IoInMux
    port map (
            O => \N__3308\,
            I => \N__3305\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3305\,
            I => \N__3302\
        );

    \I__428\ : Span4Mux_s3_v
    port map (
            O => \N__3302\,
            I => \N__3299\
        );

    \I__427\ : Odrv4
    port map (
            O => \N__3299\,
            I => \VBENn_c\
        );

    \I__426\ : InMux
    port map (
            O => \N__3296\,
            I => \N__3293\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3293\,
            I => \N__3290\
        );

    \I__424\ : Span4Mux_v
    port map (
            O => \N__3290\,
            I => \N__3287\
        );

    \I__423\ : Span4Mux_v
    port map (
            O => \N__3287\,
            I => \N__3284\
        );

    \I__422\ : Sp12to4
    port map (
            O => \N__3284\,
            I => \N__3281\
        );

    \I__421\ : Span12Mux_h
    port map (
            O => \N__3281\,
            I => \N__3278\
        );

    \I__420\ : Odrv12
    port map (
            O => \N__3278\,
            I => \A_c_14\
        );

    \I__419\ : InMux
    port map (
            O => \N__3275\,
            I => \N__3272\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3272\,
            I => \N__3269\
        );

    \I__417\ : Span4Mux_v
    port map (
            O => \N__3269\,
            I => \N__3266\
        );

    \I__416\ : Sp12to4
    port map (
            O => \N__3266\,
            I => \N__3263\
        );

    \I__415\ : Span12Mux_h
    port map (
            O => \N__3263\,
            I => \N__3260\
        );

    \I__414\ : Odrv12
    port map (
            O => \N__3260\,
            I => \A_c_10\
        );

    \I__413\ : InMux
    port map (
            O => \N__3257\,
            I => \N__3253\
        );

    \I__412\ : InMux
    port map (
            O => \N__3256\,
            I => \N__3250\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__3253\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3250\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__409\ : InMux
    port map (
            O => \N__3245\,
            I => \bfn_8_10_0_\
        );

    \I__408\ : InMux
    port map (
            O => \N__3242\,
            I => \N__3238\
        );

    \I__407\ : InMux
    port map (
            O => \N__3241\,
            I => \N__3235\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3238\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__3235\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__404\ : InMux
    port map (
            O => \N__3230\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__403\ : InMux
    port map (
            O => \N__3227\,
            I => \N__3224\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3224\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__401\ : InMux
    port map (
            O => \N__3221\,
            I => \N__3218\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3218\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__399\ : InMux
    port map (
            O => \N__3215\,
            I => \N__3208\
        );

    \I__398\ : InMux
    port map (
            O => \N__3214\,
            I => \N__3208\
        );

    \I__397\ : InMux
    port map (
            O => \N__3213\,
            I => \N__3205\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3208\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__3205\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__394\ : InMux
    port map (
            O => \N__3200\,
            I => \N__3197\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3197\,
            I => \U712_REG_SM.STATE_COUNT5\
        );

    \I__392\ : InMux
    port map (
            O => \N__3194\,
            I => \N__3191\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__3191\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\
        );

    \I__390\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3184\
        );

    \I__389\ : InMux
    port map (
            O => \N__3187\,
            I => \N__3181\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3184\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__3181\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__386\ : CascadeMux
    port map (
            O => \N__3176\,
            I => \N__3172\
        );

    \I__385\ : InMux
    port map (
            O => \N__3175\,
            I => \N__3167\
        );

    \I__384\ : InMux
    port map (
            O => \N__3172\,
            I => \N__3164\
        );

    \I__383\ : InMux
    port map (
            O => \N__3171\,
            I => \N__3159\
        );

    \I__382\ : InMux
    port map (
            O => \N__3170\,
            I => \N__3159\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__3167\,
            I => \N__3156\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__3164\,
            I => \N__3151\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__3159\,
            I => \N__3151\
        );

    \I__378\ : Span4Mux_v
    port map (
            O => \N__3156\,
            I => \N__3148\
        );

    \I__377\ : Span4Mux_h
    port map (
            O => \N__3151\,
            I => \N__3145\
        );

    \I__376\ : Span4Mux_v
    port map (
            O => \N__3148\,
            I => \N__3142\
        );

    \I__375\ : Span4Mux_h
    port map (
            O => \N__3145\,
            I => \N__3139\
        );

    \I__374\ : Sp12to4
    port map (
            O => \N__3142\,
            I => \N__3136\
        );

    \I__373\ : Sp12to4
    port map (
            O => \N__3139\,
            I => \N__3133\
        );

    \I__372\ : Span12Mux_h
    port map (
            O => \N__3136\,
            I => \N__3128\
        );

    \I__371\ : Span12Mux_v
    port map (
            O => \N__3133\,
            I => \N__3128\
        );

    \I__370\ : Odrv12
    port map (
            O => \N__3128\,
            I => \CLK40_OUT_i\
        );

    \I__369\ : InMux
    port map (
            O => \N__3125\,
            I => \N__3119\
        );

    \I__368\ : InMux
    port map (
            O => \N__3124\,
            I => \N__3112\
        );

    \I__367\ : InMux
    port map (
            O => \N__3123\,
            I => \N__3112\
        );

    \I__366\ : InMux
    port map (
            O => \N__3122\,
            I => \N__3112\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__3119\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3112\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__363\ : InMux
    port map (
            O => \N__3107\,
            I => \N__3104\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__3104\,
            I => \N__3101\
        );

    \I__361\ : Span4Mux_v
    port map (
            O => \N__3101\,
            I => \N__3098\
        );

    \I__360\ : Span4Mux_v
    port map (
            O => \N__3098\,
            I => \N__3095\
        );

    \I__359\ : Sp12to4
    port map (
            O => \N__3095\,
            I => \N__3092\
        );

    \I__358\ : Odrv12
    port map (
            O => \N__3092\,
            I => \A_c_8\
        );

    \I__357\ : CascadeMux
    port map (
            O => \N__3089\,
            I => \N__3086\
        );

    \I__356\ : InMux
    port map (
            O => \N__3086\,
            I => \N__3083\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__3083\,
            I => \N__3080\
        );

    \I__354\ : Span4Mux_v
    port map (
            O => \N__3080\,
            I => \N__3077\
        );

    \I__353\ : Span4Mux_v
    port map (
            O => \N__3077\,
            I => \N__3074\
        );

    \I__352\ : Sp12to4
    port map (
            O => \N__3074\,
            I => \N__3071\
        );

    \I__351\ : Odrv12
    port map (
            O => \N__3071\,
            I => \A_c_15\
        );

    \I__350\ : IoInMux
    port map (
            O => \N__3068\,
            I => \N__3065\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__3065\,
            I => \N__3062\
        );

    \I__348\ : Span12Mux_s10_h
    port map (
            O => \N__3062\,
            I => \N__3059\
        );

    \I__347\ : Span12Mux_h
    port map (
            O => \N__3059\,
            I => \N__3056\
        );

    \I__346\ : Odrv12
    port map (
            O => \N__3056\,
            I => \CMA_c_6\
        );

    \I__345\ : InMux
    port map (
            O => \N__3053\,
            I => \N__3050\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__3050\,
            I => \N__3047\
        );

    \I__343\ : Span12Mux_v
    port map (
            O => \N__3047\,
            I => \N__3044\
        );

    \I__342\ : Odrv12
    port map (
            O => \N__3044\,
            I => \A_c_18\
        );

    \I__341\ : InMux
    port map (
            O => \N__3041\,
            I => \N__3038\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__3038\,
            I => \N__3035\
        );

    \I__339\ : Span4Mux_v
    port map (
            O => \N__3035\,
            I => \N__3032\
        );

    \I__338\ : Span4Mux_v
    port map (
            O => \N__3032\,
            I => \N__3029\
        );

    \I__337\ : Sp12to4
    port map (
            O => \N__3029\,
            I => \N__3026\
        );

    \I__336\ : Odrv12
    port map (
            O => \N__3026\,
            I => \A_c_16\
        );

    \I__335\ : IoInMux
    port map (
            O => \N__3023\,
            I => \N__3020\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__3020\,
            I => \N__3017\
        );

    \I__333\ : Span12Mux_s10_h
    port map (
            O => \N__3017\,
            I => \N__3014\
        );

    \I__332\ : Span12Mux_h
    port map (
            O => \N__3014\,
            I => \N__3011\
        );

    \I__331\ : Odrv12
    port map (
            O => \N__3011\,
            I => \CMA_c_7\
        );

    \I__330\ : InMux
    port map (
            O => \N__3008\,
            I => \N__3005\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__3005\,
            I => \N__3002\
        );

    \I__328\ : Span4Mux_v
    port map (
            O => \N__3002\,
            I => \N__2999\
        );

    \I__327\ : Sp12to4
    port map (
            O => \N__2999\,
            I => \N__2996\
        );

    \I__326\ : Odrv12
    port map (
            O => \N__2996\,
            I => \A_c_13\
        );

    \I__325\ : CascadeMux
    port map (
            O => \N__2993\,
            I => \N__2990\
        );

    \I__324\ : InMux
    port map (
            O => \N__2990\,
            I => \N__2987\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2987\,
            I => \N__2984\
        );

    \I__322\ : Span12Mux_v
    port map (
            O => \N__2984\,
            I => \N__2981\
        );

    \I__321\ : Odrv12
    port map (
            O => \N__2981\,
            I => \A_c_6\
        );

    \I__320\ : IoInMux
    port map (
            O => \N__2978\,
            I => \N__2975\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2975\,
            I => \N__2972\
        );

    \I__318\ : Span4Mux_s1_h
    port map (
            O => \N__2972\,
            I => \N__2969\
        );

    \I__317\ : Sp12to4
    port map (
            O => \N__2969\,
            I => \N__2966\
        );

    \I__316\ : Span12Mux_s11_v
    port map (
            O => \N__2966\,
            I => \N__2963\
        );

    \I__315\ : Span12Mux_h
    port map (
            O => \N__2963\,
            I => \N__2960\
        );

    \I__314\ : Odrv12
    port map (
            O => \N__2960\,
            I => \CMA_c_4\
        );

    \I__313\ : InMux
    port map (
            O => \N__2957\,
            I => \N__2954\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2954\,
            I => \N__2951\
        );

    \I__311\ : Span4Mux_v
    port map (
            O => \N__2951\,
            I => \N__2948\
        );

    \I__310\ : Sp12to4
    port map (
            O => \N__2948\,
            I => \N__2945\
        );

    \I__309\ : Odrv12
    port map (
            O => \N__2945\,
            I => \A_c_11\
        );

    \I__308\ : CascadeMux
    port map (
            O => \N__2942\,
            I => \N__2939\
        );

    \I__307\ : InMux
    port map (
            O => \N__2939\,
            I => \N__2936\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2936\,
            I => \N__2933\
        );

    \I__305\ : Span12Mux_v
    port map (
            O => \N__2933\,
            I => \N__2930\
        );

    \I__304\ : Odrv12
    port map (
            O => \N__2930\,
            I => \A_c_4\
        );

    \I__303\ : IoInMux
    port map (
            O => \N__2927\,
            I => \N__2924\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2924\,
            I => \N__2921\
        );

    \I__301\ : Span4Mux_s1_v
    port map (
            O => \N__2921\,
            I => \N__2918\
        );

    \I__300\ : Sp12to4
    port map (
            O => \N__2918\,
            I => \N__2915\
        );

    \I__299\ : Span12Mux_h
    port map (
            O => \N__2915\,
            I => \N__2912\
        );

    \I__298\ : Span12Mux_v
    port map (
            O => \N__2912\,
            I => \N__2909\
        );

    \I__297\ : Odrv12
    port map (
            O => \N__2909\,
            I => \CMA_c_2\
        );

    \I__296\ : IoInMux
    port map (
            O => \N__2906\,
            I => \N__2903\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2903\,
            I => \N__2900\
        );

    \I__294\ : Span12Mux_s9_h
    port map (
            O => \N__2900\,
            I => \N__2897\
        );

    \I__293\ : Odrv12
    port map (
            O => \N__2897\,
            I => \CLK40_OUT_i_i\
        );

    \I__292\ : IoInMux
    port map (
            O => \N__2894\,
            I => \N__2891\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2891\,
            I => \N__2888\
        );

    \I__290\ : Span4Mux_s3_h
    port map (
            O => \N__2888\,
            I => \N__2885\
        );

    \I__289\ : Span4Mux_h
    port map (
            O => \N__2885\,
            I => \N__2882\
        );

    \I__288\ : Span4Mux_v
    port map (
            O => \N__2882\,
            I => \N__2879\
        );

    \I__287\ : Span4Mux_v
    port map (
            O => \N__2879\,
            I => \N__2875\
        );

    \I__286\ : InMux
    port map (
            O => \N__2878\,
            I => \N__2872\
        );

    \I__285\ : Odrv4
    port map (
            O => \N__2875\,
            I => \TACK_OUTn\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2872\,
            I => \TACK_OUTn\
        );

    \I__283\ : IoInMux
    port map (
            O => \N__2867\,
            I => \N__2864\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2864\,
            I => \N__2861\
        );

    \I__281\ : Span4Mux_s2_v
    port map (
            O => \N__2861\,
            I => \N__2858\
        );

    \I__280\ : Span4Mux_v
    port map (
            O => \N__2858\,
            I => \N__2855\
        );

    \I__279\ : Odrv4
    port map (
            O => \N__2855\,
            I => \CLK80_OUT_i_i\
        );

    \I__278\ : IoInMux
    port map (
            O => \N__2852\,
            I => \N__2849\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2849\,
            I => \N__2846\
        );

    \I__276\ : Span4Mux_s2_h
    port map (
            O => \N__2846\,
            I => \N__2843\
        );

    \I__275\ : Span4Mux_v
    port map (
            O => \N__2843\,
            I => \N__2840\
        );

    \I__274\ : Odrv4
    port map (
            O => \N__2840\,
            I => \N_620_i\
        );

    \I__273\ : InMux
    port map (
            O => \N__2837\,
            I => \N__2834\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2834\,
            I => \N__2831\
        );

    \I__271\ : Span4Mux_v
    port map (
            O => \N__2831\,
            I => \N__2828\
        );

    \I__270\ : Sp12to4
    port map (
            O => \N__2828\,
            I => \N__2825\
        );

    \I__269\ : Odrv12
    port map (
            O => \N__2825\,
            I => \A_c_9\
        );

    \I__268\ : CascadeMux
    port map (
            O => \N__2822\,
            I => \N__2819\
        );

    \I__267\ : InMux
    port map (
            O => \N__2819\,
            I => \N__2816\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2816\,
            I => \N__2813\
        );

    \I__265\ : Span4Mux_v
    port map (
            O => \N__2813\,
            I => \N__2810\
        );

    \I__264\ : Sp12to4
    port map (
            O => \N__2810\,
            I => \N__2807\
        );

    \I__263\ : Span12Mux_h
    port map (
            O => \N__2807\,
            I => \N__2804\
        );

    \I__262\ : Span12Mux_v
    port map (
            O => \N__2804\,
            I => \N__2801\
        );

    \I__261\ : Odrv12
    port map (
            O => \N__2801\,
            I => \A_c_2\
        );

    \I__260\ : IoInMux
    port map (
            O => \N__2798\,
            I => \N__2795\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__2795\,
            I => \N__2792\
        );

    \I__258\ : Span4Mux_s1_v
    port map (
            O => \N__2792\,
            I => \N__2789\
        );

    \I__257\ : Sp12to4
    port map (
            O => \N__2789\,
            I => \N__2786\
        );

    \I__256\ : Span12Mux_h
    port map (
            O => \N__2786\,
            I => \N__2783\
        );

    \I__255\ : Odrv12
    port map (
            O => \N__2783\,
            I => \CMA_c_0\
        );

    \I__254\ : InMux
    port map (
            O => \N__2780\,
            I => \N__2777\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__2777\,
            I => \N__2774\
        );

    \I__252\ : Span4Mux_v
    port map (
            O => \N__2774\,
            I => \N__2771\
        );

    \I__251\ : Sp12to4
    port map (
            O => \N__2771\,
            I => \N__2768\
        );

    \I__250\ : Odrv12
    port map (
            O => \N__2768\,
            I => \A_c_12\
        );

    \I__249\ : InMux
    port map (
            O => \N__2765\,
            I => \N__2762\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__2762\,
            I => \N__2759\
        );

    \I__247\ : Span4Mux_v
    port map (
            O => \N__2759\,
            I => \N__2756\
        );

    \I__246\ : Span4Mux_v
    port map (
            O => \N__2756\,
            I => \N__2753\
        );

    \I__245\ : Sp12to4
    port map (
            O => \N__2753\,
            I => \N__2750\
        );

    \I__244\ : Odrv12
    port map (
            O => \N__2750\,
            I => \A_c_5\
        );

    \I__243\ : IoInMux
    port map (
            O => \N__2747\,
            I => \N__2744\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__2744\,
            I => \N__2741\
        );

    \I__241\ : Span12Mux_s6_h
    port map (
            O => \N__2741\,
            I => \N__2738\
        );

    \I__240\ : Span12Mux_h
    port map (
            O => \N__2738\,
            I => \N__2735\
        );

    \I__239\ : Span12Mux_v
    port map (
            O => \N__2735\,
            I => \N__2732\
        );

    \I__238\ : Odrv12
    port map (
            O => \N__2732\,
            I => \CMA_c_3\
        );

    \I__237\ : IoInMux
    port map (
            O => \N__2729\,
            I => \N__2726\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2726\,
            I => \N__2723\
        );

    \I__235\ : Span4Mux_s0_v
    port map (
            O => \N__2723\,
            I => \N__2720\
        );

    \I__234\ : Span4Mux_v
    port map (
            O => \N__2720\,
            I => \N__2717\
        );

    \I__233\ : Sp12to4
    port map (
            O => \N__2717\,
            I => \N__2714\
        );

    \I__232\ : Span12Mux_h
    port map (
            O => \N__2714\,
            I => \N__2711\
        );

    \I__231\ : Span12Mux_v
    port map (
            O => \N__2711\,
            I => \N__2708\
        );

    \I__230\ : Odrv12
    port map (
            O => \N__2708\,
            I => \CLK40_IN_c\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5119\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6884\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6038\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3332\,
            lcout => \N_620_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__2837\,
            in1 => \N__4710\,
            in2 => \N__2822\,
            in3 => \N__6375\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6024\,
            ce => \N__4572\,
            sr => \N__7086\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__6374\,
            in1 => \N__2780\,
            in2 => \N__4720\,
            in3 => \N__2765\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6024\,
            ce => \N__4572\,
            sr => \N__7086\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__3107\,
            in1 => \N__6379\,
            in2 => \N__3089\,
            in3 => \N__4707\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6011\,
            ce => \N__4577\,
            sr => \N__7088\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__6378\,
            in1 => \N__3053\,
            in2 => \N__4719\,
            in3 => \N__3041\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6011\,
            ce => \N__4577\,
            sr => \N__7088\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__3008\,
            in1 => \N__6364\,
            in2 => \N__2993\,
            in3 => \N__4718\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6013\,
            ce => \N__4576\,
            sr => \N__7087\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__2957\,
            in1 => \N__6376\,
            in2 => \N__2942\,
            in3 => \N__4714\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6019\,
            ce => \N__4560\,
            sr => \N__7085\
        );

    \CLK40C_obuf_RNO_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3175\,
            lcout => \CLK40_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3188\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6030\,
            ce => 'H',
            sr => \N__7072\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3215\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6032\,
            ce => 'H',
            sr => \N__7069\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111000100"
        )
    port map (
            in0 => \N__3125\,
            in1 => \N__2878\,
            in2 => \N__3176\,
            in3 => \N__3214\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6032\,
            ce => 'H',
            sr => \N__7069\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3484\,
            in2 => \_gnd_net_\,
            in3 => \N__3499\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__3547\,
            in1 => \N__3241\,
            in2 => \N__3518\,
            in3 => \N__3256\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111111011"
        )
    port map (
            in0 => \N__3532\,
            in1 => \N__3227\,
            in2 => \N__3467\,
            in3 => \N__3221\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6025\,
            ce => 'H',
            sr => \N__7073\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3213\,
            in2 => \_gnd_net_\,
            in3 => \N__3187\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6809\,
            in2 => \_gnd_net_\,
            in3 => \N__3598\,
            lcout => \U712_REG_SM.STATE_COUNT5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__3560\,
            in1 => \N__6656\,
            in2 => \N__4399\,
            in3 => \N__3200\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6031\,
            ce => 'H',
            sr => \N__7066\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__3194\,
            in1 => \N__3369\,
            in2 => \N__3395\,
            in3 => \N__3122\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6031\,
            ce => 'H',
            sr => \N__7066\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__3123\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3171\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6031\,
            ce => 'H',
            sr => \N__7066\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000110000"
        )
    port map (
            in0 => \N__3170\,
            in1 => \N__3370\,
            in2 => \N__3356\,
            in3 => \N__3124\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6031\,
            ce => 'H',
            sr => \N__7066\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3613\,
            in2 => \_gnd_net_\,
            in3 => \N__3628\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__6970\,
            in1 => \N__3388\,
            in2 => \N__3377\,
            in3 => \N__3348\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_45_0_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__7120\,
            in1 => \_gnd_net_\,
            in2 => \N__3374\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.N_45_0_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__6971\,
            in1 => \N__3371\,
            in2 => \_gnd_net_\,
            in3 => \N__3355\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6034\,
            ce => \N__3320\,
            sr => \N__7055\
        );

    \U712_BUFFERS.un2_VBENn_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6773\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3439\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__3296\,
            in1 => \N__6328\,
            in2 => \_gnd_net_\,
            in3 => \N__4677\,
            lcout => \U712_CHIP_RAM.A_m_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__3275\,
            in1 => \N__6318\,
            in2 => \_gnd_net_\,
            in3 => \N__4661\,
            lcout => \U712_CHIP_RAM.A_m_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3257\,
            in2 => \_gnd_net_\,
            in3 => \N__3245\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__3452\,
            ce => 'H',
            sr => \N__3677\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3242\,
            in2 => \_gnd_net_\,
            in3 => \N__3230\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__3452\,
            ce => 'H',
            sr => \N__3677\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3548\,
            in2 => \_gnd_net_\,
            in3 => \N__3536\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__3452\,
            ce => 'H',
            sr => \N__3677\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3533\,
            in2 => \_gnd_net_\,
            in3 => \N__3521\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__3452\,
            ce => 'H',
            sr => \N__3677\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3517\,
            in2 => \_gnd_net_\,
            in3 => \N__3503\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__3452\,
            ce => 'H',
            sr => \N__3677\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3500\,
            in2 => \_gnd_net_\,
            in3 => \N__3488\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__3452\,
            ce => 'H',
            sr => \N__3677\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3485\,
            in2 => \_gnd_net_\,
            in3 => \N__3473\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__3452\,
            ce => 'H',
            sr => \N__3677\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3466\,
            in2 => \_gnd_net_\,
            in3 => \N__3470\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3452\,
            ce => 'H',
            sr => \N__3677\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIEJEJ2_1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5368\,
            in1 => \N__5886\,
            in2 => \N__5647\,
            in3 => \N__3875\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIDQ7S6_1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__3953\,
            in1 => \N__4365\,
            in2 => \N__3443\,
            in3 => \N__5290\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100000011"
        )
    port map (
            in0 => \N__3812\,
            in1 => \N__3602\,
            in2 => \N__3440\,
            in3 => \N__3947\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6022\,
            ce => 'H',
            sr => \N__7070\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3659\,
            in2 => \_gnd_net_\,
            in3 => \N__3810\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6026\,
            ce => 'H',
            sr => \N__7067\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4235\,
            in2 => \_gnd_net_\,
            in3 => \N__5703\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6026\,
            ce => 'H',
            sr => \N__7067\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4213\,
            lcout => \U712_REG_SM_DBR_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6026\,
            ce => 'H',
            sr => \N__7067\
        );

    \U712_CHIP_RAM.DBR_SYNC_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3653\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM_DBR_SYNC_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6026\,
            ce => 'H',
            sr => \N__7067\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__4052\,
            in1 => \N__4070\,
            in2 => \N__3632\,
            in3 => \N__4046\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6028\,
            ce => 'H',
            sr => \N__7059\
        );

    \U712_REG_SM.REG_TACK_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000011111011"
        )
    port map (
            in0 => \N__6156\,
            in1 => \N__3994\,
            in2 => \N__3617\,
            in3 => \N__4028\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6028\,
            ce => 'H',
            sr => \N__7059\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__3591\,
            in1 => \N__3559\,
            in2 => \N__6821\,
            in3 => \N__4163\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6028\,
            ce => 'H',
            sr => \N__7059\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__5039\,
            in1 => \N__5006\,
            in2 => \N__3995\,
            in3 => \N__4412\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6028\,
            ce => 'H',
            sr => \N__7059\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001011111010"
        )
    port map (
            in0 => \N__4037\,
            in1 => \N__6125\,
            in2 => \N__6161\,
            in3 => \N__6091\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6028\,
            ce => 'H',
            sr => \N__7059\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_4_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101010101"
        )
    port map (
            in0 => \N__4011\,
            in1 => \N__4187\,
            in2 => \N__4217\,
            in3 => \N__5455\,
            lcout => \U712_REG_SM.N_160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_0_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000011010"
        )
    port map (
            in0 => \N__6559\,
            in1 => \N__4840\,
            in2 => \N__4820\,
            in3 => \N__6609\,
            lcout => \CLLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001010001"
        )
    port map (
            in0 => \N__3767\,
            in1 => \N__5503\,
            in2 => \N__4958\,
            in3 => \N__5459\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6033\,
            ce => 'H',
            sr => \N__7050\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011101111"
        )
    port map (
            in0 => \N__3761\,
            in1 => \N__3755\,
            in2 => \N__6365\,
            in3 => \N__6225\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6007\,
            ce => \N__4553\,
            sr => \N__7080\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011101111"
        )
    port map (
            in0 => \N__3716\,
            in1 => \N__3710\,
            in2 => \N__6358\,
            in3 => \N__6224\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6012\,
            ce => \N__4551\,
            sr => \N__7078\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6292\,
            in1 => \N__4645\,
            in2 => \N__6217\,
            in3 => \N__6413\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011000101"
        )
    port map (
            in0 => \N__4286\,
            in1 => \N__4646\,
            in2 => \N__3836\,
            in3 => \N__3851\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6014\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__4271\,
            in1 => \N__3835\,
            in2 => \N__6327\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6014\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISSMN4_2_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6967\,
            in1 => \N__5630\,
            in2 => \N__5888\,
            in3 => \N__3970\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_80_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIUTL6G_2_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__3668\,
            in1 => \N__6969\,
            in2 => \N__3662\,
            in3 => \N__4228\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000001"
        )
    port map (
            in0 => \N__4295\,
            in1 => \N__3844\,
            in2 => \N__3857\,
            in3 => \N__6216\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI5DTJ_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__3935\,
            in1 => \N__3908\,
            in2 => \_gnd_net_\,
            in3 => \N__5352\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_2\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__5884\,
            in1 => \N__6736\,
            in2 => \N__3854\,
            in3 => \N__4376\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIT4P84_0_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__3971\,
            in1 => \N__6968\,
            in2 => \_gnd_net_\,
            in3 => \N__5883\,
            lcout => \U712_CHIP_RAM.N_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110100000001"
        )
    port map (
            in0 => \N__3845\,
            in1 => \N__3831\,
            in2 => \N__4244\,
            in3 => \N__6420\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4371\,
            in1 => \N__3788\,
            in2 => \_gnd_net_\,
            in3 => \N__3877\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__3811\,
            in1 => \N__3794\,
            in2 => \N__3815\,
            in3 => \N__3980\,
            lcout => \U712_CHIP_RAM.CPU_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6020\,
            ce => 'H',
            sr => \N__7068\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNO_1_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__4063\,
            in1 => \N__5871\,
            in2 => \N__5646\,
            in3 => \N__3878\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_4_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5361\,
            in1 => \N__5411\,
            in2 => \N__5218\,
            in3 => \N__5281\,
            lcout => \U712_CHIP_RAM.N_110\,
            ltout => \U712_CHIP_RAM.N_110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3904\,
            in2 => \N__3983\,
            in3 => \N__3933\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLE_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5360\,
            in1 => \N__5784\,
            in2 => \N__5217\,
            in3 => \N__5280\,
            lcout => \U712_CHIP_RAM.N_58\,
            ltout => \U712_CHIP_RAM.N_58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIA5V93_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__5699\,
            in1 => \N__3903\,
            in2 => \N__3974\,
            in3 => \N__3932\,
            lcout => \U712_CHIP_RAM.N_118\,
            ltout => \U712_CHIP_RAM.N_118_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__3934\,
            in1 => \N__5887\,
            in2 => \N__3962\,
            in3 => \N__3959\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6020\,
            ce => 'H',
            sr => \N__7068\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__3902\,
            in1 => \N__6966\,
            in2 => \N__5729\,
            in3 => \N__3931\,
            lcout => \U712_CHIP_RAM.N_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIU1NR1_3_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__5201\,
            in1 => \N__5781\,
            in2 => \N__5639\,
            in3 => \N__5354\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_o2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIKEL61_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4208\,
            in1 => \N__4182\,
            in2 => \_gnd_net_\,
            in3 => \N__3946\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__3930\,
            in1 => \N__3901\,
            in2 => \_gnd_net_\,
            in3 => \N__5717\,
            lcout => \U712_CHIP_RAM.N_40\,
            ltout => \U712_CHIP_RAM.N_40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIC55U3_2_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001101"
        )
    port map (
            in0 => \N__5629\,
            in1 => \N__4076\,
            in2 => \N__3881\,
            in3 => \N__3876\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_10_u_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINN5O1_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111001110"
        )
    port map (
            in0 => \N__5625\,
            in1 => \N__5782\,
            in2 => \N__5727\,
            in3 => \N__5852\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_10_u_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4307\,
            in1 => \N__4337\,
            in2 => \_gnd_net_\,
            in3 => \N__5299\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5202\,
            in1 => \N__5783\,
            in2 => \N__5300\,
            in3 => \N__4064\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__5648\,
            in1 => \N__5873\,
            in2 => \_gnd_net_\,
            in3 => \N__5369\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_6_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4882\,
            in1 => \N__4936\,
            in2 => \N__5084\,
            in3 => \N__5063\,
            lcout => \U712_REG_SM.N_148_0\,
            ltout => \U712_REG_SM.N_148_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI1VLC2_5_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4021\,
            in1 => \N__5037\,
            in2 => \N__4040\,
            in3 => \N__4998\,
            lcout => \U712_REG_SM.N_157_0\,
            ltout => \U712_REG_SM.N_157_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100001111"
        )
    port map (
            in0 => \N__4012\,
            in1 => \_gnd_net_\,
            in2 => \N__4031\,
            in3 => \N__6722\,
            lcout => \U712_REG_SM.REG_TACK_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIFFKI2_5_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__4022\,
            in1 => \N__4013\,
            in2 => \N__4950\,
            in3 => \N__5499\,
            lcout => \U712_REG_SM.un1_STATE_COUNT_3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4209\,
            in1 => \N__4186\,
            in2 => \_gnd_net_\,
            in3 => \N__4937\,
            lcout => \U712_REG_SM.STATE_COUNT_srsts_i_a3_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5082\,
            in2 => \_gnd_net_\,
            in3 => \N__4883\,
            lcout => \U712_REG_SM.N_146_0\,
            ltout => \U712_REG_SM.N_146_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6151\,
            in2 => \N__4166\,
            in3 => \N__6114\,
            lcout => \U712_REG_SM.DS_EN_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI1FQR1_2_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5038\,
            in1 => \N__4996\,
            in2 => \_gnd_net_\,
            in3 => \N__5045\,
            lcout => \U712_REG_SM.N_149_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_2_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4997\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6029\,
            ce => 'H',
            sr => \N__7051\
        );

    \U712_REG_SM.C3_SYNC_1_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4886\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6029\,
            ce => 'H',
            sr => \N__7051\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4157\,
            in1 => \N__6380\,
            in2 => \_gnd_net_\,
            in3 => \N__4708\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6004\,
            ce => \N__4570\,
            sr => \N__7083\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4124\,
            in1 => \N__6363\,
            in2 => \_gnd_net_\,
            in3 => \N__4700\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6006\,
            ce => \N__4552\,
            sr => \N__7081\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7121\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4082\,
            lcout => \U712_CHIP_RAM.un1_CMA21_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100111"
        )
    port map (
            in0 => \N__6296\,
            in1 => \N__6204\,
            in2 => \N__4676\,
            in3 => \N__6414\,
            lcout => \U712_CHIP_RAM.un1_CMA21_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__4313\,
            in1 => \N__4285\,
            in2 => \N__5429\,
            in3 => \N__5363\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_29_i_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISUCO3_4_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6959\,
            in1 => \N__5219\,
            in2 => \N__5410\,
            in3 => \N__5282\,
            lcout => \U712_CHIP_RAM.N_116\,
            ltout => \U712_CHIP_RAM.N_116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINFP34_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4289\,
            in3 => \N__5730\,
            lcout => \U712_CHIP_RAM.N_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001100"
        )
    port map (
            in0 => \N__5362\,
            in1 => \N__4263\,
            in2 => \N__5735\,
            in3 => \N__5425\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_67_i_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__4333\,
            in1 => \N__4375\,
            in2 => \N__4274\,
            in3 => \N__5885\,
            lcout => \U712_CHIP_RAM.N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__5734\,
            in1 => \N__4264\,
            in2 => \_gnd_net_\,
            in3 => \N__5424\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__4332\,
            in1 => \N__4265\,
            in2 => \N__4247\,
            in3 => \N__4367\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4466\,
            in2 => \_gnd_net_\,
            in3 => \N__5240\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5215\,
            in1 => \N__5156\,
            in2 => \_gnd_net_\,
            in3 => \N__7119\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4366\,
            in1 => \N__4331\,
            in2 => \_gnd_net_\,
            in3 => \N__5859\,
            lcout => \U712_CHIP_RAM.N_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4478\,
            in1 => \N__5387\,
            in2 => \_gnd_net_\,
            in3 => \N__5638\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5367\,
            in1 => \N__5860\,
            in2 => \_gnd_net_\,
            in3 => \N__4477\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5899\,
            in1 => \N__5913\,
            in2 => \_gnd_net_\,
            in3 => \N__5136\,
            lcout => \U712_CHIP_RAM.N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5619\,
            in1 => \N__5850\,
            in2 => \N__5786\,
            in3 => \N__5200\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIMKLS1_3_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__6958\,
            in1 => \N__5773\,
            in2 => \N__5216\,
            in3 => \N__5617\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_a5_0_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIERVM2_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5704\,
            in2 => \N__4301\,
            in3 => \N__5848\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_a5_0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011010100000"
        )
    port map (
            in0 => \N__5851\,
            in1 => \N__5409\,
            in2 => \N__5246\,
            in3 => \N__4487\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__5242\,
            in1 => \N__7117\,
            in2 => \N__4298\,
            in3 => \N__5558\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6021\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAKMO6_2_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__7118\,
            in1 => \N__4486\,
            in2 => \_gnd_net_\,
            in3 => \N__5241\,
            lcout => \U712_CHIP_RAM.N_13\,
            ltout => \U712_CHIP_RAM.N_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__5778\,
            in1 => \_gnd_net_\,
            in2 => \N__4469\,
            in3 => \N__5378\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6021\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNINN5O1_0_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5849\,
            in1 => \N__5774\,
            in2 => \N__5726\,
            in3 => \N__5618\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNICU4F1_1_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4991\,
            in1 => \N__5066\,
            in2 => \N__4951\,
            in3 => \N__5035\,
            lcout => \U712_REG_SM.N_182\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__4946\,
            in1 => \N__6723\,
            in2 => \_gnd_net_\,
            in3 => \N__4885\,
            lcout => \U712_REG_SM.DS_EN_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_23_i_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011100000"
        )
    port map (
            in0 => \N__4858\,
            in1 => \N__6632\,
            in2 => \N__6587\,
            in3 => \N__4811\,
            lcout => \N_23_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_0_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111000000"
        )
    port map (
            in0 => \N__6633\,
            in1 => \N__4859\,
            in2 => \N__4819\,
            in3 => \N__6586\,
            lcout => \CUMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4411\,
            in1 => \N__5034\,
            in2 => \N__5002\,
            in3 => \N__4400\,
            lcout => \U712_REG_SM.N_155_0\,
            ltout => \U712_REG_SM.N_155_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIVQBP4_6_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__6090\,
            in1 => \N__6152\,
            in2 => \N__4379\,
            in3 => \N__6113\,
            lcout => \U712_REG_SM.STATE_COUNT_RNIVQBP4Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_1_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4945\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6027\,
            ce => 'H',
            sr => \N__7046\
        );

    \U712_REG_SM.C1_SYNC_2_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5065\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6027\,
            ce => 'H',
            sr => \N__7046\
        );

    \U712_REG_SM.C1_SYNC_0_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5120\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6027\,
            ce => 'H',
            sr => \N__7046\
        );

    \U712_REG_SM.C1_SYNC_RNIOEF21_2_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5083\,
            in1 => \N__4884\,
            in2 => \_gnd_net_\,
            in3 => \N__5064\,
            lcout => \U712_REG_SM.N_145_0\,
            ltout => \U712_REG_SM.N_145_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5036\,
            in1 => \N__4995\,
            in2 => \N__4961\,
            in3 => \N__4944\,
            lcout => \U712_REG_SM.N_152_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4904\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6027\,
            ce => 'H',
            sr => \N__7046\
        );

    \U712_BYTE_ENABLE.N_22_i_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110110000"
        )
    port map (
            in0 => \N__6631\,
            in1 => \N__4852\,
            in2 => \N__4818\,
            in3 => \N__6581\,
            lcout => \N_22_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4709\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6003\,
            ce => 'H',
            sr => \N__7082\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6362\,
            in1 => \N__6226\,
            in2 => \N__4721\,
            in3 => \N__6436\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6005\,
            ce => \N__4571\,
            sr => \N__7079\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5283\,
            in1 => \N__5435\,
            in2 => \_gnd_net_\,
            in3 => \N__5356\,
            lcout => \U712_CHIP_RAM.N_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIS6PC1_3_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5846\,
            in1 => \N__5779\,
            in2 => \_gnd_net_\,
            in3 => \N__5620\,
            lcout => \U712_CHIP_RAM.N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5355\,
            in2 => \_gnd_net_\,
            in3 => \N__5847\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_ac0_1_out\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_ac0_1_out_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5381\,
            in3 => \N__5621\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_ac0_3_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_ac0_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__5780\,
            in1 => \_gnd_net_\,
            in2 => \N__5372\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI85LA2_4_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5353\,
            in1 => \N__5203\,
            in2 => \_gnd_net_\,
            in3 => \N__5279\,
            lcout => \U712_CHIP_RAM.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5204\,
            in1 => \N__5154\,
            in2 => \_gnd_net_\,
            in3 => \N__5137\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_c6\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_11_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__7115\,
            in1 => \_gnd_net_\,
            in2 => \N__5222\,
            in3 => \N__5914\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__5205\,
            in1 => \N__5155\,
            in2 => \N__5141\,
            in3 => \N__7114\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__7116\,
            in1 => \N__5900\,
            in2 => \N__5924\,
            in3 => \N__5915\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011111111111"
        )
    port map (
            in0 => \N__5872\,
            in1 => \N__5785\,
            in2 => \N__5728\,
            in3 => \N__5637\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER19_i_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_1_ess_RNO_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7113\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5521\,
            lcout => \U712_REG_SM.N_177_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIURLC2_2_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5536\,
            in2 => \_gnd_net_\,
            in3 => \N__5551\,
            lcout => \U712_REG_SM.N_156_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__5540\,
            in1 => \N__6653\,
            in2 => \_gnd_net_\,
            in3 => \N__5552\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6023\,
            ce => 'H',
            sr => \N__7045\
        );

    \U712_REG_SM.LDS_OUT_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110001010"
        )
    port map (
            in0 => \N__6655\,
            in1 => \N__6634\,
            in2 => \N__6535\,
            in3 => \N__6520\,
            lcout => \U712_REG_SM.LDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6023\,
            ce => 'H',
            sr => \N__7045\
        );

    \U712_REG_SM.DS_EN_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010011111110"
        )
    port map (
            in0 => \N__5468\,
            in1 => \N__6468\,
            in2 => \N__5525\,
            in3 => \N__5510\,
            lcout => \U712_REG_SM.DS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6023\,
            ce => 'H',
            sr => \N__7045\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111100101010"
        )
    port map (
            in0 => \N__5454\,
            in1 => \N__5504\,
            in2 => \N__5483\,
            in3 => \N__5467\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6023\,
            ce => 'H',
            sr => \N__7045\
        );

    \U712_REG_SM.UDS_OUT_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100101010"
        )
    port map (
            in0 => \N__6654\,
            in1 => \N__6635\,
            in2 => \N__6536\,
            in3 => \N__6484\,
            lcout => \U712_REG_SM.UDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6023\,
            ce => 'H',
            sr => \N__7045\
        );

    \U712_REG_SM.LDS_OUT_2_0_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6582\,
            in2 => \_gnd_net_\,
            in3 => \N__6718\,
            lcout => \U712_REG_SM.LDS_OUT_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDS_OUT_RNIL31J_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6521\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6469\,
            lcout => \U712_REG_SM_un1_LDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_RNIUP9B_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6488\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6473\,
            lcout => \U712_REG_SM_un1_UDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CRCSn_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6437\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6000\,
            ce => 'H',
            sr => \N__7084\
        );

    \U712_CHIP_RAM.RASn_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6377\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6001\,
            ce => 'H',
            sr => \N__7077\
        );

    \U712_CHIP_RAM.CASn_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6227\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6002\,
            ce => 'H',
            sr => \N__7071\
        );

    \U712_REG_SM.REGENn_1_ess_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6160\,
            in1 => \N__6121\,
            in2 => \_gnd_net_\,
            in3 => \N__6095\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6015\,
            ce => \N__5930\,
            sr => \N__7044\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6947\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_13_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDDIR_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6820\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6737\,
            lcout => \DRDDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 9 2025 19:17:52

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    DBRn : in std_logic;
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__12127\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \DBRn_c_i_cascade_\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \U712_CYCLE_TERM_TCIn_0_i\ : std_logic;
signal \U712_CYCLE_TERM.RAM_CYCLEZ0\ : std_logic;
signal \U712_REG_SM.N_486_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_6_0_a3_0_a2_1\ : std_logic;
signal \N_490\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_554_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_a2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_373\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0\ : std_logic;
signal \U712_CHIP_RAM.N_409\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1\ : std_logic;
signal \U712_CYCLE_TERM.N_565\ : std_logic;
signal \U712_CYCLE_TERM.N_407\ : std_logic;
signal \U712_CYCLE_TERM.N_534\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.N_371_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_375_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_498\ : std_logic;
signal \U712_CHIP_RAM.N_547_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_501_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_a2_0_cascade_\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.N_666_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_393_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_6_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0_cascade_\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\ : std_logic;
signal \U712_CHIP_RAM.N_504\ : std_logic;
signal \U712_CYCLE_TERM.N_539_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \A_c_14\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.N_669_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_520_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_560\ : std_logic;
signal \U712_CHIP_RAM.N_501\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1\ : std_logic;
signal \U712_CHIP_RAM.N_515\ : std_logic;
signal \U712_CHIP_RAM.N_516\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_519\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_78\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_559_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_665\ : std_logic;
signal \U712_CHIP_RAM.N_665_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_471\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.N_506_cascade_\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \U712_CHIP_RAM.N_375\ : std_logic;
signal \U712_CHIP_RAM.N_547\ : std_logic;
signal \U712_CHIP_RAM.N_522\ : std_logic;
signal \U712_CHIP_RAM.N_523_cascade_\ : std_logic;
signal \U712_CHIP_RAM.BANK0_9\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.N_545_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_549\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_666\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_557\ : std_logic;
signal \U712_CHIP_RAM.N_393\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_557_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_31\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_566\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \ASn_c\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_1\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_REG_SM.N_447\ : std_logic;
signal \U712_REG_SM.N_447_cascade_\ : std_logic;
signal \U712_REG_SM.REG_TACK_RNOZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_478\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.N_379_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.N_517\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_a2_1_0\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_567\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_562\ : std_logic;
signal \U712_CHIP_RAM.N_502\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_545\ : std_logic;
signal \U712_CHIP_RAM.N_572\ : std_logic;
signal \U712_CHIP_RAM.N_518_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_a2_0_0\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \U712_CHIP_RAM.N_492_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_0_0_a2_0_0_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_374\ : std_logic;
signal \U712_REG_SM.N_374_cascade_\ : std_logic;
signal \U712_REG_SM.N_417\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.DS_EN_RNOZ0Z_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \RASn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_8\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_REG_SM.N_477_cascade_\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.N_422\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.N_445\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.START_RSTZ0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN_RNOZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.un13_0\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \U712_REG_SM.N_661\ : std_logic;
signal \U712_REG_SM.N_389\ : std_logic;
signal \U712_REG_SM.N_475_cascade_\ : std_logic;
signal \N_57_i\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_449_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.START_RST_0_sqmuxa\ : std_logic;
signal \U712_REG_SM.N_396_cascade_\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_4_i_i_0_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_2\ : std_logic;
signal \U712_REG_SM.N_479\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \U712_CHIP_RAM.un3_DMA_CYCLE_START\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \N_295_i\ : std_logic;
signal \N_299_i\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \N_297_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_528\ : std_logic;
signal \U712_BYTE_ENABLE.N_377_cascade_\ : std_logic;
signal \U712_BYTE_ENABLE.N_508\ : std_logic;
signal \U712_BYTE_ENABLE.N_377\ : std_logic;
signal \U712_BYTE_ENABLE.N_530\ : std_logic;
signal \U712_BYTE_ENABLE.N_532\ : std_logic;
signal \U712_BYTE_ENABLE.N_364_i\ : std_logic;
signal \DMA_LATCH_EN_c\ : std_logic;
signal \N_403_i\ : std_logic;
signal \CASn_c\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\ : std_logic;
signal \U712_CHIP_RAM.N_379\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ1Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \N_402_i\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \N_291\ : std_logic;
signal \N_400_i\ : std_logic;
signal \DS_ENm\ : std_logic;
signal \N_293\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \N_401_i\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \WRITE_CYCLEm\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \N_450\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    TBIn <= \TBIn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    TCIn <= \TCIn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4089\,
            RESETB => \N__4938\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12127\,
            DIN => \N__12126\,
            DOUT => \N__12125\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12127\,
            PADOUT => \N__12126\,
            PADIN => \N__12125\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8718\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12118\,
            DIN => \N__12117\,
            DOUT => \N__12116\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12118\,
            PADOUT => \N__12117\,
            PADIN => \N__12116\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12109\,
            DIN => \N__12108\,
            DOUT => \N__12107\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12109\,
            PADOUT => \N__12108\,
            PADIN => \N__12107\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9240\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12100\,
            DIN => \N__12099\,
            DOUT => \N__12098\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12100\,
            PADOUT => \N__12099\,
            PADIN => \N__12098\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11121\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12091\,
            DIN => \N__12090\,
            DOUT => \N__12089\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12091\,
            PADOUT => \N__12090\,
            PADIN => \N__12089\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12082\,
            DIN => \N__12081\,
            DOUT => \N__12080\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12082\,
            PADOUT => \N__12081\,
            PADIN => \N__12080\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12073\,
            DIN => \N__12072\,
            DOUT => \N__12071\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12073\,
            PADOUT => \N__12072\,
            PADIN => \N__12071\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12064\,
            DIN => \N__12063\,
            DOUT => \N__12062\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12064\,
            PADOUT => \N__12063\,
            PADIN => \N__12062\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12055\,
            DIN => \N__12054\,
            DOUT => \N__12053\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12055\,
            PADOUT => \N__12054\,
            PADIN => \N__12053\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12046\,
            DIN => \N__12045\,
            DOUT => \N__12044\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12046\,
            PADOUT => \N__12045\,
            PADIN => \N__12044\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12037\,
            DIN => \N__12036\,
            DOUT => \N__12035\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12037\,
            PADOUT => \N__12036\,
            PADIN => \N__12035\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5616\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12028\,
            DIN => \N__12027\,
            DOUT => \N__12026\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12028\,
            PADOUT => \N__12027\,
            PADIN => \N__12026\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9252\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12019\,
            DIN => \N__12018\,
            DOUT => \N__12017\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12019\,
            PADOUT => \N__12018\,
            PADIN => \N__12017\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12010\,
            DIN => \N__12009\,
            DOUT => \N__12008\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12010\,
            PADOUT => \N__12009\,
            PADIN => \N__12008\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6485\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12001\,
            DIN => \N__12000\,
            DOUT => \N__11999\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12001\,
            PADOUT => \N__12000\,
            PADIN => \N__11999\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11992\,
            DIN => \N__11991\,
            DOUT => \N__11990\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11992\,
            PADOUT => \N__11991\,
            PADIN => \N__11990\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11983\,
            DIN => \N__11982\,
            DOUT => \N__11981\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11983\,
            PADOUT => \N__11982\,
            PADIN => \N__11981\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4200\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11974\,
            DIN => \N__11973\,
            DOUT => \N__11972\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11974\,
            PADOUT => \N__11973\,
            PADIN => \N__11972\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11965\,
            DIN => \N__11964\,
            DOUT => \N__11963\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11965\,
            PADOUT => \N__11964\,
            PADIN => \N__11963\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11956\,
            DIN => \N__11955\,
            DOUT => \N__11954\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11956\,
            PADOUT => \N__11955\,
            PADIN => \N__11954\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8841\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11947\,
            DIN => \N__11946\,
            DOUT => \N__11945\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11947\,
            PADOUT => \N__11946\,
            PADIN => \N__11945\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11938\,
            DIN => \N__11937\,
            DOUT => \N__11936\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11938\,
            PADOUT => \N__11937\,
            PADIN => \N__11936\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7332\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11929\,
            DIN => \N__11928\,
            DOUT => \N__11927\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11929\,
            PADOUT => \N__11928\,
            PADIN => \N__11927\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11920\,
            DIN => \N__11919\,
            DOUT => \N__11918\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11920\,
            PADOUT => \N__11919\,
            PADIN => \N__11918\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10746\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11911\,
            DIN => \N__11910\,
            DOUT => \N__11909\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11911\,
            PADOUT => \N__11910\,
            PADIN => \N__11909\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7425\,
            DIN0 => OPEN,
            DOUT0 => \N__5292\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11902\,
            DIN => \N__11901\,
            DOUT => \N__11900\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11902\,
            PADOUT => \N__11901\,
            PADIN => \N__11900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11893\,
            DIN => \N__11892\,
            DOUT => \N__11891\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11893\,
            PADOUT => \N__11892\,
            PADIN => \N__11891\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11884\,
            DIN => \N__11883\,
            DOUT => \N__11882\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11884\,
            PADOUT => \N__11883\,
            PADIN => \N__11882\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11875\,
            DIN => \N__11874\,
            DOUT => \N__11873\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11875\,
            PADOUT => \N__11874\,
            PADIN => \N__11873\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11866\,
            DIN => \N__11865\,
            DOUT => \N__11864\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11866\,
            PADOUT => \N__11865\,
            PADIN => \N__11864\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11857\,
            DIN => \N__11856\,
            DOUT => \N__11855\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11857\,
            PADOUT => \N__11856\,
            PADIN => \N__11855\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9270\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11848\,
            DIN => \N__11847\,
            DOUT => \N__11846\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11848\,
            PADOUT => \N__11847\,
            PADIN => \N__11846\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11839\,
            DIN => \N__11838\,
            DOUT => \N__11837\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11839\,
            PADOUT => \N__11838\,
            PADIN => \N__11837\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11830\,
            DIN => \N__11829\,
            DOUT => \N__11828\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11830\,
            PADOUT => \N__11829\,
            PADIN => \N__11828\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11821\,
            DIN => \N__11820\,
            DOUT => \N__11819\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11821\,
            PADOUT => \N__11820\,
            PADIN => \N__11819\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11812\,
            DIN => \N__11811\,
            DOUT => \N__11810\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11812\,
            PADOUT => \N__11811\,
            PADIN => \N__11810\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4128\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11803\,
            DIN => \N__11802\,
            DOUT => \N__11801\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11803\,
            PADOUT => \N__11802\,
            PADIN => \N__11801\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11794\,
            DIN => \N__11793\,
            DOUT => \N__11792\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11794\,
            PADOUT => \N__11793\,
            PADIN => \N__11792\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6921\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11785\,
            DIN => \N__11784\,
            DOUT => \N__11783\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11785\,
            PADOUT => \N__11784\,
            PADIN => \N__11783\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5112\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11776\,
            DIN => \N__11775\,
            DOUT => \N__11774\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11776\,
            PADOUT => \N__11775\,
            PADIN => \N__11774\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8003\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11767\,
            DIN => \N__11766\,
            DOUT => \N__11765\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11767\,
            PADOUT => \N__11766\,
            PADIN => \N__11765\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4170\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11758\,
            DIN => \N__11757\,
            DOUT => \N__11756\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11758\,
            PADOUT => \N__11757\,
            PADIN => \N__11756\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11749\,
            DIN => \N__11748\,
            DOUT => \N__11747\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11749\,
            PADOUT => \N__11748\,
            PADIN => \N__11747\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5820\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11740\,
            DIN => \N__11739\,
            DOUT => \N__11738\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11740\,
            PADOUT => \N__11739\,
            PADIN => \N__11738\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6429\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11731\,
            DIN => \N__11730\,
            DOUT => \N__11729\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11731\,
            PADOUT => \N__11730\,
            PADIN => \N__11729\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8301\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11722\,
            DIN => \N__11721\,
            DOUT => \N__11720\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11722\,
            PADOUT => \N__11721\,
            PADIN => \N__11720\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11713\,
            DIN => \N__11712\,
            DOUT => \N__11711\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11713\,
            PADOUT => \N__11712\,
            PADIN => \N__11711\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11704\,
            DIN => \N__11703\,
            DOUT => \N__11702\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11704\,
            PADOUT => \N__11703\,
            PADIN => \N__11702\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11695\,
            DIN => \N__11694\,
            DOUT => \N__11693\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11695\,
            PADOUT => \N__11694\,
            PADIN => \N__11693\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11686\,
            DIN => \N__11685\,
            DOUT => \N__11684\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11686\,
            PADOUT => \N__11685\,
            PADIN => \N__11684\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7179\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11677\,
            DIN => \N__11676\,
            DOUT => \N__11675\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11677\,
            PADOUT => \N__11676\,
            PADIN => \N__11675\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11668\,
            DIN => \N__11667\,
            DOUT => \N__11666\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11668\,
            PADOUT => \N__11667\,
            PADIN => \N__11666\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8002\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11659\,
            DIN => \N__11658\,
            DOUT => \N__11657\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11659\,
            PADOUT => \N__11658\,
            PADIN => \N__11657\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9219\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11650\,
            DIN => \N__11649\,
            DOUT => \N__11648\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11650\,
            PADOUT => \N__11649\,
            PADIN => \N__11648\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10101\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11641\,
            DIN => \N__11640\,
            DOUT => \N__11639\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11641\,
            PADOUT => \N__11640\,
            PADIN => \N__11639\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7860\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11632\,
            DIN => \N__11631\,
            DOUT => \N__11630\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11632\,
            PADOUT => \N__11631\,
            PADIN => \N__11630\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7296\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11623\,
            DIN => \N__11622\,
            DOUT => \N__11621\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11623\,
            PADOUT => \N__11622\,
            PADIN => \N__11621\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5816\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11614\,
            DIN => \N__11613\,
            DOUT => \N__11612\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11614\,
            PADOUT => \N__11613\,
            PADIN => \N__11612\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11605\,
            DIN => \N__11604\,
            DOUT => \N__11603\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11605\,
            PADOUT => \N__11604\,
            PADIN => \N__11603\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11596\,
            DIN => \N__11595\,
            DOUT => \N__11594\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11596\,
            PADOUT => \N__11595\,
            PADIN => \N__11594\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8739\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11587\,
            DIN => \N__11586\,
            DOUT => \N__11585\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11587\,
            PADOUT => \N__11586\,
            PADIN => \N__11585\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7356\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11578\,
            DIN => \N__11577\,
            DOUT => \N__11576\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11578\,
            PADOUT => \N__11577\,
            PADIN => \N__11576\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5703\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11569\,
            DIN => \N__11568\,
            DOUT => \N__11567\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11569\,
            PADOUT => \N__11568\,
            PADIN => \N__11567\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8592\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11560\,
            DIN => \N__11559\,
            DOUT => \N__11558\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11560\,
            PADOUT => \N__11559\,
            PADIN => \N__11558\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11551\,
            DIN => \N__11550\,
            DOUT => \N__11549\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11551\,
            PADOUT => \N__11550\,
            PADIN => \N__11549\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11542\,
            DIN => \N__11541\,
            DOUT => \N__11540\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11542\,
            PADOUT => \N__11541\,
            PADIN => \N__11540\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5904\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11533\,
            DIN => \N__11532\,
            DOUT => \N__11531\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11533\,
            PADOUT => \N__11532\,
            PADIN => \N__11531\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11524\,
            DIN => \N__11523\,
            DOUT => \N__11522\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11524\,
            PADOUT => \N__11523\,
            PADIN => \N__11522\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11515\,
            DIN => \N__11514\,
            DOUT => \N__11513\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11515\,
            PADOUT => \N__11514\,
            PADIN => \N__11513\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7233\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11506\,
            DIN => \N__11505\,
            DOUT => \N__11504\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11506\,
            PADOUT => \N__11505\,
            PADIN => \N__11504\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9507\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11497\,
            DIN => \N__11496\,
            DOUT => \N__11495\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11497\,
            PADOUT => \N__11496\,
            PADIN => \N__11495\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11488\,
            DIN => \N__11487\,
            DOUT => \N__11486\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11488\,
            PADOUT => \N__11487\,
            PADIN => \N__11486\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8760\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11479\,
            DIN => \N__11478\,
            DOUT => \N__11477\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11479\,
            PADOUT => \N__11478\,
            PADIN => \N__11477\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7418\,
            DIN0 => OPEN,
            DOUT0 => \N__5291\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11470\,
            DIN => \N__11469\,
            DOUT => \N__11468\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11470\,
            PADOUT => \N__11469\,
            PADIN => \N__11468\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7158\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11461\,
            DIN => \N__11460\,
            DOUT => \N__11459\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11461\,
            PADOUT => \N__11460\,
            PADIN => \N__11459\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11452\,
            DIN => \N__11451\,
            DOUT => \N__11450\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11452\,
            PADOUT => \N__11451\,
            PADIN => \N__11450\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11443\,
            DIN => \N__11442\,
            DOUT => \N__11441\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11443\,
            PADOUT => \N__11442\,
            PADIN => \N__11441\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7257\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11434\,
            DIN => \N__11433\,
            DOUT => \N__11432\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11434\,
            PADOUT => \N__11433\,
            PADIN => \N__11432\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11425\,
            DIN => \N__11424\,
            DOUT => \N__11423\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11425\,
            PADOUT => \N__11424\,
            PADIN => \N__11423\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11416\,
            DIN => \N__11415\,
            DOUT => \N__11414\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11416\,
            PADOUT => \N__11415\,
            PADIN => \N__11414\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7587\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11407\,
            DIN => \N__11406\,
            DOUT => \N__11405\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11407\,
            PADOUT => \N__11406\,
            PADIN => \N__11405\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11398\,
            DIN => \N__11397\,
            DOUT => \N__11396\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11398\,
            PADOUT => \N__11397\,
            PADIN => \N__11396\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11389\,
            DIN => \N__11388\,
            DOUT => \N__11387\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11389\,
            PADOUT => \N__11388\,
            PADIN => \N__11387\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5646\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11380\,
            DIN => \N__11379\,
            DOUT => \N__11378\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11380\,
            PADOUT => \N__11379\,
            PADIN => \N__11378\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11109\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11371\,
            DIN => \N__11370\,
            DOUT => \N__11369\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11371\,
            PADOUT => \N__11370\,
            PADIN => \N__11369\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11091\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11362\,
            DIN => \N__11361\,
            DOUT => \N__11360\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11362\,
            PADOUT => \N__11361\,
            PADIN => \N__11360\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4443\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11353\,
            DIN => \N__11352\,
            DOUT => \N__11351\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11353\,
            PADOUT => \N__11352\,
            PADIN => \N__11351\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11344\,
            DIN => \N__11343\,
            DOUT => \N__11342\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11344\,
            PADOUT => \N__11343\,
            PADIN => \N__11342\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11335\,
            DIN => \N__11334\,
            DOUT => \N__11333\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11335\,
            PADOUT => \N__11334\,
            PADIN => \N__11333\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9060\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11326\,
            DIN => \N__11325\,
            DOUT => \N__11324\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11326\,
            PADOUT => \N__11325\,
            PADIN => \N__11324\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11317\,
            DIN => \N__11316\,
            DOUT => \N__11315\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11317\,
            PADOUT => \N__11316\,
            PADIN => \N__11315\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11308\,
            DIN => \N__11307\,
            DOUT => \N__11306\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11308\,
            PADOUT => \N__11307\,
            PADIN => \N__11306\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5427\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11299\,
            DIN => \N__11298\,
            DOUT => \N__11297\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11299\,
            PADOUT => \N__11298\,
            PADIN => \N__11297\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11043\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11290\,
            DIN => \N__11289\,
            DOUT => \N__11288\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11290\,
            PADOUT => \N__11289\,
            PADIN => \N__11288\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8004\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11281\,
            DIN => \N__11280\,
            DOUT => \N__11279\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11281\,
            PADOUT => \N__11280\,
            PADIN => \N__11279\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2749\ : CascadeMux
    port map (
            O => \N__11262\,
            I => \N__11259\
        );

    \I__2748\ : InMux
    port map (
            O => \N__11259\,
            I => \N__11256\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__11256\,
            I => \N__11252\
        );

    \I__2746\ : InMux
    port map (
            O => \N__11255\,
            I => \N__11249\
        );

    \I__2745\ : Span4Mux_v
    port map (
            O => \N__11252\,
            I => \N__11246\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__11249\,
            I => \N__11243\
        );

    \I__2743\ : Span4Mux_h
    port map (
            O => \N__11246\,
            I => \N__11239\
        );

    \I__2742\ : Span4Mux_v
    port map (
            O => \N__11243\,
            I => \N__11236\
        );

    \I__2741\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11232\
        );

    \I__2740\ : Sp12to4
    port map (
            O => \N__11239\,
            I => \N__11226\
        );

    \I__2739\ : Sp12to4
    port map (
            O => \N__11236\,
            I => \N__11226\
        );

    \I__2738\ : InMux
    port map (
            O => \N__11235\,
            I => \N__11223\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__11232\,
            I => \N__11220\
        );

    \I__2736\ : InMux
    port map (
            O => \N__11231\,
            I => \N__11217\
        );

    \I__2735\ : Span12Mux_h
    port map (
            O => \N__11226\,
            I => \N__11210\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__11223\,
            I => \N__11207\
        );

    \I__2733\ : Span4Mux_h
    port map (
            O => \N__11220\,
            I => \N__11202\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__11217\,
            I => \N__11202\
        );

    \I__2731\ : InMux
    port map (
            O => \N__11216\,
            I => \N__11199\
        );

    \I__2730\ : InMux
    port map (
            O => \N__11215\,
            I => \N__11196\
        );

    \I__2729\ : InMux
    port map (
            O => \N__11214\,
            I => \N__11191\
        );

    \I__2728\ : InMux
    port map (
            O => \N__11213\,
            I => \N__11191\
        );

    \I__2727\ : Odrv12
    port map (
            O => \N__11210\,
            I => \WRITE_CYCLEm\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__11207\,
            I => \WRITE_CYCLEm\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__11202\,
            I => \WRITE_CYCLEm\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__11199\,
            I => \WRITE_CYCLEm\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__11196\,
            I => \WRITE_CYCLEm\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__11191\,
            I => \WRITE_CYCLEm\
        );

    \I__2721\ : InMux
    port map (
            O => \N__11178\,
            I => \N__11175\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__11175\,
            I => \N__11171\
        );

    \I__2719\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11166\
        );

    \I__2718\ : Span4Mux_h
    port map (
            O => \N__11171\,
            I => \N__11163\
        );

    \I__2717\ : InMux
    port map (
            O => \N__11170\,
            I => \N__11160\
        );

    \I__2716\ : InMux
    port map (
            O => \N__11169\,
            I => \N__11157\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__11166\,
            I => \N__11152\
        );

    \I__2714\ : Span4Mux_v
    port map (
            O => \N__11163\,
            I => \N__11149\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__11160\,
            I => \N__11144\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__11157\,
            I => \N__11144\
        );

    \I__2711\ : InMux
    port map (
            O => \N__11156\,
            I => \N__11139\
        );

    \I__2710\ : InMux
    port map (
            O => \N__11155\,
            I => \N__11139\
        );

    \I__2709\ : Span12Mux_v
    port map (
            O => \N__11152\,
            I => \N__11134\
        );

    \I__2708\ : Sp12to4
    port map (
            O => \N__11149\,
            I => \N__11134\
        );

    \I__2707\ : Span12Mux_h
    port map (
            O => \N__11144\,
            I => \N__11129\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__11139\,
            I => \N__11129\
        );

    \I__2705\ : Span12Mux_h
    port map (
            O => \N__11134\,
            I => \N__11124\
        );

    \I__2704\ : Span12Mux_v
    port map (
            O => \N__11129\,
            I => \N__11124\
        );

    \I__2703\ : Odrv12
    port map (
            O => \N__11124\,
            I => \CASLn_c\
        );

    \I__2702\ : IoInMux
    port map (
            O => \N__11121\,
            I => \N__11118\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__11118\,
            I => \N__11115\
        );

    \I__2700\ : Span12Mux_s4_h
    port map (
            O => \N__11115\,
            I => \N__11112\
        );

    \I__2699\ : Odrv12
    port map (
            O => \N__11112\,
            I => \N_450\
        );

    \I__2698\ : IoInMux
    port map (
            O => \N__11109\,
            I => \N__11106\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__11106\,
            I => \N__11103\
        );

    \I__2696\ : Span4Mux_s3_v
    port map (
            O => \N__11103\,
            I => \N__11100\
        );

    \I__2695\ : Span4Mux_h
    port map (
            O => \N__11100\,
            I => \N__11097\
        );

    \I__2694\ : Span4Mux_v
    port map (
            O => \N__11097\,
            I => \N__11094\
        );

    \I__2693\ : Odrv4
    port map (
            O => \N__11094\,
            I => \N_291\
        );

    \I__2692\ : IoInMux
    port map (
            O => \N__11091\,
            I => \N__11088\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__11088\,
            I => \N__11085\
        );

    \I__2690\ : IoSpan4Mux
    port map (
            O => \N__11085\,
            I => \N__11082\
        );

    \I__2689\ : Span4Mux_s2_v
    port map (
            O => \N__11082\,
            I => \N__11079\
        );

    \I__2688\ : Span4Mux_v
    port map (
            O => \N__11079\,
            I => \N__11076\
        );

    \I__2687\ : Odrv4
    port map (
            O => \N__11076\,
            I => \N_400_i\
        );

    \I__2686\ : InMux
    port map (
            O => \N__11073\,
            I => \N__11070\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__11070\,
            I => \N__11066\
        );

    \I__2684\ : InMux
    port map (
            O => \N__11069\,
            I => \N__11063\
        );

    \I__2683\ : Span4Mux_v
    port map (
            O => \N__11066\,
            I => \N__11058\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__11063\,
            I => \N__11058\
        );

    \I__2681\ : Span4Mux_v
    port map (
            O => \N__11058\,
            I => \N__11055\
        );

    \I__2680\ : Sp12to4
    port map (
            O => \N__11055\,
            I => \N__11051\
        );

    \I__2679\ : InMux
    port map (
            O => \N__11054\,
            I => \N__11048\
        );

    \I__2678\ : Odrv12
    port map (
            O => \N__11051\,
            I => \DS_ENm\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11048\,
            I => \DS_ENm\
        );

    \I__2676\ : IoInMux
    port map (
            O => \N__11043\,
            I => \N__11040\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__11040\,
            I => \N__11037\
        );

    \I__2674\ : Span4Mux_s2_v
    port map (
            O => \N__11037\,
            I => \N__11034\
        );

    \I__2673\ : Span4Mux_h
    port map (
            O => \N__11034\,
            I => \N__11031\
        );

    \I__2672\ : Span4Mux_v
    port map (
            O => \N__11031\,
            I => \N__11028\
        );

    \I__2671\ : Odrv4
    port map (
            O => \N__11028\,
            I => \N_293\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__11025\,
            I => \N__11020\
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__11024\,
            I => \N__11015\
        );

    \I__2668\ : InMux
    port map (
            O => \N__11023\,
            I => \N__11011\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11020\,
            I => \N__11004\
        );

    \I__2666\ : InMux
    port map (
            O => \N__11019\,
            I => \N__11004\
        );

    \I__2665\ : InMux
    port map (
            O => \N__11018\,
            I => \N__11004\
        );

    \I__2664\ : InMux
    port map (
            O => \N__11015\,
            I => \N__11001\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__11014\,
            I => \N__10998\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__11011\,
            I => \N__10995\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__11004\,
            I => \N__10990\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__11001\,
            I => \N__10990\
        );

    \I__2659\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10987\
        );

    \I__2658\ : Span4Mux_v
    port map (
            O => \N__10995\,
            I => \N__10979\
        );

    \I__2657\ : Span4Mux_h
    port map (
            O => \N__10990\,
            I => \N__10979\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__10987\,
            I => \N__10979\
        );

    \I__2655\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10976\
        );

    \I__2654\ : Span4Mux_h
    port map (
            O => \N__10979\,
            I => \N__10973\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__10976\,
            I => \N__10970\
        );

    \I__2652\ : Span4Mux_v
    port map (
            O => \N__10973\,
            I => \N__10967\
        );

    \I__2651\ : Span12Mux_v
    port map (
            O => \N__10970\,
            I => \N__10964\
        );

    \I__2650\ : Span4Mux_h
    port map (
            O => \N__10967\,
            I => \N__10961\
        );

    \I__2649\ : Span12Mux_h
    port map (
            O => \N__10964\,
            I => \N__10958\
        );

    \I__2648\ : Sp12to4
    port map (
            O => \N__10961\,
            I => \N__10955\
        );

    \I__2647\ : Odrv12
    port map (
            O => \N__10958\,
            I => \SIZ_c_0\
        );

    \I__2646\ : Odrv12
    port map (
            O => \N__10955\,
            I => \SIZ_c_0\
        );

    \I__2645\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10940\
        );

    \I__2644\ : InMux
    port map (
            O => \N__10949\,
            I => \N__10940\
        );

    \I__2643\ : InMux
    port map (
            O => \N__10948\,
            I => \N__10940\
        );

    \I__2642\ : InMux
    port map (
            O => \N__10947\,
            I => \N__10937\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__10940\,
            I => \N__10928\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__10937\,
            I => \N__10928\
        );

    \I__2639\ : InMux
    port map (
            O => \N__10936\,
            I => \N__10925\
        );

    \I__2638\ : InMux
    port map (
            O => \N__10935\,
            I => \N__10922\
        );

    \I__2637\ : InMux
    port map (
            O => \N__10934\,
            I => \N__10917\
        );

    \I__2636\ : InMux
    port map (
            O => \N__10933\,
            I => \N__10917\
        );

    \I__2635\ : Span4Mux_v
    port map (
            O => \N__10928\,
            I => \N__10914\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__10925\,
            I => \N__10909\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__10922\,
            I => \N__10909\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__10917\,
            I => \N__10906\
        );

    \I__2631\ : Span4Mux_v
    port map (
            O => \N__10914\,
            I => \N__10901\
        );

    \I__2630\ : Span4Mux_v
    port map (
            O => \N__10909\,
            I => \N__10901\
        );

    \I__2629\ : Span12Mux_s7_v
    port map (
            O => \N__10906\,
            I => \N__10898\
        );

    \I__2628\ : Sp12to4
    port map (
            O => \N__10901\,
            I => \N__10895\
        );

    \I__2627\ : Span12Mux_h
    port map (
            O => \N__10898\,
            I => \N__10892\
        );

    \I__2626\ : Span12Mux_h
    port map (
            O => \N__10895\,
            I => \N__10889\
        );

    \I__2625\ : Odrv12
    port map (
            O => \N__10892\,
            I => \A_c_1\
        );

    \I__2624\ : Odrv12
    port map (
            O => \N__10889\,
            I => \A_c_1\
        );

    \I__2623\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10878\
        );

    \I__2622\ : InMux
    port map (
            O => \N__10883\,
            I => \N__10875\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__10882\,
            I => \N__10870\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__10881\,
            I => \N__10866\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__10878\,
            I => \N__10859\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__10875\,
            I => \N__10859\
        );

    \I__2617\ : InMux
    port map (
            O => \N__10874\,
            I => \N__10854\
        );

    \I__2616\ : InMux
    port map (
            O => \N__10873\,
            I => \N__10854\
        );

    \I__2615\ : InMux
    port map (
            O => \N__10870\,
            I => \N__10851\
        );

    \I__2614\ : InMux
    port map (
            O => \N__10869\,
            I => \N__10844\
        );

    \I__2613\ : InMux
    port map (
            O => \N__10866\,
            I => \N__10844\
        );

    \I__2612\ : InMux
    port map (
            O => \N__10865\,
            I => \N__10844\
        );

    \I__2611\ : InMux
    port map (
            O => \N__10864\,
            I => \N__10841\
        );

    \I__2610\ : Span4Mux_v
    port map (
            O => \N__10859\,
            I => \N__10834\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__10854\,
            I => \N__10834\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__10851\,
            I => \N__10834\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__10844\,
            I => \N__10829\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__10841\,
            I => \N__10829\
        );

    \I__2605\ : Span4Mux_v
    port map (
            O => \N__10834\,
            I => \N__10826\
        );

    \I__2604\ : Span12Mux_s10_v
    port map (
            O => \N__10829\,
            I => \N__10821\
        );

    \I__2603\ : Sp12to4
    port map (
            O => \N__10826\,
            I => \N__10821\
        );

    \I__2602\ : Span12Mux_h
    port map (
            O => \N__10821\,
            I => \N__10818\
        );

    \I__2601\ : Odrv12
    port map (
            O => \N__10818\,
            I => \A_c_0\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__10815\,
            I => \N__10812\
        );

    \I__2599\ : InMux
    port map (
            O => \N__10812\,
            I => \N__10808\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__10811\,
            I => \N__10803\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__10808\,
            I => \N__10799\
        );

    \I__2596\ : InMux
    port map (
            O => \N__10807\,
            I => \N__10792\
        );

    \I__2595\ : InMux
    port map (
            O => \N__10806\,
            I => \N__10792\
        );

    \I__2594\ : InMux
    port map (
            O => \N__10803\,
            I => \N__10792\
        );

    \I__2593\ : InMux
    port map (
            O => \N__10802\,
            I => \N__10789\
        );

    \I__2592\ : Span4Mux_v
    port map (
            O => \N__10799\,
            I => \N__10782\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__10792\,
            I => \N__10782\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__10789\,
            I => \N__10782\
        );

    \I__2589\ : Span4Mux_h
    port map (
            O => \N__10782\,
            I => \N__10776\
        );

    \I__2588\ : InMux
    port map (
            O => \N__10781\,
            I => \N__10773\
        );

    \I__2587\ : InMux
    port map (
            O => \N__10780\,
            I => \N__10770\
        );

    \I__2586\ : InMux
    port map (
            O => \N__10779\,
            I => \N__10767\
        );

    \I__2585\ : Span4Mux_v
    port map (
            O => \N__10776\,
            I => \N__10764\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__10773\,
            I => \N__10757\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__10770\,
            I => \N__10757\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__10767\,
            I => \N__10757\
        );

    \I__2581\ : Sp12to4
    port map (
            O => \N__10764\,
            I => \N__10752\
        );

    \I__2580\ : Span12Mux_v
    port map (
            O => \N__10757\,
            I => \N__10752\
        );

    \I__2579\ : Span12Mux_h
    port map (
            O => \N__10752\,
            I => \N__10749\
        );

    \I__2578\ : Odrv12
    port map (
            O => \N__10749\,
            I => \SIZ_c_1\
        );

    \I__2577\ : IoInMux
    port map (
            O => \N__10746\,
            I => \N__10743\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__10743\,
            I => \N__10740\
        );

    \I__2575\ : Odrv12
    port map (
            O => \N__10740\,
            I => \N_401_i\
        );

    \I__2574\ : InMux
    port map (
            O => \N__10737\,
            I => \N__10733\
        );

    \I__2573\ : InMux
    port map (
            O => \N__10736\,
            I => \N__10730\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__10733\,
            I => \N__10725\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__10730\,
            I => \N__10722\
        );

    \I__2570\ : InMux
    port map (
            O => \N__10729\,
            I => \N__10719\
        );

    \I__2569\ : InMux
    port map (
            O => \N__10728\,
            I => \N__10716\
        );

    \I__2568\ : Span4Mux_v
    port map (
            O => \N__10725\,
            I => \N__10713\
        );

    \I__2567\ : Span4Mux_v
    port map (
            O => \N__10722\,
            I => \N__10710\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__10719\,
            I => \N__10707\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__10716\,
            I => \N__10702\
        );

    \I__2564\ : Sp12to4
    port map (
            O => \N__10713\,
            I => \N__10702\
        );

    \I__2563\ : Span4Mux_h
    port map (
            O => \N__10710\,
            I => \N__10697\
        );

    \I__2562\ : Span4Mux_v
    port map (
            O => \N__10707\,
            I => \N__10697\
        );

    \I__2561\ : Span12Mux_h
    port map (
            O => \N__10702\,
            I => \N__10694\
        );

    \I__2560\ : Sp12to4
    port map (
            O => \N__10697\,
            I => \N__10691\
        );

    \I__2559\ : Odrv12
    port map (
            O => \N__10694\,
            I => \DRA_c_8\
        );

    \I__2558\ : Odrv12
    port map (
            O => \N__10691\,
            I => \DRA_c_8\
        );

    \I__2557\ : InMux
    port map (
            O => \N__10686\,
            I => \N__10681\
        );

    \I__2556\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10677\
        );

    \I__2555\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10674\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__10681\,
            I => \N__10671\
        );

    \I__2553\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10668\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10677\,
            I => \N__10663\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__10674\,
            I => \N__10663\
        );

    \I__2550\ : Span4Mux_v
    port map (
            O => \N__10671\,
            I => \N__10660\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__10668\,
            I => \N__10657\
        );

    \I__2548\ : Span4Mux_v
    port map (
            O => \N__10663\,
            I => \N__10654\
        );

    \I__2547\ : Sp12to4
    port map (
            O => \N__10660\,
            I => \N__10647\
        );

    \I__2546\ : Span12Mux_v
    port map (
            O => \N__10657\,
            I => \N__10647\
        );

    \I__2545\ : Sp12to4
    port map (
            O => \N__10654\,
            I => \N__10647\
        );

    \I__2544\ : Span12Mux_h
    port map (
            O => \N__10647\,
            I => \N__10644\
        );

    \I__2543\ : Odrv12
    port map (
            O => \N__10644\,
            I => \DRA_c_7\
        );

    \I__2542\ : InMux
    port map (
            O => \N__10641\,
            I => \N__10638\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__10638\,
            I => \N__10635\
        );

    \I__2540\ : Span4Mux_h
    port map (
            O => \N__10635\,
            I => \N__10632\
        );

    \I__2539\ : Odrv4
    port map (
            O => \N__10632\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2538\ : InMux
    port map (
            O => \N__10629\,
            I => \N__10625\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__10628\,
            I => \N__10620\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10625\,
            I => \N__10616\
        );

    \I__2535\ : InMux
    port map (
            O => \N__10624\,
            I => \N__10613\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__10623\,
            I => \N__10604\
        );

    \I__2533\ : InMux
    port map (
            O => \N__10620\,
            I => \N__10593\
        );

    \I__2532\ : InMux
    port map (
            O => \N__10619\,
            I => \N__10593\
        );

    \I__2531\ : Span4Mux_v
    port map (
            O => \N__10616\,
            I => \N__10590\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__10613\,
            I => \N__10587\
        );

    \I__2529\ : InMux
    port map (
            O => \N__10612\,
            I => \N__10584\
        );

    \I__2528\ : InMux
    port map (
            O => \N__10611\,
            I => \N__10581\
        );

    \I__2527\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10578\
        );

    \I__2526\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10573\
        );

    \I__2525\ : InMux
    port map (
            O => \N__10608\,
            I => \N__10573\
        );

    \I__2524\ : InMux
    port map (
            O => \N__10607\,
            I => \N__10569\
        );

    \I__2523\ : InMux
    port map (
            O => \N__10604\,
            I => \N__10564\
        );

    \I__2522\ : InMux
    port map (
            O => \N__10603\,
            I => \N__10564\
        );

    \I__2521\ : InMux
    port map (
            O => \N__10602\,
            I => \N__10561\
        );

    \I__2520\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10556\
        );

    \I__2519\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10556\
        );

    \I__2518\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10551\
        );

    \I__2517\ : InMux
    port map (
            O => \N__10598\,
            I => \N__10551\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__10593\,
            I => \N__10546\
        );

    \I__2515\ : Span4Mux_h
    port map (
            O => \N__10590\,
            I => \N__10540\
        );

    \I__2514\ : Span4Mux_v
    port map (
            O => \N__10587\,
            I => \N__10540\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__10584\,
            I => \N__10537\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__10581\,
            I => \N__10532\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__10578\,
            I => \N__10532\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__10573\,
            I => \N__10529\
        );

    \I__2509\ : InMux
    port map (
            O => \N__10572\,
            I => \N__10526\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10569\,
            I => \N__10523\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__10564\,
            I => \N__10518\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__10561\,
            I => \N__10518\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__10556\,
            I => \N__10513\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__10551\,
            I => \N__10513\
        );

    \I__2503\ : InMux
    port map (
            O => \N__10550\,
            I => \N__10510\
        );

    \I__2502\ : InMux
    port map (
            O => \N__10549\,
            I => \N__10507\
        );

    \I__2501\ : Span4Mux_v
    port map (
            O => \N__10546\,
            I => \N__10504\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10501\
        );

    \I__2499\ : Span4Mux_h
    port map (
            O => \N__10540\,
            I => \N__10488\
        );

    \I__2498\ : Span4Mux_v
    port map (
            O => \N__10537\,
            I => \N__10488\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__10532\,
            I => \N__10488\
        );

    \I__2496\ : Span4Mux_h
    port map (
            O => \N__10529\,
            I => \N__10488\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__10526\,
            I => \N__10488\
        );

    \I__2494\ : Span4Mux_v
    port map (
            O => \N__10523\,
            I => \N__10488\
        );

    \I__2493\ : Sp12to4
    port map (
            O => \N__10518\,
            I => \N__10483\
        );

    \I__2492\ : Sp12to4
    port map (
            O => \N__10513\,
            I => \N__10483\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__10510\,
            I => \N__10478\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10507\,
            I => \N__10478\
        );

    \I__2489\ : Sp12to4
    port map (
            O => \N__10504\,
            I => \N__10471\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__10501\,
            I => \N__10471\
        );

    \I__2487\ : Sp12to4
    port map (
            O => \N__10488\,
            I => \N__10471\
        );

    \I__2486\ : Span12Mux_v
    port map (
            O => \N__10483\,
            I => \N__10468\
        );

    \I__2485\ : Span12Mux_h
    port map (
            O => \N__10478\,
            I => \N__10465\
        );

    \I__2484\ : Span12Mux_h
    port map (
            O => \N__10471\,
            I => \N__10462\
        );

    \I__2483\ : Span12Mux_h
    port map (
            O => \N__10468\,
            I => \N__10457\
        );

    \I__2482\ : Span12Mux_v
    port map (
            O => \N__10465\,
            I => \N__10457\
        );

    \I__2481\ : Span12Mux_v
    port map (
            O => \N__10462\,
            I => \N__10454\
        );

    \I__2480\ : Odrv12
    port map (
            O => \N__10457\,
            I => \AGNUS_REV_c\
        );

    \I__2479\ : Odrv12
    port map (
            O => \N__10454\,
            I => \AGNUS_REV_c\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10449\,
            I => \N__10446\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__10446\,
            I => \N__10443\
        );

    \I__2476\ : Span4Mux_v
    port map (
            O => \N__10443\,
            I => \N__10440\
        );

    \I__2475\ : Sp12to4
    port map (
            O => \N__10440\,
            I => \N__10437\
        );

    \I__2474\ : Odrv12
    port map (
            O => \N__10437\,
            I => \RAS0n_c\
        );

    \I__2473\ : InMux
    port map (
            O => \N__10434\,
            I => \N__10430\
        );

    \I__2472\ : InMux
    port map (
            O => \N__10433\,
            I => \N__10426\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__10430\,
            I => \N__10423\
        );

    \I__2470\ : InMux
    port map (
            O => \N__10429\,
            I => \N__10420\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__10426\,
            I => \N__10417\
        );

    \I__2468\ : Span4Mux_v
    port map (
            O => \N__10423\,
            I => \N__10411\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__10420\,
            I => \N__10411\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__10417\,
            I => \N__10408\
        );

    \I__2465\ : InMux
    port map (
            O => \N__10416\,
            I => \N__10405\
        );

    \I__2464\ : Span4Mux_v
    port map (
            O => \N__10411\,
            I => \N__10402\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__10408\,
            I => \N__10399\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__10405\,
            I => \N__10396\
        );

    \I__2461\ : Sp12to4
    port map (
            O => \N__10402\,
            I => \N__10391\
        );

    \I__2460\ : Sp12to4
    port map (
            O => \N__10399\,
            I => \N__10391\
        );

    \I__2459\ : Span12Mux_h
    port map (
            O => \N__10396\,
            I => \N__10388\
        );

    \I__2458\ : Span12Mux_h
    port map (
            O => \N__10391\,
            I => \N__10385\
        );

    \I__2457\ : Span12Mux_v
    port map (
            O => \N__10388\,
            I => \N__10382\
        );

    \I__2456\ : Span12Mux_v
    port map (
            O => \N__10385\,
            I => \N__10379\
        );

    \I__2455\ : Odrv12
    port map (
            O => \N__10382\,
            I => \DRA_c_9\
        );

    \I__2454\ : Odrv12
    port map (
            O => \N__10379\,
            I => \DRA_c_9\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10374\,
            I => \N__10371\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__10371\,
            I => \N__10368\
        );

    \I__2451\ : Odrv12
    port map (
            O => \N__10368\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2450\ : ClkMux
    port map (
            O => \N__10365\,
            I => \N__10344\
        );

    \I__2449\ : ClkMux
    port map (
            O => \N__10364\,
            I => \N__10344\
        );

    \I__2448\ : ClkMux
    port map (
            O => \N__10363\,
            I => \N__10344\
        );

    \I__2447\ : ClkMux
    port map (
            O => \N__10362\,
            I => \N__10344\
        );

    \I__2446\ : ClkMux
    port map (
            O => \N__10361\,
            I => \N__10344\
        );

    \I__2445\ : ClkMux
    port map (
            O => \N__10360\,
            I => \N__10344\
        );

    \I__2444\ : ClkMux
    port map (
            O => \N__10359\,
            I => \N__10344\
        );

    \I__2443\ : GlobalMux
    port map (
            O => \N__10344\,
            I => \N__10341\
        );

    \I__2442\ : gio2CtrlBuf
    port map (
            O => \N__10341\,
            I => \C3_c_g\
        );

    \I__2441\ : CEMux
    port map (
            O => \N__10338\,
            I => \N__10299\
        );

    \I__2440\ : CEMux
    port map (
            O => \N__10337\,
            I => \N__10299\
        );

    \I__2439\ : CEMux
    port map (
            O => \N__10336\,
            I => \N__10299\
        );

    \I__2438\ : CEMux
    port map (
            O => \N__10335\,
            I => \N__10299\
        );

    \I__2437\ : CEMux
    port map (
            O => \N__10334\,
            I => \N__10299\
        );

    \I__2436\ : CEMux
    port map (
            O => \N__10333\,
            I => \N__10299\
        );

    \I__2435\ : CEMux
    port map (
            O => \N__10332\,
            I => \N__10299\
        );

    \I__2434\ : CEMux
    port map (
            O => \N__10331\,
            I => \N__10299\
        );

    \I__2433\ : CEMux
    port map (
            O => \N__10330\,
            I => \N__10299\
        );

    \I__2432\ : CEMux
    port map (
            O => \N__10329\,
            I => \N__10299\
        );

    \I__2431\ : CEMux
    port map (
            O => \N__10328\,
            I => \N__10299\
        );

    \I__2430\ : CEMux
    port map (
            O => \N__10327\,
            I => \N__10299\
        );

    \I__2429\ : CEMux
    port map (
            O => \N__10326\,
            I => \N__10299\
        );

    \I__2428\ : GlobalMux
    port map (
            O => \N__10299\,
            I => \N__10296\
        );

    \I__2427\ : gio2CtrlBuf
    port map (
            O => \N__10296\,
            I => \DBRn_c_i_0_g\
        );

    \I__2426\ : InMux
    port map (
            O => \N__10293\,
            I => \N__10286\
        );

    \I__2425\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10283\
        );

    \I__2424\ : InMux
    port map (
            O => \N__10291\,
            I => \N__10280\
        );

    \I__2423\ : InMux
    port map (
            O => \N__10290\,
            I => \N__10277\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10289\,
            I => \N__10274\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__10286\,
            I => \N__10265\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__10283\,
            I => \N__10262\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__10280\,
            I => \N__10250\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__10277\,
            I => \N__10240\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__10274\,
            I => \N__10233\
        );

    \I__2416\ : SRMux
    port map (
            O => \N__10273\,
            I => \N__10146\
        );

    \I__2415\ : SRMux
    port map (
            O => \N__10272\,
            I => \N__10146\
        );

    \I__2414\ : SRMux
    port map (
            O => \N__10271\,
            I => \N__10146\
        );

    \I__2413\ : SRMux
    port map (
            O => \N__10270\,
            I => \N__10146\
        );

    \I__2412\ : SRMux
    port map (
            O => \N__10269\,
            I => \N__10146\
        );

    \I__2411\ : SRMux
    port map (
            O => \N__10268\,
            I => \N__10146\
        );

    \I__2410\ : Glb2LocalMux
    port map (
            O => \N__10265\,
            I => \N__10146\
        );

    \I__2409\ : Glb2LocalMux
    port map (
            O => \N__10262\,
            I => \N__10146\
        );

    \I__2408\ : SRMux
    port map (
            O => \N__10261\,
            I => \N__10146\
        );

    \I__2407\ : SRMux
    port map (
            O => \N__10260\,
            I => \N__10146\
        );

    \I__2406\ : SRMux
    port map (
            O => \N__10259\,
            I => \N__10146\
        );

    \I__2405\ : SRMux
    port map (
            O => \N__10258\,
            I => \N__10146\
        );

    \I__2404\ : SRMux
    port map (
            O => \N__10257\,
            I => \N__10146\
        );

    \I__2403\ : SRMux
    port map (
            O => \N__10256\,
            I => \N__10146\
        );

    \I__2402\ : SRMux
    port map (
            O => \N__10255\,
            I => \N__10146\
        );

    \I__2401\ : SRMux
    port map (
            O => \N__10254\,
            I => \N__10146\
        );

    \I__2400\ : SRMux
    port map (
            O => \N__10253\,
            I => \N__10146\
        );

    \I__2399\ : Glb2LocalMux
    port map (
            O => \N__10250\,
            I => \N__10146\
        );

    \I__2398\ : SRMux
    port map (
            O => \N__10249\,
            I => \N__10146\
        );

    \I__2397\ : SRMux
    port map (
            O => \N__10248\,
            I => \N__10146\
        );

    \I__2396\ : SRMux
    port map (
            O => \N__10247\,
            I => \N__10146\
        );

    \I__2395\ : SRMux
    port map (
            O => \N__10246\,
            I => \N__10146\
        );

    \I__2394\ : SRMux
    port map (
            O => \N__10245\,
            I => \N__10146\
        );

    \I__2393\ : SRMux
    port map (
            O => \N__10244\,
            I => \N__10146\
        );

    \I__2392\ : SRMux
    port map (
            O => \N__10243\,
            I => \N__10146\
        );

    \I__2391\ : Glb2LocalMux
    port map (
            O => \N__10240\,
            I => \N__10146\
        );

    \I__2390\ : SRMux
    port map (
            O => \N__10239\,
            I => \N__10146\
        );

    \I__2389\ : SRMux
    port map (
            O => \N__10238\,
            I => \N__10146\
        );

    \I__2388\ : SRMux
    port map (
            O => \N__10237\,
            I => \N__10146\
        );

    \I__2387\ : SRMux
    port map (
            O => \N__10236\,
            I => \N__10146\
        );

    \I__2386\ : Glb2LocalMux
    port map (
            O => \N__10233\,
            I => \N__10146\
        );

    \I__2385\ : SRMux
    port map (
            O => \N__10232\,
            I => \N__10146\
        );

    \I__2384\ : SRMux
    port map (
            O => \N__10231\,
            I => \N__10146\
        );

    \I__2383\ : SRMux
    port map (
            O => \N__10230\,
            I => \N__10146\
        );

    \I__2382\ : SRMux
    port map (
            O => \N__10229\,
            I => \N__10146\
        );

    \I__2381\ : SRMux
    port map (
            O => \N__10228\,
            I => \N__10146\
        );

    \I__2380\ : SRMux
    port map (
            O => \N__10227\,
            I => \N__10146\
        );

    \I__2379\ : SRMux
    port map (
            O => \N__10226\,
            I => \N__10146\
        );

    \I__2378\ : SRMux
    port map (
            O => \N__10225\,
            I => \N__10146\
        );

    \I__2377\ : GlobalMux
    port map (
            O => \N__10146\,
            I => \N__10143\
        );

    \I__2376\ : gio2CtrlBuf
    port map (
            O => \N__10143\,
            I => \RESETn_c_i_g\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10140\,
            I => \N__10137\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__10137\,
            I => \N__10134\
        );

    \I__2373\ : Span4Mux_v
    port map (
            O => \N__10134\,
            I => \N__10131\
        );

    \I__2372\ : Span4Mux_h
    port map (
            O => \N__10131\,
            I => \N__10127\
        );

    \I__2371\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10124\
        );

    \I__2370\ : Sp12to4
    port map (
            O => \N__10127\,
            I => \N__10121\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__10124\,
            I => \N__10118\
        );

    \I__2368\ : Span12Mux_h
    port map (
            O => \N__10121\,
            I => \N__10114\
        );

    \I__2367\ : Span4Mux_v
    port map (
            O => \N__10118\,
            I => \N__10111\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10117\,
            I => \N__10108\
        );

    \I__2365\ : Odrv12
    port map (
            O => \N__10114\,
            I => \REG_CYCLEm\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__10111\,
            I => \REG_CYCLEm\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__10108\,
            I => \REG_CYCLEm\
        );

    \I__2362\ : IoInMux
    port map (
            O => \N__10101\,
            I => \N__10098\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__10098\,
            I => \N__10095\
        );

    \I__2360\ : Span4Mux_s2_v
    port map (
            O => \N__10095\,
            I => \N__10092\
        );

    \I__2359\ : Span4Mux_v
    port map (
            O => \N__10092\,
            I => \N__10089\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__10089\,
            I => \DRDENn_c\
        );

    \I__2357\ : InMux
    port map (
            O => \N__10086\,
            I => \N__10083\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10083\,
            I => \N__10079\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10076\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__10079\,
            I => \N__10073\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__10076\,
            I => \N__10069\
        );

    \I__2352\ : Span4Mux_v
    port map (
            O => \N__10073\,
            I => \N__10065\
        );

    \I__2351\ : InMux
    port map (
            O => \N__10072\,
            I => \N__10062\
        );

    \I__2350\ : Span4Mux_v
    port map (
            O => \N__10069\,
            I => \N__10059\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10068\,
            I => \N__10056\
        );

    \I__2348\ : Sp12to4
    port map (
            O => \N__10065\,
            I => \N__10053\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__10062\,
            I => \N__10050\
        );

    \I__2346\ : Sp12to4
    port map (
            O => \N__10059\,
            I => \N__10045\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10056\,
            I => \N__10045\
        );

    \I__2344\ : Span12Mux_h
    port map (
            O => \N__10053\,
            I => \N__10040\
        );

    \I__2343\ : Span12Mux_v
    port map (
            O => \N__10050\,
            I => \N__10040\
        );

    \I__2342\ : Span12Mux_h
    port map (
            O => \N__10045\,
            I => \N__10037\
        );

    \I__2341\ : Span12Mux_h
    port map (
            O => \N__10040\,
            I => \N__10032\
        );

    \I__2340\ : Span12Mux_v
    port map (
            O => \N__10037\,
            I => \N__10032\
        );

    \I__2339\ : Odrv12
    port map (
            O => \N__10032\,
            I => \RnW_c\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10029\,
            I => \N__10025\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__10028\,
            I => \N__10021\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__10025\,
            I => \N__10016\
        );

    \I__2335\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10011\
        );

    \I__2334\ : InMux
    port map (
            O => \N__10021\,
            I => \N__10011\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10008\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__10019\,
            I => \N__10005\
        );

    \I__2331\ : Sp12to4
    port map (
            O => \N__10016\,
            I => \N__9997\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__10011\,
            I => \N__9997\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10008\,
            I => \N__9997\
        );

    \I__2328\ : InMux
    port map (
            O => \N__10005\,
            I => \N__9992\
        );

    \I__2327\ : InMux
    port map (
            O => \N__10004\,
            I => \N__9992\
        );

    \I__2326\ : Span12Mux_v
    port map (
            O => \N__9997\,
            I => \N__9989\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__9992\,
            I => \N__9986\
        );

    \I__2324\ : Span12Mux_h
    port map (
            O => \N__9989\,
            I => \N__9983\
        );

    \I__2323\ : Span4Mux_v
    port map (
            O => \N__9986\,
            I => \N__9980\
        );

    \I__2322\ : Odrv12
    port map (
            O => \N__9983\,
            I => \CASUn_c\
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__9980\,
            I => \CASUn_c\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__9975\,
            I => \N__9971\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__9974\,
            I => \N__9968\
        );

    \I__2318\ : InMux
    port map (
            O => \N__9971\,
            I => \N__9954\
        );

    \I__2317\ : InMux
    port map (
            O => \N__9968\,
            I => \N__9954\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__9967\,
            I => \N__9947\
        );

    \I__2315\ : InMux
    port map (
            O => \N__9966\,
            I => \N__9942\
        );

    \I__2314\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9939\
        );

    \I__2313\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9933\
        );

    \I__2312\ : InMux
    port map (
            O => \N__9963\,
            I => \N__9925\
        );

    \I__2311\ : InMux
    port map (
            O => \N__9962\,
            I => \N__9925\
        );

    \I__2310\ : InMux
    port map (
            O => \N__9961\,
            I => \N__9925\
        );

    \I__2309\ : InMux
    port map (
            O => \N__9960\,
            I => \N__9922\
        );

    \I__2308\ : CascadeMux
    port map (
            O => \N__9959\,
            I => \N__9919\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__9954\,
            I => \N__9915\
        );

    \I__2306\ : InMux
    port map (
            O => \N__9953\,
            I => \N__9908\
        );

    \I__2305\ : InMux
    port map (
            O => \N__9952\,
            I => \N__9908\
        );

    \I__2304\ : InMux
    port map (
            O => \N__9951\,
            I => \N__9908\
        );

    \I__2303\ : InMux
    port map (
            O => \N__9950\,
            I => \N__9905\
        );

    \I__2302\ : InMux
    port map (
            O => \N__9947\,
            I => \N__9902\
        );

    \I__2301\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9899\
        );

    \I__2300\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9896\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__9942\,
            I => \N__9892\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__9939\,
            I => \N__9889\
        );

    \I__2297\ : InMux
    port map (
            O => \N__9938\,
            I => \N__9886\
        );

    \I__2296\ : InMux
    port map (
            O => \N__9937\,
            I => \N__9881\
        );

    \I__2295\ : InMux
    port map (
            O => \N__9936\,
            I => \N__9881\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__9933\,
            I => \N__9878\
        );

    \I__2293\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9875\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__9925\,
            I => \N__9872\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__9922\,
            I => \N__9869\
        );

    \I__2290\ : InMux
    port map (
            O => \N__9919\,
            I => \N__9866\
        );

    \I__2289\ : InMux
    port map (
            O => \N__9918\,
            I => \N__9863\
        );

    \I__2288\ : Span4Mux_v
    port map (
            O => \N__9915\,
            I => \N__9854\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__9908\,
            I => \N__9854\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__9905\,
            I => \N__9854\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__9902\,
            I => \N__9854\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__9899\,
            I => \N__9849\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__9896\,
            I => \N__9849\
        );

    \I__2282\ : InMux
    port map (
            O => \N__9895\,
            I => \N__9846\
        );

    \I__2281\ : Span4Mux_h
    port map (
            O => \N__9892\,
            I => \N__9839\
        );

    \I__2280\ : Span4Mux_v
    port map (
            O => \N__9889\,
            I => \N__9839\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__9886\,
            I => \N__9839\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__9881\,
            I => \N__9836\
        );

    \I__2277\ : Span4Mux_h
    port map (
            O => \N__9878\,
            I => \N__9831\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__9875\,
            I => \N__9831\
        );

    \I__2275\ : Span4Mux_v
    port map (
            O => \N__9872\,
            I => \N__9822\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__9869\,
            I => \N__9822\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__9866\,
            I => \N__9822\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__9863\,
            I => \N__9822\
        );

    \I__2271\ : Span4Mux_h
    port map (
            O => \N__9854\,
            I => \N__9819\
        );

    \I__2270\ : Span12Mux_h
    port map (
            O => \N__9849\,
            I => \N__9814\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__9846\,
            I => \N__9814\
        );

    \I__2268\ : Span4Mux_v
    port map (
            O => \N__9839\,
            I => \N__9805\
        );

    \I__2267\ : Span4Mux_h
    port map (
            O => \N__9836\,
            I => \N__9805\
        );

    \I__2266\ : Span4Mux_v
    port map (
            O => \N__9831\,
            I => \N__9805\
        );

    \I__2265\ : Span4Mux_h
    port map (
            O => \N__9822\,
            I => \N__9805\
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__9819\,
            I => \CPU_CYCLEm\
        );

    \I__2263\ : Odrv12
    port map (
            O => \N__9814\,
            I => \CPU_CYCLEm\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__9805\,
            I => \CPU_CYCLEm\
        );

    \I__2261\ : InMux
    port map (
            O => \N__9798\,
            I => \N__9795\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__9795\,
            I => \N__9792\
        );

    \I__2259\ : Odrv12
    port map (
            O => \N__9792\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__9789\,
            I => \N__9783\
        );

    \I__2257\ : InMux
    port map (
            O => \N__9788\,
            I => \N__9776\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__9787\,
            I => \N__9773\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__9786\,
            I => \N__9770\
        );

    \I__2254\ : InMux
    port map (
            O => \N__9783\,
            I => \N__9765\
        );

    \I__2253\ : InMux
    port map (
            O => \N__9782\,
            I => \N__9765\
        );

    \I__2252\ : InMux
    port map (
            O => \N__9781\,
            I => \N__9760\
        );

    \I__2251\ : InMux
    port map (
            O => \N__9780\,
            I => \N__9760\
        );

    \I__2250\ : CascadeMux
    port map (
            O => \N__9779\,
            I => \N__9755\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__9776\,
            I => \N__9752\
        );

    \I__2248\ : InMux
    port map (
            O => \N__9773\,
            I => \N__9749\
        );

    \I__2247\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9746\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__9765\,
            I => \N__9733\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__9760\,
            I => \N__9733\
        );

    \I__2244\ : InMux
    port map (
            O => \N__9759\,
            I => \N__9726\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9758\,
            I => \N__9726\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9726\
        );

    \I__2241\ : Span4Mux_v
    port map (
            O => \N__9752\,
            I => \N__9721\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__9749\,
            I => \N__9721\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__9746\,
            I => \N__9718\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9745\,
            I => \N__9714\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9744\,
            I => \N__9711\
        );

    \I__2236\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9706\
        );

    \I__2235\ : InMux
    port map (
            O => \N__9742\,
            I => \N__9706\
        );

    \I__2234\ : InMux
    port map (
            O => \N__9741\,
            I => \N__9699\
        );

    \I__2233\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9699\
        );

    \I__2232\ : InMux
    port map (
            O => \N__9739\,
            I => \N__9699\
        );

    \I__2231\ : InMux
    port map (
            O => \N__9738\,
            I => \N__9691\
        );

    \I__2230\ : Span4Mux_v
    port map (
            O => \N__9733\,
            I => \N__9688\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__9726\,
            I => \N__9683\
        );

    \I__2228\ : Span4Mux_h
    port map (
            O => \N__9721\,
            I => \N__9683\
        );

    \I__2227\ : Span12Mux_v
    port map (
            O => \N__9718\,
            I => \N__9680\
        );

    \I__2226\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9677\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__9714\,
            I => \N__9672\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__9711\,
            I => \N__9672\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__9706\,
            I => \N__9667\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__9699\,
            I => \N__9667\
        );

    \I__2221\ : InMux
    port map (
            O => \N__9698\,
            I => \N__9662\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9697\,
            I => \N__9662\
        );

    \I__2219\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9657\
        );

    \I__2218\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9657\
        );

    \I__2217\ : InMux
    port map (
            O => \N__9694\,
            I => \N__9654\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__9691\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_1\
        );

    \I__2215\ : Odrv4
    port map (
            O => \N__9688\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_1\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__9683\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_1\
        );

    \I__2213\ : Odrv12
    port map (
            O => \N__9680\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_1\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__9677\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_1\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__9672\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_1\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__9667\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_1\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__9662\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_1\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__9657\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_1\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__9654\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_1\
        );

    \I__2206\ : InMux
    port map (
            O => \N__9633\,
            I => \N__9630\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__9630\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__2204\ : InMux
    port map (
            O => \N__9627\,
            I => \N__9624\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__9624\,
            I => \N__9621\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__9621\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2201\ : InMux
    port map (
            O => \N__9618\,
            I => \N__9615\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__9615\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__9612\,
            I => \N__9609\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9609\,
            I => \N__9606\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__9606\,
            I => \N__9603\
        );

    \I__2196\ : Span4Mux_h
    port map (
            O => \N__9603\,
            I => \N__9600\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__9600\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9597\,
            I => \N__9594\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__9594\,
            I => \N__9591\
        );

    \I__2192\ : Odrv4
    port map (
            O => \N__9591\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9583\
        );

    \I__2190\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9579\
        );

    \I__2189\ : InMux
    port map (
            O => \N__9586\,
            I => \N__9576\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__9583\,
            I => \N__9573\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9582\,
            I => \N__9570\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9579\,
            I => \N__9565\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__9576\,
            I => \N__9565\
        );

    \I__2184\ : Span4Mux_v
    port map (
            O => \N__9573\,
            I => \N__9560\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__9570\,
            I => \N__9560\
        );

    \I__2182\ : Span4Mux_h
    port map (
            O => \N__9565\,
            I => \N__9557\
        );

    \I__2181\ : Span4Mux_h
    port map (
            O => \N__9560\,
            I => \N__9554\
        );

    \I__2180\ : Sp12to4
    port map (
            O => \N__9557\,
            I => \N__9549\
        );

    \I__2179\ : Sp12to4
    port map (
            O => \N__9554\,
            I => \N__9549\
        );

    \I__2178\ : Span12Mux_v
    port map (
            O => \N__9549\,
            I => \N__9546\
        );

    \I__2177\ : Odrv12
    port map (
            O => \N__9546\,
            I => \DRA_c_1\
        );

    \I__2176\ : InMux
    port map (
            O => \N__9543\,
            I => \N__9540\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__9540\,
            I => \N__9536\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9533\
        );

    \I__2173\ : Span4Mux_v
    port map (
            O => \N__9536\,
            I => \N__9528\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9533\,
            I => \N__9528\
        );

    \I__2171\ : Sp12to4
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__2170\ : Span12Mux_v
    port map (
            O => \N__9525\,
            I => \N__9522\
        );

    \I__2169\ : Span12Mux_h
    port map (
            O => \N__9522\,
            I => \N__9519\
        );

    \I__2168\ : Odrv12
    port map (
            O => \N__9519\,
            I => \DRA_c_0\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9516\,
            I => \N__9513\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__9513\,
            I => \N__9510\
        );

    \I__2165\ : Odrv12
    port map (
            O => \N__9510\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2164\ : IoInMux
    port map (
            O => \N__9507\,
            I => \N__9504\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__9504\,
            I => \N__9501\
        );

    \I__2162\ : Span4Mux_s3_v
    port map (
            O => \N__9501\,
            I => \N__9498\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__9498\,
            I => \N_402_i\
        );

    \I__2160\ : InMux
    port map (
            O => \N__9495\,
            I => \N__9490\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9487\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9493\,
            I => \N__9483\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9490\,
            I => \N__9478\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__9487\,
            I => \N__9478\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9475\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9483\,
            I => \N__9472\
        );

    \I__2153\ : Span4Mux_v
    port map (
            O => \N__9478\,
            I => \N__9467\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__9475\,
            I => \N__9467\
        );

    \I__2151\ : Span4Mux_v
    port map (
            O => \N__9472\,
            I => \N__9464\
        );

    \I__2150\ : Span4Mux_h
    port map (
            O => \N__9467\,
            I => \N__9461\
        );

    \I__2149\ : Span4Mux_v
    port map (
            O => \N__9464\,
            I => \N__9458\
        );

    \I__2148\ : Span4Mux_v
    port map (
            O => \N__9461\,
            I => \N__9455\
        );

    \I__2147\ : Sp12to4
    port map (
            O => \N__9458\,
            I => \N__9450\
        );

    \I__2146\ : Sp12to4
    port map (
            O => \N__9455\,
            I => \N__9450\
        );

    \I__2145\ : Odrv12
    port map (
            O => \N__9450\,
            I => \DRA_c_6\
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__9447\,
            I => \N__9444\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9444\,
            I => \N__9441\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9441\,
            I => \N__9438\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__9438\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9435\,
            I => \N__9432\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__9432\,
            I => \N__9426\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9423\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9430\,
            I => \N__9420\
        );

    \I__2136\ : InMux
    port map (
            O => \N__9429\,
            I => \N__9417\
        );

    \I__2135\ : Span4Mux_h
    port map (
            O => \N__9426\,
            I => \N__9410\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9423\,
            I => \N__9410\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__9420\,
            I => \N__9410\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9417\,
            I => \N__9407\
        );

    \I__2131\ : Span4Mux_h
    port map (
            O => \N__9410\,
            I => \N__9404\
        );

    \I__2130\ : Span4Mux_v
    port map (
            O => \N__9407\,
            I => \N__9401\
        );

    \I__2129\ : Sp12to4
    port map (
            O => \N__9404\,
            I => \N__9398\
        );

    \I__2128\ : Span4Mux_v
    port map (
            O => \N__9401\,
            I => \N__9395\
        );

    \I__2127\ : Span12Mux_v
    port map (
            O => \N__9398\,
            I => \N__9390\
        );

    \I__2126\ : Sp12to4
    port map (
            O => \N__9395\,
            I => \N__9390\
        );

    \I__2125\ : Odrv12
    port map (
            O => \N__9390\,
            I => \DRA_c_5\
        );

    \I__2124\ : InMux
    port map (
            O => \N__9387\,
            I => \N__9383\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9386\,
            I => \N__9379\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9383\,
            I => \N__9376\
        );

    \I__2121\ : InMux
    port map (
            O => \N__9382\,
            I => \N__9373\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9379\,
            I => \N__9370\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__9376\,
            I => \N__9364\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9373\,
            I => \N__9364\
        );

    \I__2117\ : Span4Mux_v
    port map (
            O => \N__9370\,
            I => \N__9361\
        );

    \I__2116\ : InMux
    port map (
            O => \N__9369\,
            I => \N__9358\
        );

    \I__2115\ : Span4Mux_h
    port map (
            O => \N__9364\,
            I => \N__9355\
        );

    \I__2114\ : Span4Mux_v
    port map (
            O => \N__9361\,
            I => \N__9352\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__9358\,
            I => \N__9349\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__9355\,
            I => \N__9346\
        );

    \I__2111\ : Sp12to4
    port map (
            O => \N__9352\,
            I => \N__9339\
        );

    \I__2110\ : Span12Mux_v
    port map (
            O => \N__9349\,
            I => \N__9339\
        );

    \I__2109\ : Sp12to4
    port map (
            O => \N__9346\,
            I => \N__9339\
        );

    \I__2108\ : Span12Mux_h
    port map (
            O => \N__9339\,
            I => \N__9336\
        );

    \I__2107\ : Odrv12
    port map (
            O => \N__9336\,
            I => \DRA_c_4\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9333\,
            I => \N__9330\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__9330\,
            I => \N__9327\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__9327\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__9324\,
            I => \N__9321\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9321\,
            I => \N__9318\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9318\,
            I => \U712_BYTE_ENABLE.N_377\
        );

    \I__2100\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9312\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9312\,
            I => \U712_BYTE_ENABLE.N_530\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9309\,
            I => \N__9306\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__9306\,
            I => \N__9303\
        );

    \I__2096\ : Odrv4
    port map (
            O => \N__9303\,
            I => \U712_BYTE_ENABLE.N_532\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__9300\,
            I => \N__9297\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9291\
        );

    \I__2093\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9286\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9286\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9294\,
            I => \N__9283\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9291\,
            I => \N__9278\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__9286\,
            I => \N__9278\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__9283\,
            I => \N__9275\
        );

    \I__2087\ : Odrv12
    port map (
            O => \N__9278\,
            I => \U712_BYTE_ENABLE.N_364_i\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__9275\,
            I => \U712_BYTE_ENABLE.N_364_i\
        );

    \I__2085\ : IoInMux
    port map (
            O => \N__9270\,
            I => \N__9267\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__9267\,
            I => \N__9264\
        );

    \I__2083\ : Span4Mux_s1_v
    port map (
            O => \N__9264\,
            I => \N__9261\
        );

    \I__2082\ : Sp12to4
    port map (
            O => \N__9261\,
            I => \N__9258\
        );

    \I__2081\ : Span12Mux_h
    port map (
            O => \N__9258\,
            I => \N__9255\
        );

    \I__2080\ : Odrv12
    port map (
            O => \N__9255\,
            I => \DMA_LATCH_EN_c\
        );

    \I__2079\ : IoInMux
    port map (
            O => \N__9252\,
            I => \N__9249\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__9249\,
            I => \N__9246\
        );

    \I__2077\ : Span4Mux_s3_v
    port map (
            O => \N__9246\,
            I => \N__9243\
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__9243\,
            I => \N_403_i\
        );

    \I__2075\ : IoInMux
    port map (
            O => \N__9240\,
            I => \N__9237\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__9237\,
            I => \N__9234\
        );

    \I__2073\ : Span4Mux_s1_v
    port map (
            O => \N__9234\,
            I => \N__9231\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__9231\,
            I => \N__9228\
        );

    \I__2071\ : Span4Mux_v
    port map (
            O => \N__9228\,
            I => \N__9225\
        );

    \I__2070\ : Sp12to4
    port map (
            O => \N__9225\,
            I => \N__9222\
        );

    \I__2069\ : Odrv12
    port map (
            O => \N__9222\,
            I => \CASn_c\
        );

    \I__2068\ : IoInMux
    port map (
            O => \N__9219\,
            I => \N__9216\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__9216\,
            I => \N__9213\
        );

    \I__2066\ : IoSpan4Mux
    port map (
            O => \N__9213\,
            I => \N__9210\
        );

    \I__2065\ : Span4Mux_s3_v
    port map (
            O => \N__9210\,
            I => \N__9207\
        );

    \I__2064\ : Span4Mux_v
    port map (
            O => \N__9207\,
            I => \N__9204\
        );

    \I__2063\ : Sp12to4
    port map (
            O => \N__9204\,
            I => \N__9201\
        );

    \I__2062\ : Span12Mux_h
    port map (
            O => \N__9201\,
            I => \N__9198\
        );

    \I__2061\ : Odrv12
    port map (
            O => \N__9198\,
            I => \CMA_c_4\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__9195\,
            I => \N__9188\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__9194\,
            I => \N__9185\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__9193\,
            I => \N__9182\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__9192\,
            I => \N__9179\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9191\,
            I => \N__9174\
        );

    \I__2055\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9174\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9170\
        );

    \I__2053\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9167\
        );

    \I__2052\ : InMux
    port map (
            O => \N__9179\,
            I => \N__9164\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__9174\,
            I => \N__9161\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__9173\,
            I => \N__9158\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9170\,
            I => \N__9155\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9167\,
            I => \N__9148\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9164\,
            I => \N__9148\
        );

    \I__2046\ : Span4Mux_h
    port map (
            O => \N__9161\,
            I => \N__9148\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9145\
        );

    \I__2044\ : Span4Mux_h
    port map (
            O => \N__9155\,
            I => \N__9142\
        );

    \I__2043\ : Span4Mux_v
    port map (
            O => \N__9148\,
            I => \N__9139\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9145\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__9142\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__9139\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9132\,
            I => \N__9128\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__9131\,
            I => \N__9122\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__9128\,
            I => \N__9118\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9127\,
            I => \N__9113\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9126\,
            I => \N__9113\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9125\,
            I => \N__9109\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9104\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9121\,
            I => \N__9104\
        );

    \I__2031\ : Span4Mux_v
    port map (
            O => \N__9118\,
            I => \N__9099\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9113\,
            I => \N__9099\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9112\,
            I => \N__9096\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9109\,
            I => \N__9085\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__9104\,
            I => \N__9085\
        );

    \I__2026\ : Span4Mux_v
    port map (
            O => \N__9099\,
            I => \N__9085\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__9096\,
            I => \N__9085\
        );

    \I__2024\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9082\
        );

    \I__2023\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9079\
        );

    \I__2022\ : Span4Mux_h
    port map (
            O => \N__9085\,
            I => \N__9076\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9082\,
            I => \U712_CHIP_RAM.N_379\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__9079\,
            I => \U712_CHIP_RAM.N_379\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__9076\,
            I => \U712_CHIP_RAM.N_379\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9069\,
            I => \N__9066\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__9066\,
            I => \N__9063\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__9063\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__2015\ : IoInMux
    port map (
            O => \N__9060\,
            I => \N__9057\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__9057\,
            I => \N__9054\
        );

    \I__2013\ : Span4Mux_s3_h
    port map (
            O => \N__9054\,
            I => \N__9051\
        );

    \I__2012\ : Sp12to4
    port map (
            O => \N__9051\,
            I => \N__9048\
        );

    \I__2011\ : Span12Mux_s11_v
    port map (
            O => \N__9048\,
            I => \N__9045\
        );

    \I__2010\ : Odrv12
    port map (
            O => \N__9045\,
            I => \CMA_c_6\
        );

    \I__2009\ : InMux
    port map (
            O => \N__9042\,
            I => \N__9039\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__9039\,
            I => \N__9006\
        );

    \I__2007\ : ClkMux
    port map (
            O => \N__9038\,
            I => \N__8916\
        );

    \I__2006\ : ClkMux
    port map (
            O => \N__9037\,
            I => \N__8916\
        );

    \I__2005\ : ClkMux
    port map (
            O => \N__9036\,
            I => \N__8916\
        );

    \I__2004\ : ClkMux
    port map (
            O => \N__9035\,
            I => \N__8916\
        );

    \I__2003\ : ClkMux
    port map (
            O => \N__9034\,
            I => \N__8916\
        );

    \I__2002\ : ClkMux
    port map (
            O => \N__9033\,
            I => \N__8916\
        );

    \I__2001\ : ClkMux
    port map (
            O => \N__9032\,
            I => \N__8916\
        );

    \I__2000\ : ClkMux
    port map (
            O => \N__9031\,
            I => \N__8916\
        );

    \I__1999\ : ClkMux
    port map (
            O => \N__9030\,
            I => \N__8916\
        );

    \I__1998\ : ClkMux
    port map (
            O => \N__9029\,
            I => \N__8916\
        );

    \I__1997\ : ClkMux
    port map (
            O => \N__9028\,
            I => \N__8916\
        );

    \I__1996\ : ClkMux
    port map (
            O => \N__9027\,
            I => \N__8916\
        );

    \I__1995\ : ClkMux
    port map (
            O => \N__9026\,
            I => \N__8916\
        );

    \I__1994\ : ClkMux
    port map (
            O => \N__9025\,
            I => \N__8916\
        );

    \I__1993\ : ClkMux
    port map (
            O => \N__9024\,
            I => \N__8916\
        );

    \I__1992\ : ClkMux
    port map (
            O => \N__9023\,
            I => \N__8916\
        );

    \I__1991\ : ClkMux
    port map (
            O => \N__9022\,
            I => \N__8916\
        );

    \I__1990\ : ClkMux
    port map (
            O => \N__9021\,
            I => \N__8916\
        );

    \I__1989\ : ClkMux
    port map (
            O => \N__9020\,
            I => \N__8916\
        );

    \I__1988\ : ClkMux
    port map (
            O => \N__9019\,
            I => \N__8916\
        );

    \I__1987\ : ClkMux
    port map (
            O => \N__9018\,
            I => \N__8916\
        );

    \I__1986\ : ClkMux
    port map (
            O => \N__9017\,
            I => \N__8916\
        );

    \I__1985\ : ClkMux
    port map (
            O => \N__9016\,
            I => \N__8916\
        );

    \I__1984\ : ClkMux
    port map (
            O => \N__9015\,
            I => \N__8916\
        );

    \I__1983\ : ClkMux
    port map (
            O => \N__9014\,
            I => \N__8916\
        );

    \I__1982\ : ClkMux
    port map (
            O => \N__9013\,
            I => \N__8916\
        );

    \I__1981\ : ClkMux
    port map (
            O => \N__9012\,
            I => \N__8916\
        );

    \I__1980\ : ClkMux
    port map (
            O => \N__9011\,
            I => \N__8916\
        );

    \I__1979\ : ClkMux
    port map (
            O => \N__9010\,
            I => \N__8916\
        );

    \I__1978\ : ClkMux
    port map (
            O => \N__9009\,
            I => \N__8916\
        );

    \I__1977\ : Glb2LocalMux
    port map (
            O => \N__9006\,
            I => \N__8916\
        );

    \I__1976\ : ClkMux
    port map (
            O => \N__9005\,
            I => \N__8916\
        );

    \I__1975\ : ClkMux
    port map (
            O => \N__9004\,
            I => \N__8916\
        );

    \I__1974\ : ClkMux
    port map (
            O => \N__9003\,
            I => \N__8916\
        );

    \I__1973\ : ClkMux
    port map (
            O => \N__9002\,
            I => \N__8916\
        );

    \I__1972\ : ClkMux
    port map (
            O => \N__9001\,
            I => \N__8916\
        );

    \I__1971\ : ClkMux
    port map (
            O => \N__9000\,
            I => \N__8916\
        );

    \I__1970\ : ClkMux
    port map (
            O => \N__8999\,
            I => \N__8916\
        );

    \I__1969\ : ClkMux
    port map (
            O => \N__8998\,
            I => \N__8916\
        );

    \I__1968\ : ClkMux
    port map (
            O => \N__8997\,
            I => \N__8916\
        );

    \I__1967\ : GlobalMux
    port map (
            O => \N__8916\,
            I => \CLK80_PLL\
        );

    \I__1966\ : CEMux
    port map (
            O => \N__8913\,
            I => \N__8909\
        );

    \I__1965\ : CEMux
    port map (
            O => \N__8912\,
            I => \N__8904\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__8909\,
            I => \N__8901\
        );

    \I__1963\ : CEMux
    port map (
            O => \N__8908\,
            I => \N__8898\
        );

    \I__1962\ : CEMux
    port map (
            O => \N__8907\,
            I => \N__8895\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__8904\,
            I => \N__8892\
        );

    \I__1960\ : Span4Mux_v
    port map (
            O => \N__8901\,
            I => \N__8888\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__8898\,
            I => \N__8885\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__8895\,
            I => \N__8880\
        );

    \I__1957\ : Span4Mux_v
    port map (
            O => \N__8892\,
            I => \N__8880\
        );

    \I__1956\ : CEMux
    port map (
            O => \N__8891\,
            I => \N__8877\
        );

    \I__1955\ : Span4Mux_h
    port map (
            O => \N__8888\,
            I => \N__8872\
        );

    \I__1954\ : Span4Mux_v
    port map (
            O => \N__8885\,
            I => \N__8872\
        );

    \I__1953\ : Span4Mux_h
    port map (
            O => \N__8880\,
            I => \N__8869\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__8877\,
            I => \N__8866\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__8872\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__8869\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1949\ : Odrv12
    port map (
            O => \N__8866\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1948\ : InMux
    port map (
            O => \N__8859\,
            I => \N__8853\
        );

    \I__1947\ : InMux
    port map (
            O => \N__8858\,
            I => \N__8853\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__8853\,
            I => \N__8850\
        );

    \I__1945\ : Odrv12
    port map (
            O => \N__8850\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8844\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__8844\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1942\ : IoInMux
    port map (
            O => \N__8841\,
            I => \N__8838\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__8838\,
            I => \N__8835\
        );

    \I__1940\ : Span4Mux_s3_v
    port map (
            O => \N__8835\,
            I => \N__8832\
        );

    \I__1939\ : Span4Mux_v
    port map (
            O => \N__8832\,
            I => \N__8829\
        );

    \I__1938\ : Span4Mux_v
    port map (
            O => \N__8829\,
            I => \N__8826\
        );

    \I__1937\ : Span4Mux_h
    port map (
            O => \N__8826\,
            I => \N__8823\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__8823\,
            I => \CMA_c_0\
        );

    \I__1935\ : InMux
    port map (
            O => \N__8820\,
            I => \N__8817\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__8817\,
            I => \N__8813\
        );

    \I__1933\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8810\
        );

    \I__1932\ : Span4Mux_v
    port map (
            O => \N__8813\,
            I => \N__8804\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__8810\,
            I => \N__8804\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8809\,
            I => \N__8801\
        );

    \I__1929\ : Span4Mux_h
    port map (
            O => \N__8804\,
            I => \N__8796\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__8801\,
            I => \N__8796\
        );

    \I__1927\ : Span4Mux_v
    port map (
            O => \N__8796\,
            I => \N__8792\
        );

    \I__1926\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8789\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__8792\,
            I => \N__8786\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8789\,
            I => \N__8783\
        );

    \I__1923\ : Sp12to4
    port map (
            O => \N__8786\,
            I => \N__8778\
        );

    \I__1922\ : Span12Mux_v
    port map (
            O => \N__8783\,
            I => \N__8778\
        );

    \I__1921\ : Span12Mux_h
    port map (
            O => \N__8778\,
            I => \N__8775\
        );

    \I__1920\ : Odrv12
    port map (
            O => \N__8775\,
            I => \DRA_c_2\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8772\,
            I => \N__8769\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__8769\,
            I => \N__8766\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__8766\,
            I => \N__8763\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__8763\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1915\ : IoInMux
    port map (
            O => \N__8760\,
            I => \N__8757\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__8757\,
            I => \N__8754\
        );

    \I__1913\ : Span4Mux_s2_h
    port map (
            O => \N__8754\,
            I => \N__8751\
        );

    \I__1912\ : Sp12to4
    port map (
            O => \N__8751\,
            I => \N__8748\
        );

    \I__1911\ : Span12Mux_v
    port map (
            O => \N__8748\,
            I => \N__8745\
        );

    \I__1910\ : Span12Mux_h
    port map (
            O => \N__8745\,
            I => \N__8742\
        );

    \I__1909\ : Odrv12
    port map (
            O => \N__8742\,
            I => \N_295_i\
        );

    \I__1908\ : IoInMux
    port map (
            O => \N__8739\,
            I => \N__8736\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8736\,
            I => \N__8733\
        );

    \I__1906\ : Span4Mux_s2_h
    port map (
            O => \N__8733\,
            I => \N__8730\
        );

    \I__1905\ : Sp12to4
    port map (
            O => \N__8730\,
            I => \N__8727\
        );

    \I__1904\ : Span12Mux_s11_v
    port map (
            O => \N__8727\,
            I => \N__8724\
        );

    \I__1903\ : Span12Mux_h
    port map (
            O => \N__8724\,
            I => \N__8721\
        );

    \I__1902\ : Odrv12
    port map (
            O => \N__8721\,
            I => \N_299_i\
        );

    \I__1901\ : IoInMux
    port map (
            O => \N__8718\,
            I => \N__8715\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__8715\,
            I => \N__8712\
        );

    \I__1899\ : IoSpan4Mux
    port map (
            O => \N__8712\,
            I => \N__8709\
        );

    \I__1898\ : Span4Mux_s3_v
    port map (
            O => \N__8709\,
            I => \N__8703\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8696\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8707\,
            I => \N__8696\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8696\
        );

    \I__1894\ : Span4Mux_v
    port map (
            O => \N__8703\,
            I => \N__8693\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__8696\,
            I => \N__8690\
        );

    \I__1892\ : Sp12to4
    port map (
            O => \N__8693\,
            I => \N__8686\
        );

    \I__1891\ : Span4Mux_v
    port map (
            O => \N__8690\,
            I => \N__8683\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8689\,
            I => \N__8680\
        );

    \I__1889\ : Span12Mux_v
    port map (
            O => \N__8686\,
            I => \N__8672\
        );

    \I__1888\ : Sp12to4
    port map (
            O => \N__8683\,
            I => \N__8672\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8680\,
            I => \N__8672\
        );

    \I__1886\ : InMux
    port map (
            O => \N__8679\,
            I => \N__8669\
        );

    \I__1885\ : Odrv12
    port map (
            O => \N__8672\,
            I => \DBENn_c\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__8669\,
            I => \DBENn_c\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__8664\,
            I => \N__8659\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__8663\,
            I => \N__8656\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__8662\,
            I => \N__8652\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8659\,
            I => \N__8649\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8656\,
            I => \N__8644\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8644\
        );

    \I__1877\ : InMux
    port map (
            O => \N__8652\,
            I => \N__8641\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__8649\,
            I => \N__8635\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8644\,
            I => \N__8635\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__8641\,
            I => \N__8632\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8640\,
            I => \N__8629\
        );

    \I__1872\ : Span4Mux_h
    port map (
            O => \N__8635\,
            I => \N__8621\
        );

    \I__1871\ : Span4Mux_v
    port map (
            O => \N__8632\,
            I => \N__8621\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8629\,
            I => \N__8621\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8628\,
            I => \N__8615\
        );

    \I__1868\ : Span4Mux_h
    port map (
            O => \N__8621\,
            I => \N__8612\
        );

    \I__1867\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8609\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8604\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8618\,
            I => \N__8604\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8615\,
            I => \N__8601\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__8612\,
            I => \DMA_CYCLEm\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8609\,
            I => \DMA_CYCLEm\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8604\,
            I => \DMA_CYCLEm\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__8601\,
            I => \DMA_CYCLEm\
        );

    \I__1859\ : IoInMux
    port map (
            O => \N__8592\,
            I => \N__8589\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__8589\,
            I => \N__8586\
        );

    \I__1857\ : Span12Mux_s2_h
    port map (
            O => \N__8586\,
            I => \N__8583\
        );

    \I__1856\ : Span12Mux_h
    port map (
            O => \N__8583\,
            I => \N__8580\
        );

    \I__1855\ : Span12Mux_v
    port map (
            O => \N__8580\,
            I => \N__8577\
        );

    \I__1854\ : Odrv12
    port map (
            O => \N__8577\,
            I => \N_297_i\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8571\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__8571\,
            I => \U712_BYTE_ENABLE.N_528\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__8568\,
            I => \U712_BYTE_ENABLE.N_377_cascade_\
        );

    \I__1850\ : InMux
    port map (
            O => \N__8565\,
            I => \N__8562\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__1848\ : Odrv4
    port map (
            O => \N__8559\,
            I => \U712_BYTE_ENABLE.N_508\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8556\,
            I => \N__8553\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__8553\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1845\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8547\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__8547\,
            I => \N__8544\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__8544\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1842\ : InMux
    port map (
            O => \N__8541\,
            I => \N__8538\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8538\,
            I => \N__8535\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__8535\,
            I => \U712_CHIP_RAM.un3_DMA_CYCLE_START\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8532\,
            I => \N__8526\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8526\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__8526\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__8523\,
            I => \N__8512\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8507\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8507\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8520\,
            I => \N__8498\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8498\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8518\,
            I => \N__8489\
        );

    \I__1830\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8486\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8483\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8515\,
            I => \N__8476\
        );

    \I__1827\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8476\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__8507\,
            I => \N__8473\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8506\,
            I => \N__8470\
        );

    \I__1824\ : InMux
    port map (
            O => \N__8505\,
            I => \N__8467\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8504\,
            I => \N__8462\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8503\,
            I => \N__8462\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8498\,
            I => \N__8459\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8497\,
            I => \N__8456\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8453\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8448\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8494\,
            I => \N__8448\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8493\,
            I => \N__8443\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8443\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8489\,
            I => \N__8436\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8486\,
            I => \N__8436\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8483\,
            I => \N__8436\
        );

    \I__1811\ : InMux
    port map (
            O => \N__8482\,
            I => \N__8433\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8481\,
            I => \N__8422\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__8476\,
            I => \N__8419\
        );

    \I__1808\ : Span4Mux_h
    port map (
            O => \N__8473\,
            I => \N__8410\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8470\,
            I => \N__8410\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__8467\,
            I => \N__8410\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__8462\,
            I => \N__8410\
        );

    \I__1804\ : Span4Mux_v
    port map (
            O => \N__8459\,
            I => \N__8407\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8456\,
            I => \N__8404\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8453\,
            I => \N__8397\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8448\,
            I => \N__8397\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__8443\,
            I => \N__8397\
        );

    \I__1799\ : Sp12to4
    port map (
            O => \N__8436\,
            I => \N__8392\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8433\,
            I => \N__8392\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8432\,
            I => \N__8385\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8431\,
            I => \N__8385\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8385\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8378\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8428\,
            I => \N__8378\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8378\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8373\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8425\,
            I => \N__8373\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__8422\,
            I => \N__8370\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__8419\,
            I => \N__8365\
        );

    \I__1787\ : Span4Mux_v
    port map (
            O => \N__8410\,
            I => \N__8365\
        );

    \I__1786\ : Span4Mux_h
    port map (
            O => \N__8407\,
            I => \N__8358\
        );

    \I__1785\ : Span4Mux_v
    port map (
            O => \N__8404\,
            I => \N__8358\
        );

    \I__1784\ : Span4Mux_v
    port map (
            O => \N__8397\,
            I => \N__8358\
        );

    \I__1783\ : Span12Mux_v
    port map (
            O => \N__8392\,
            I => \N__8349\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8385\,
            I => \N__8349\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__8378\,
            I => \N__8349\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8373\,
            I => \N__8349\
        );

    \I__1779\ : Span12Mux_v
    port map (
            O => \N__8370\,
            I => \N__8342\
        );

    \I__1778\ : Sp12to4
    port map (
            O => \N__8365\,
            I => \N__8342\
        );

    \I__1777\ : Sp12to4
    port map (
            O => \N__8358\,
            I => \N__8342\
        );

    \I__1776\ : Span12Mux_h
    port map (
            O => \N__8349\,
            I => \N__8339\
        );

    \I__1775\ : Span12Mux_h
    port map (
            O => \N__8342\,
            I => \N__8336\
        );

    \I__1774\ : Odrv12
    port map (
            O => \N__8339\,
            I => \RESETn_c\
        );

    \I__1773\ : Odrv12
    port map (
            O => \N__8336\,
            I => \RESETn_c\
        );

    \I__1772\ : InMux
    port map (
            O => \N__8331\,
            I => \N__8328\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__8328\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8325\,
            I => \N__8322\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__8322\,
            I => \N__8319\
        );

    \I__1768\ : Span4Mux_v
    port map (
            O => \N__8319\,
            I => \N__8316\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__8316\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8313\,
            I => \N__8310\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__8310\,
            I => \N__8307\
        );

    \I__1764\ : Span4Mux_h
    port map (
            O => \N__8307\,
            I => \N__8304\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__8304\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1762\ : IoInMux
    port map (
            O => \N__8301\,
            I => \N__8298\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8298\,
            I => \N__8295\
        );

    \I__1760\ : IoSpan4Mux
    port map (
            O => \N__8295\,
            I => \N__8292\
        );

    \I__1759\ : Span4Mux_s3_h
    port map (
            O => \N__8292\,
            I => \N__8289\
        );

    \I__1758\ : Sp12to4
    port map (
            O => \N__8289\,
            I => \N__8286\
        );

    \I__1757\ : Span12Mux_h
    port map (
            O => \N__8286\,
            I => \N__8283\
        );

    \I__1756\ : Odrv12
    port map (
            O => \N__8283\,
            I => \CMA_c_3\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8276\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8273\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__8276\,
            I => \N__8268\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__8273\,
            I => \N__8265\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8272\,
            I => \N__8262\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8271\,
            I => \N__8259\
        );

    \I__1749\ : Span4Mux_v
    port map (
            O => \N__8268\,
            I => \N__8252\
        );

    \I__1748\ : Span4Mux_h
    port map (
            O => \N__8265\,
            I => \N__8252\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8262\,
            I => \N__8252\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__8259\,
            I => \N__8247\
        );

    \I__1745\ : Sp12to4
    port map (
            O => \N__8252\,
            I => \N__8247\
        );

    \I__1744\ : Span12Mux_v
    port map (
            O => \N__8247\,
            I => \N__8244\
        );

    \I__1743\ : Span12Mux_h
    port map (
            O => \N__8244\,
            I => \N__8241\
        );

    \I__1742\ : Odrv12
    port map (
            O => \N__8241\,
            I => \DRA_c_3\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8238\,
            I => \N__8235\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__8235\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1739\ : InMux
    port map (
            O => \N__8232\,
            I => \N__8228\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8231\,
            I => \N__8221\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__8228\,
            I => \N__8218\
        );

    \I__1736\ : InMux
    port map (
            O => \N__8227\,
            I => \N__8213\
        );

    \I__1735\ : InMux
    port map (
            O => \N__8226\,
            I => \N__8213\
        );

    \I__1734\ : InMux
    port map (
            O => \N__8225\,
            I => \N__8208\
        );

    \I__1733\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8208\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__8221\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__8218\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__8213\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8208\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__8199\,
            I => \N__8189\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8198\,
            I => \N__8180\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8197\,
            I => \N__8180\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8196\,
            I => \N__8180\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8175\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8194\,
            I => \N__8172\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8193\,
            I => \N__8169\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8192\,
            I => \N__8164\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8189\,
            I => \N__8164\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8188\,
            I => \N__8159\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8187\,
            I => \N__8159\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8180\,
            I => \N__8156\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8179\,
            I => \N__8151\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8178\,
            I => \N__8151\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8175\,
            I => \N__8148\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__8172\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__8169\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8164\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__8159\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__8156\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__8151\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__8148\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__8133\,
            I => \N__8129\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8132\,
            I => \N__8121\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8129\,
            I => \N__8118\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8128\,
            I => \N__8109\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8127\,
            I => \N__8109\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8126\,
            I => \N__8109\
        );

    \I__1700\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8109\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8106\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__8121\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__8118\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__8109\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8106\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8090\
        );

    \I__1693\ : InMux
    port map (
            O => \N__8096\,
            I => \N__8083\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8083\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8094\,
            I => \N__8078\
        );

    \I__1690\ : InMux
    port map (
            O => \N__8093\,
            I => \N__8078\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__8090\,
            I => \N__8075\
        );

    \I__1688\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8070\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8070\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8083\,
            I => \N__8067\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8078\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1684\ : Odrv12
    port map (
            O => \N__8075\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8070\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1682\ : Odrv4
    port map (
            O => \N__8067\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__8058\,
            I => \N__8055\
        );

    \I__1680\ : InMux
    port map (
            O => \N__8055\,
            I => \N__8052\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8052\,
            I => \U712_REG_SM.N_479\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__8049\,
            I => \N__8044\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8048\,
            I => \N__8038\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8047\,
            I => \N__8038\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8044\,
            I => \N__8035\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8043\,
            I => \N__8032\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__8038\,
            I => \N__8027\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8035\,
            I => \N__8027\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__8032\,
            I => \N__8024\
        );

    \I__1670\ : Span4Mux_v
    port map (
            O => \N__8027\,
            I => \N__8021\
        );

    \I__1669\ : Sp12to4
    port map (
            O => \N__8024\,
            I => \N__8018\
        );

    \I__1668\ : Sp12to4
    port map (
            O => \N__8021\,
            I => \N__8015\
        );

    \I__1667\ : Span12Mux_v
    port map (
            O => \N__8018\,
            I => \N__8010\
        );

    \I__1666\ : Span12Mux_h
    port map (
            O => \N__8015\,
            I => \N__8010\
        );

    \I__1665\ : Span12Mux_v
    port map (
            O => \N__8010\,
            I => \N__8007\
        );

    \I__1664\ : Odrv12
    port map (
            O => \N__8007\,
            I => \CLK40_PLL_i\
        );

    \I__1663\ : IoInMux
    port map (
            O => \N__8004\,
            I => \N__7999\
        );

    \I__1662\ : IoInMux
    port map (
            O => \N__8003\,
            I => \N__7996\
        );

    \I__1661\ : IoInMux
    port map (
            O => \N__8002\,
            I => \N__7993\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7999\,
            I => \N__7988\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__7996\,
            I => \N__7988\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__7993\,
            I => \N__7985\
        );

    \I__1657\ : IoSpan4Mux
    port map (
            O => \N__7988\,
            I => \N__7982\
        );

    \I__1656\ : Span4Mux_s3_h
    port map (
            O => \N__7985\,
            I => \N__7979\
        );

    \I__1655\ : Span4Mux_s1_v
    port map (
            O => \N__7982\,
            I => \N__7976\
        );

    \I__1654\ : Sp12to4
    port map (
            O => \N__7979\,
            I => \N__7973\
        );

    \I__1653\ : Sp12to4
    port map (
            O => \N__7976\,
            I => \N__7970\
        );

    \I__1652\ : Span12Mux_v
    port map (
            O => \N__7973\,
            I => \N__7967\
        );

    \I__1651\ : Span12Mux_h
    port map (
            O => \N__7970\,
            I => \N__7962\
        );

    \I__1650\ : Span12Mux_h
    port map (
            O => \N__7967\,
            I => \N__7962\
        );

    \I__1649\ : Odrv12
    port map (
            O => \N__7962\,
            I => \CLK40_PLL_i_i\
        );

    \I__1648\ : IoInMux
    port map (
            O => \N__7959\,
            I => \N__7956\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__7956\,
            I => \N__7953\
        );

    \I__1646\ : Span12Mux_s5_v
    port map (
            O => \N__7953\,
            I => \N__7950\
        );

    \I__1645\ : Odrv12
    port map (
            O => \N__7950\,
            I => \RESETn_c_i\
        );

    \I__1644\ : InMux
    port map (
            O => \N__7947\,
            I => \N__7944\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7944\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1642\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7938\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7938\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1640\ : InMux
    port map (
            O => \N__7935\,
            I => \N__7932\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__7932\,
            I => \N__7929\
        );

    \I__1638\ : Odrv4
    port map (
            O => \N__7929\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1637\ : InMux
    port map (
            O => \N__7926\,
            I => \N__7923\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__7923\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1635\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7917\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__7917\,
            I => \N__7914\
        );

    \I__1633\ : Span4Mux_h
    port map (
            O => \N__7914\,
            I => \N__7911\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__7911\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1631\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7905\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__7905\,
            I => \N__7902\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__7902\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7895\
        );

    \I__1627\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7892\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__7895\,
            I => \N__7889\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__7892\,
            I => \N__7886\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__7889\,
            I => \U712_REG_SM.N_661\
        );

    \I__1623\ : Odrv12
    port map (
            O => \N__7886\,
            I => \U712_REG_SM.N_661\
        );

    \I__1622\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7876\
        );

    \I__1621\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7873\
        );

    \I__1620\ : InMux
    port map (
            O => \N__7879\,
            I => \N__7870\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7876\,
            I => \U712_REG_SM.N_389\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__7873\,
            I => \U712_REG_SM.N_389\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__7870\,
            I => \U712_REG_SM.N_389\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__7863\,
            I => \U712_REG_SM.N_475_cascade_\
        );

    \I__1615\ : IoInMux
    port map (
            O => \N__7860\,
            I => \N__7857\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__7857\,
            I => \N__7854\
        );

    \I__1613\ : Span4Mux_s2_v
    port map (
            O => \N__7854\,
            I => \N__7851\
        );

    \I__1612\ : Span4Mux_h
    port map (
            O => \N__7851\,
            I => \N__7848\
        );

    \I__1611\ : Sp12to4
    port map (
            O => \N__7848\,
            I => \N__7845\
        );

    \I__1610\ : Span12Mux_s9_v
    port map (
            O => \N__7845\,
            I => \N__7842\
        );

    \I__1609\ : Odrv12
    port map (
            O => \N__7842\,
            I => \N_57_i\
        );

    \I__1608\ : InMux
    port map (
            O => \N__7839\,
            I => \N__7835\
        );

    \I__1607\ : InMux
    port map (
            O => \N__7838\,
            I => \N__7832\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__7835\,
            I => \N__7826\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__7832\,
            I => \N__7826\
        );

    \I__1604\ : InMux
    port map (
            O => \N__7831\,
            I => \N__7823\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__7826\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__7823\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7818\,
            I => \N__7815\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7815\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__7812\,
            I => \N__7809\
        );

    \I__1598\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7804\
        );

    \I__1597\ : InMux
    port map (
            O => \N__7808\,
            I => \N__7801\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7807\,
            I => \N__7798\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7804\,
            I => \N__7790\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__7801\,
            I => \N__7790\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__7798\,
            I => \N__7790\
        );

    \I__1592\ : InMux
    port map (
            O => \N__7797\,
            I => \N__7787\
        );

    \I__1591\ : Odrv4
    port map (
            O => \N__7790\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__7787\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__7782\,
            I => \U712_REG_SM.N_449_cascade_\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7779\,
            I => \N__7773\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7778\,
            I => \N__7773\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__7773\,
            I => \N__7766\
        );

    \I__1585\ : InMux
    port map (
            O => \N__7772\,
            I => \N__7763\
        );

    \I__1584\ : InMux
    port map (
            O => \N__7771\,
            I => \N__7758\
        );

    \I__1583\ : InMux
    port map (
            O => \N__7770\,
            I => \N__7758\
        );

    \I__1582\ : InMux
    port map (
            O => \N__7769\,
            I => \N__7755\
        );

    \I__1581\ : Span4Mux_h
    port map (
            O => \N__7766\,
            I => \N__7752\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__7763\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__7758\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__7755\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__7752\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__1576\ : InMux
    port map (
            O => \N__7743\,
            I => \N__7739\
        );

    \I__1575\ : InMux
    port map (
            O => \N__7742\,
            I => \N__7736\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__7739\,
            I => \U712_REG_SM.START_RST_0_sqmuxa\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7736\,
            I => \U712_REG_SM.START_RST_0_sqmuxa\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__7731\,
            I => \U712_REG_SM.N_396_cascade_\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__7728\,
            I => \N__7725\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7725\,
            I => \N__7720\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__7724\,
            I => \N__7717\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__7723\,
            I => \N__7713\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__7720\,
            I => \N__7709\
        );

    \I__1566\ : InMux
    port map (
            O => \N__7717\,
            I => \N__7702\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7716\,
            I => \N__7702\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7713\,
            I => \N__7702\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7712\,
            I => \N__7697\
        );

    \I__1562\ : Span4Mux_v
    port map (
            O => \N__7709\,
            I => \N__7690\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7702\,
            I => \N__7690\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7701\,
            I => \N__7685\
        );

    \I__1559\ : InMux
    port map (
            O => \N__7700\,
            I => \N__7682\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7697\,
            I => \N__7679\
        );

    \I__1557\ : InMux
    port map (
            O => \N__7696\,
            I => \N__7676\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7695\,
            I => \N__7673\
        );

    \I__1555\ : Span4Mux_h
    port map (
            O => \N__7690\,
            I => \N__7670\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7689\,
            I => \N__7665\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7688\,
            I => \N__7665\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7685\,
            I => \N__7662\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7682\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1550\ : Odrv4
    port map (
            O => \N__7679\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7676\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7673\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__7670\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__7665\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1545\ : Odrv4
    port map (
            O => \N__7662\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7647\,
            I => \N__7644\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__7644\,
            I => \U712_REG_SM.un1_STATE_COUNT_4_i_i_0_0\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7641\,
            I => \N__7637\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7634\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7637\,
            I => \N__7631\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__7634\,
            I => \N__7628\
        );

    \I__1538\ : Span4Mux_v
    port map (
            O => \N__7631\,
            I => \N__7623\
        );

    \I__1537\ : Span4Mux_v
    port map (
            O => \N__7628\,
            I => \N__7623\
        );

    \I__1536\ : Span4Mux_v
    port map (
            O => \N__7623\,
            I => \N__7620\
        );

    \I__1535\ : Sp12to4
    port map (
            O => \N__7620\,
            I => \N__7617\
        );

    \I__1534\ : Span12Mux_h
    port map (
            O => \N__7617\,
            I => \N__7614\
        );

    \I__1533\ : Odrv12
    port map (
            O => \N__7614\,
            I => \TSn_c\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__7611\,
            I => \U712_REG_SM.N_477_cascade_\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7608\,
            I => \N__7605\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7605\,
            I => \N__7602\
        );

    \I__1529\ : Span4Mux_v
    port map (
            O => \N__7602\,
            I => \N__7599\
        );

    \I__1528\ : Sp12to4
    port map (
            O => \N__7599\,
            I => \N__7596\
        );

    \I__1527\ : Span12Mux_h
    port map (
            O => \N__7596\,
            I => \N__7593\
        );

    \I__1526\ : Span12Mux_v
    port map (
            O => \N__7593\,
            I => \N__7590\
        );

    \I__1525\ : Odrv12
    port map (
            O => \N__7590\,
            I => \REGSPACEn_c\
        );

    \I__1524\ : IoInMux
    port map (
            O => \N__7587\,
            I => \N__7584\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7584\,
            I => \N__7581\
        );

    \I__1522\ : Span4Mux_s0_v
    port map (
            O => \N__7581\,
            I => \N__7578\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__7578\,
            I => \N__7574\
        );

    \I__1520\ : InMux
    port map (
            O => \N__7577\,
            I => \N__7571\
        );

    \I__1519\ : Span4Mux_v
    port map (
            O => \N__7574\,
            I => \N__7568\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7571\,
            I => \N__7565\
        );

    \I__1517\ : Sp12to4
    port map (
            O => \N__7568\,
            I => \N__7562\
        );

    \I__1516\ : Span4Mux_v
    port map (
            O => \N__7565\,
            I => \N__7559\
        );

    \I__1515\ : Span12Mux_h
    port map (
            O => \N__7562\,
            I => \N__7556\
        );

    \I__1514\ : Sp12to4
    port map (
            O => \N__7559\,
            I => \N__7553\
        );

    \I__1513\ : Span12Mux_v
    port map (
            O => \N__7556\,
            I => \N__7548\
        );

    \I__1512\ : Span12Mux_h
    port map (
            O => \N__7553\,
            I => \N__7548\
        );

    \I__1511\ : Odrv12
    port map (
            O => \N__7548\,
            I => \A_c_10\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7542\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__7542\,
            I => \N__7539\
        );

    \I__1508\ : Odrv4
    port map (
            O => \N__7539\,
            I => \U712_CHIP_RAM.N_422\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7536\,
            I => \N__7533\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7533\,
            I => \N__7530\
        );

    \I__1505\ : Span4Mux_v
    port map (
            O => \N__7530\,
            I => \N__7527\
        );

    \I__1504\ : Sp12to4
    port map (
            O => \N__7527\,
            I => \N__7524\
        );

    \I__1503\ : Span12Mux_h
    port map (
            O => \N__7524\,
            I => \N__7521\
        );

    \I__1502\ : Span12Mux_v
    port map (
            O => \N__7521\,
            I => \N__7518\
        );

    \I__1501\ : Odrv12
    port map (
            O => \N__7518\,
            I => \A_c_3\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7515\,
            I => \N__7512\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__7512\,
            I => \N__7509\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__7509\,
            I => \U712_CHIP_RAM.N_445\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7503\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__7503\,
            I => \N__7500\
        );

    \I__1495\ : Span4Mux_h
    port map (
            O => \N__7500\,
            I => \N__7496\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7499\,
            I => \N__7493\
        );

    \I__1493\ : Span4Mux_h
    port map (
            O => \N__7496\,
            I => \N__7488\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7493\,
            I => \N__7488\
        );

    \I__1491\ : Span4Mux_v
    port map (
            O => \N__7488\,
            I => \N__7485\
        );

    \I__1490\ : Span4Mux_h
    port map (
            O => \N__7485\,
            I => \N__7482\
        );

    \I__1489\ : Sp12to4
    port map (
            O => \N__7482\,
            I => \N__7479\
        );

    \I__1488\ : Odrv12
    port map (
            O => \N__7479\,
            I => \DBRn_c\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7476\,
            I => \N__7473\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7473\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7470\,
            I => \N__7466\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7469\,
            I => \N__7463\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7466\,
            I => \N__7460\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7463\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__7460\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7455\,
            I => \N__7452\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7452\,
            I => \N__7449\
        );

    \I__1478\ : Span4Mux_h
    port map (
            O => \N__7449\,
            I => \N__7446\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__7446\,
            I => \U712_CYCLE_TERM.TACK_EN_RNOZ0Z_0\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7443\,
            I => \N__7439\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7442\,
            I => \N__7436\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7439\,
            I => \N__7433\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7436\,
            I => \N__7428\
        );

    \I__1472\ : Span4Mux_h
    port map (
            O => \N__7433\,
            I => \N__7428\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__7428\,
            I => \U712_CYCLE_TERM.un13_0\
        );

    \I__1470\ : IoInMux
    port map (
            O => \N__7425\,
            I => \N__7422\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__7422\,
            I => \N__7419\
        );

    \I__1468\ : IoSpan4Mux
    port map (
            O => \N__7419\,
            I => \N__7415\
        );

    \I__1467\ : IoInMux
    port map (
            O => \N__7418\,
            I => \N__7412\
        );

    \I__1466\ : Span4Mux_s1_v
    port map (
            O => \N__7415\,
            I => \N__7409\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7412\,
            I => \N__7406\
        );

    \I__1464\ : Span4Mux_v
    port map (
            O => \N__7409\,
            I => \N__7403\
        );

    \I__1463\ : IoSpan4Mux
    port map (
            O => \N__7406\,
            I => \N__7400\
        );

    \I__1462\ : Span4Mux_v
    port map (
            O => \N__7403\,
            I => \N__7397\
        );

    \I__1461\ : Span4Mux_s2_h
    port map (
            O => \N__7400\,
            I => \N__7393\
        );

    \I__1460\ : Span4Mux_v
    port map (
            O => \N__7397\,
            I => \N__7390\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7396\,
            I => \N__7387\
        );

    \I__1458\ : Sp12to4
    port map (
            O => \N__7393\,
            I => \N__7384\
        );

    \I__1457\ : Span4Mux_h
    port map (
            O => \N__7390\,
            I => \N__7379\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7387\,
            I => \N__7379\
        );

    \I__1455\ : Span12Mux_h
    port map (
            O => \N__7384\,
            I => \N__7376\
        );

    \I__1454\ : Span4Mux_v
    port map (
            O => \N__7379\,
            I => \N__7373\
        );

    \I__1453\ : Span12Mux_v
    port map (
            O => \N__7376\,
            I => \N__7369\
        );

    \I__1452\ : Span4Mux_h
    port map (
            O => \N__7373\,
            I => \N__7366\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7372\,
            I => \N__7363\
        );

    \I__1450\ : Odrv12
    port map (
            O => \N__7369\,
            I => \TACK_EN\
        );

    \I__1449\ : Odrv4
    port map (
            O => \N__7366\,
            I => \TACK_EN\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7363\,
            I => \TACK_EN\
        );

    \I__1447\ : IoInMux
    port map (
            O => \N__7356\,
            I => \N__7353\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7353\,
            I => \N__7350\
        );

    \I__1445\ : IoSpan4Mux
    port map (
            O => \N__7350\,
            I => \N__7347\
        );

    \I__1444\ : IoSpan4Mux
    port map (
            O => \N__7347\,
            I => \N__7344\
        );

    \I__1443\ : Sp12to4
    port map (
            O => \N__7344\,
            I => \N__7341\
        );

    \I__1442\ : Span12Mux_s7_v
    port map (
            O => \N__7341\,
            I => \N__7338\
        );

    \I__1441\ : Span12Mux_h
    port map (
            O => \N__7338\,
            I => \N__7335\
        );

    \I__1440\ : Odrv12
    port map (
            O => \N__7335\,
            I => \WEn_c\
        );

    \I__1439\ : IoInMux
    port map (
            O => \N__7332\,
            I => \N__7329\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__7329\,
            I => \N__7326\
        );

    \I__1437\ : Span4Mux_s0_v
    port map (
            O => \N__7326\,
            I => \N__7323\
        );

    \I__1436\ : Sp12to4
    port map (
            O => \N__7323\,
            I => \N__7320\
        );

    \I__1435\ : Span12Mux_h
    port map (
            O => \N__7320\,
            I => \N__7317\
        );

    \I__1434\ : Odrv12
    port map (
            O => \N__7317\,
            I => \CRCSn_c\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7314\,
            I => \N__7311\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7311\,
            I => \N__7308\
        );

    \I__1431\ : Sp12to4
    port map (
            O => \N__7308\,
            I => \N__7305\
        );

    \I__1430\ : Span12Mux_v
    port map (
            O => \N__7305\,
            I => \N__7302\
        );

    \I__1429\ : Span12Mux_h
    port map (
            O => \N__7302\,
            I => \N__7299\
        );

    \I__1428\ : Odrv12
    port map (
            O => \N__7299\,
            I => \A_c_19\
        );

    \I__1427\ : IoInMux
    port map (
            O => \N__7296\,
            I => \N__7293\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__7293\,
            I => \N__7290\
        );

    \I__1425\ : IoSpan4Mux
    port map (
            O => \N__7290\,
            I => \N__7287\
        );

    \I__1424\ : Span4Mux_s3_h
    port map (
            O => \N__7287\,
            I => \N__7284\
        );

    \I__1423\ : Span4Mux_v
    port map (
            O => \N__7284\,
            I => \N__7281\
        );

    \I__1422\ : Span4Mux_h
    port map (
            O => \N__7281\,
            I => \N__7278\
        );

    \I__1421\ : Sp12to4
    port map (
            O => \N__7278\,
            I => \N__7275\
        );

    \I__1420\ : Odrv12
    port map (
            O => \N__7275\,
            I => \CMA_c_9\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7272\,
            I => \N__7269\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__7269\,
            I => \N__7266\
        );

    \I__1417\ : Span12Mux_v
    port map (
            O => \N__7266\,
            I => \N__7263\
        );

    \I__1416\ : Span12Mux_h
    port map (
            O => \N__7263\,
            I => \N__7260\
        );

    \I__1415\ : Odrv12
    port map (
            O => \N__7260\,
            I => \A_c_17\
        );

    \I__1414\ : IoInMux
    port map (
            O => \N__7257\,
            I => \N__7254\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__7254\,
            I => \N__7251\
        );

    \I__1412\ : Span4Mux_s0_h
    port map (
            O => \N__7251\,
            I => \N__7248\
        );

    \I__1411\ : Span4Mux_h
    port map (
            O => \N__7248\,
            I => \N__7245\
        );

    \I__1410\ : Sp12to4
    port map (
            O => \N__7245\,
            I => \N__7242\
        );

    \I__1409\ : Span12Mux_s10_v
    port map (
            O => \N__7242\,
            I => \N__7239\
        );

    \I__1408\ : Span12Mux_h
    port map (
            O => \N__7239\,
            I => \N__7236\
        );

    \I__1407\ : Odrv12
    port map (
            O => \N__7236\,
            I => \CMA_c_8\
        );

    \I__1406\ : IoInMux
    port map (
            O => \N__7233\,
            I => \N__7230\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7230\,
            I => \N__7227\
        );

    \I__1404\ : Span12Mux_s11_v
    port map (
            O => \N__7227\,
            I => \N__7224\
        );

    \I__1403\ : Odrv12
    port map (
            O => \N__7224\,
            I => \CMA_c_1\
        );

    \I__1402\ : InMux
    port map (
            O => \N__7221\,
            I => \N__7217\
        );

    \I__1401\ : InMux
    port map (
            O => \N__7220\,
            I => \N__7213\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7217\,
            I => \N__7209\
        );

    \I__1399\ : InMux
    port map (
            O => \N__7216\,
            I => \N__7206\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__7213\,
            I => \N__7203\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__7212\,
            I => \N__7199\
        );

    \I__1396\ : Span4Mux_h
    port map (
            O => \N__7209\,
            I => \N__7196\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7206\,
            I => \N__7191\
        );

    \I__1394\ : Span4Mux_h
    port map (
            O => \N__7203\,
            I => \N__7191\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7202\,
            I => \N__7186\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7199\,
            I => \N__7186\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__7196\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__7191\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__7186\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1388\ : IoInMux
    port map (
            O => \N__7179\,
            I => \N__7176\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7176\,
            I => \N__7173\
        );

    \I__1386\ : Span4Mux_s1_v
    port map (
            O => \N__7173\,
            I => \N__7170\
        );

    \I__1385\ : Span4Mux_v
    port map (
            O => \N__7170\,
            I => \N__7167\
        );

    \I__1384\ : Sp12to4
    port map (
            O => \N__7167\,
            I => \N__7164\
        );

    \I__1383\ : Span12Mux_h
    port map (
            O => \N__7164\,
            I => \N__7161\
        );

    \I__1382\ : Odrv12
    port map (
            O => \N__7161\,
            I => \CMA_c_10\
        );

    \I__1381\ : IoInMux
    port map (
            O => \N__7158\,
            I => \N__7155\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7155\,
            I => \N__7152\
        );

    \I__1379\ : IoSpan4Mux
    port map (
            O => \N__7152\,
            I => \N__7149\
        );

    \I__1378\ : Sp12to4
    port map (
            O => \N__7149\,
            I => \N__7146\
        );

    \I__1377\ : Span12Mux_s7_v
    port map (
            O => \N__7146\,
            I => \N__7143\
        );

    \I__1376\ : Odrv12
    port map (
            O => \N__7143\,
            I => \CMA_c_2\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7137\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7137\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7134\,
            I => \N__7131\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7131\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1371\ : InMux
    port map (
            O => \N__7128\,
            I => \N__7125\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__7125\,
            I => \N__7122\
        );

    \I__1369\ : Span4Mux_h
    port map (
            O => \N__7122\,
            I => \N__7117\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7121\,
            I => \N__7114\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7120\,
            I => \N__7110\
        );

    \I__1366\ : Span4Mux_v
    port map (
            O => \N__7117\,
            I => \N__7107\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__7114\,
            I => \N__7104\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7113\,
            I => \N__7101\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__7110\,
            I => \N__7094\
        );

    \I__1362\ : Span4Mux_v
    port map (
            O => \N__7107\,
            I => \N__7094\
        );

    \I__1361\ : Span4Mux_h
    port map (
            O => \N__7104\,
            I => \N__7091\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__7101\,
            I => \N__7088\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7085\
        );

    \I__1358\ : InMux
    port map (
            O => \N__7099\,
            I => \N__7082\
        );

    \I__1357\ : Odrv4
    port map (
            O => \N__7094\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1356\ : Odrv4
    port map (
            O => \N__7091\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__7088\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7085\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__7082\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1352\ : InMux
    port map (
            O => \N__7071\,
            I => \N__7067\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__7070\,
            I => \N__7062\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__7067\,
            I => \N__7059\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7066\,
            I => \N__7056\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7065\,
            I => \N__7053\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7062\,
            I => \N__7049\
        );

    \I__1346\ : Span4Mux_v
    port map (
            O => \N__7059\,
            I => \N__7044\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__7056\,
            I => \N__7044\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7053\,
            I => \N__7041\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7052\,
            I => \N__7038\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7049\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1341\ : Odrv4
    port map (
            O => \N__7044\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1340\ : Odrv4
    port map (
            O => \N__7041\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__7038\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7029\,
            I => \N__7023\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7028\,
            I => \N__7023\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7023\,
            I => \U712_CHIP_RAM.CMA_5_i_0_8\
        );

    \I__1335\ : CascadeMux
    port map (
            O => \N__7020\,
            I => \U712_REG_SM.N_374_cascade_\
        );

    \I__1334\ : InMux
    port map (
            O => \N__7017\,
            I => \N__7014\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__7014\,
            I => \U712_REG_SM.N_417\
        );

    \I__1332\ : IoInMux
    port map (
            O => \N__7011\,
            I => \N__7008\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__7008\,
            I => \N__7005\
        );

    \I__1330\ : IoSpan4Mux
    port map (
            O => \N__7005\,
            I => \N__7002\
        );

    \I__1329\ : Span4Mux_s3_h
    port map (
            O => \N__7002\,
            I => \N__6999\
        );

    \I__1328\ : Span4Mux_v
    port map (
            O => \N__6999\,
            I => \N__6996\
        );

    \I__1327\ : Span4Mux_h
    port map (
            O => \N__6996\,
            I => \N__6993\
        );

    \I__1326\ : Sp12to4
    port map (
            O => \N__6993\,
            I => \N__6989\
        );

    \I__1325\ : InMux
    port map (
            O => \N__6992\,
            I => \N__6986\
        );

    \I__1324\ : Span12Mux_h
    port map (
            O => \N__6989\,
            I => \N__6981\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__6986\,
            I => \N__6981\
        );

    \I__1322\ : Span12Mux_h
    port map (
            O => \N__6981\,
            I => \N__6978\
        );

    \I__1321\ : Odrv12
    port map (
            O => \N__6978\,
            I => \C3_c\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6975\,
            I => \N__6972\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6972\,
            I => \U712_REG_SM.DS_EN_RNOZ0Z_0\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6969\,
            I => \N__6966\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6966\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6963\,
            I => \N__6959\
        );

    \I__1315\ : IoInMux
    port map (
            O => \N__6962\,
            I => \N__6956\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__6959\,
            I => \N__6953\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6956\,
            I => \N__6950\
        );

    \I__1312\ : Sp12to4
    port map (
            O => \N__6953\,
            I => \N__6947\
        );

    \I__1311\ : IoSpan4Mux
    port map (
            O => \N__6950\,
            I => \N__6944\
        );

    \I__1310\ : Span12Mux_v
    port map (
            O => \N__6947\,
            I => \N__6941\
        );

    \I__1309\ : IoSpan4Mux
    port map (
            O => \N__6944\,
            I => \N__6938\
        );

    \I__1308\ : Span12Mux_h
    port map (
            O => \N__6941\,
            I => \N__6935\
        );

    \I__1307\ : IoSpan4Mux
    port map (
            O => \N__6938\,
            I => \N__6932\
        );

    \I__1306\ : Odrv12
    port map (
            O => \N__6935\,
            I => \C1_c\
        );

    \I__1305\ : Odrv4
    port map (
            O => \N__6932\,
            I => \C1_c\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6927\,
            I => \N__6924\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6924\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1302\ : IoInMux
    port map (
            O => \N__6921\,
            I => \N__6918\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__6918\,
            I => \N__6915\
        );

    \I__1300\ : Span4Mux_s3_v
    port map (
            O => \N__6915\,
            I => \N__6912\
        );

    \I__1299\ : Span4Mux_v
    port map (
            O => \N__6912\,
            I => \N__6909\
        );

    \I__1298\ : Sp12to4
    port map (
            O => \N__6909\,
            I => \N__6906\
        );

    \I__1297\ : Odrv12
    port map (
            O => \N__6906\,
            I => \RASn_c\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6903\,
            I => \N__6893\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__6902\,
            I => \N__6890\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6901\,
            I => \N__6885\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6885\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__6899\,
            I => \N__6882\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6898\,
            I => \N__6878\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6897\,
            I => \N__6875\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6896\,
            I => \N__6872\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6893\,
            I => \N__6869\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6890\,
            I => \N__6866\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__6885\,
            I => \N__6863\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6882\,
            I => \N__6858\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6855\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6878\,
            I => \N__6852\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__6875\,
            I => \N__6847\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6872\,
            I => \N__6847\
        );

    \I__1280\ : Span4Mux_h
    port map (
            O => \N__6869\,
            I => \N__6844\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6866\,
            I => \N__6839\
        );

    \I__1278\ : Span4Mux_h
    port map (
            O => \N__6863\,
            I => \N__6839\
        );

    \I__1277\ : InMux
    port map (
            O => \N__6862\,
            I => \N__6836\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6861\,
            I => \N__6833\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6858\,
            I => \N__6824\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__6855\,
            I => \N__6824\
        );

    \I__1273\ : Span4Mux_v
    port map (
            O => \N__6852\,
            I => \N__6824\
        );

    \I__1272\ : Span4Mux_v
    port map (
            O => \N__6847\,
            I => \N__6824\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__6844\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__6839\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__6836\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6833\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__6824\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6813\,
            I => \N__6803\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6812\,
            I => \N__6796\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6811\,
            I => \N__6796\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6810\,
            I => \N__6796\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6809\,
            I => \N__6793\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__6808\,
            I => \N__6786\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6807\,
            I => \N__6781\
        );

    \I__1259\ : InMux
    port map (
            O => \N__6806\,
            I => \N__6778\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__6803\,
            I => \N__6775\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6796\,
            I => \N__6769\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__6793\,
            I => \N__6769\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6792\,
            I => \N__6762\
        );

    \I__1254\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6757\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6790\,
            I => \N__6757\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6789\,
            I => \N__6754\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6786\,
            I => \N__6749\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6785\,
            I => \N__6749\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6784\,
            I => \N__6746\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6781\,
            I => \N__6743\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6778\,
            I => \N__6740\
        );

    \I__1246\ : Span4Mux_v
    port map (
            O => \N__6775\,
            I => \N__6737\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6734\
        );

    \I__1244\ : Span4Mux_h
    port map (
            O => \N__6769\,
            I => \N__6731\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6728\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6767\,
            I => \N__6721\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6766\,
            I => \N__6721\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6721\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__6762\,
            I => \N__6714\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6757\,
            I => \N__6714\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6754\,
            I => \N__6714\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6749\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6746\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1234\ : Odrv4
    port map (
            O => \N__6743\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1233\ : Odrv4
    port map (
            O => \N__6740\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1232\ : Odrv4
    port map (
            O => \N__6737\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__6734\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1230\ : Odrv4
    port map (
            O => \N__6731\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__6728\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__6721\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1227\ : Odrv12
    port map (
            O => \N__6714\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__6693\,
            I => \N__6684\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__6692\,
            I => \N__6681\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6675\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6690\,
            I => \N__6672\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6689\,
            I => \N__6667\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6688\,
            I => \N__6667\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6687\,
            I => \N__6660\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6684\,
            I => \N__6660\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6681\,
            I => \N__6660\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__6680\,
            I => \N__6654\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6648\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6678\,
            I => \N__6645\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6675\,
            I => \N__6642\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__6672\,
            I => \N__6639\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6667\,
            I => \N__6634\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6660\,
            I => \N__6634\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6659\,
            I => \N__6631\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6658\,
            I => \N__6626\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6657\,
            I => \N__6626\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6654\,
            I => \N__6619\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6619\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6652\,
            I => \N__6619\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6616\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6648\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__6645\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__6642\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1200\ : Odrv4
    port map (
            O => \N__6639\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1199\ : Odrv4
    port map (
            O => \N__6634\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6631\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6626\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__6619\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__6616\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__6597\,
            I => \N__6591\
        );

    \I__1193\ : CascadeMux
    port map (
            O => \N__6596\,
            I => \N__6588\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6583\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6580\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6591\,
            I => \N__6572\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6588\,
            I => \N__6572\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__6587\,
            I => \N__6568\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6562\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6583\,
            I => \N__6557\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6580\,
            I => \N__6557\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6579\,
            I => \N__6554\
        );

    \I__1183\ : InMux
    port map (
            O => \N__6578\,
            I => \N__6551\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__6577\,
            I => \N__6548\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6572\,
            I => \N__6543\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6540\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6568\,
            I => \N__6533\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6567\,
            I => \N__6533\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6566\,
            I => \N__6533\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6565\,
            I => \N__6530\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6562\,
            I => \N__6527\
        );

    \I__1174\ : Span4Mux_v
    port map (
            O => \N__6557\,
            I => \N__6520\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__6554\,
            I => \N__6520\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6551\,
            I => \N__6520\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6548\,
            I => \N__6513\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6513\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6546\,
            I => \N__6513\
        );

    \I__1168\ : Odrv4
    port map (
            O => \N__6543\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__6540\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6533\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6530\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1164\ : Odrv4
    port map (
            O => \N__6527\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__6520\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__6513\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6495\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__6495\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_a2_0_0\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6489\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6489\,
            I => \N__6486\
        );

    \I__1157\ : Span4Mux_v
    port map (
            O => \N__6486\,
            I => \N__6482\
        );

    \I__1156\ : IoInMux
    port map (
            O => \N__6485\,
            I => \N__6479\
        );

    \I__1155\ : Span4Mux_h
    port map (
            O => \N__6482\,
            I => \N__6476\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6479\,
            I => \N__6473\
        );

    \I__1153\ : Sp12to4
    port map (
            O => \N__6476\,
            I => \N__6470\
        );

    \I__1152\ : IoSpan4Mux
    port map (
            O => \N__6473\,
            I => \N__6467\
        );

    \I__1151\ : Odrv12
    port map (
            O => \N__6470\,
            I => \RAMENn_c\
        );

    \I__1150\ : Odrv4
    port map (
            O => \N__6467\,
            I => \RAMENn_c\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__6462\,
            I => \U712_CHIP_RAM.N_492_cascade_\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6459\,
            I => \N__6454\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6458\,
            I => \N__6449\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6457\,
            I => \N__6449\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6454\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6449\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__6444\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_0_0_a2_0_0_0_cascade_\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6441\,
            I => \N__6438\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__6438\,
            I => \U712_REG_SM.N_374\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6435\,
            I => \N__6432\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6432\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_a2_1_0\
        );

    \I__1138\ : IoInMux
    port map (
            O => \N__6429\,
            I => \N__6426\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6426\,
            I => \N__6423\
        );

    \I__1136\ : Span12Mux_s4_v
    port map (
            O => \N__6423\,
            I => \N__6419\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6422\,
            I => \N__6416\
        );

    \I__1134\ : Span12Mux_h
    port map (
            O => \N__6419\,
            I => \N__6413\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6416\,
            I => \N__6410\
        );

    \I__1132\ : Span12Mux_v
    port map (
            O => \N__6413\,
            I => \N__6407\
        );

    \I__1131\ : Span12Mux_h
    port map (
            O => \N__6410\,
            I => \N__6404\
        );

    \I__1130\ : Odrv12
    port map (
            O => \N__6407\,
            I => \A_c_9\
        );

    \I__1129\ : Odrv12
    port map (
            O => \N__6404\,
            I => \A_c_9\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6399\,
            I => \N__6396\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__6396\,
            I => \N__6393\
        );

    \I__1126\ : Sp12to4
    port map (
            O => \N__6393\,
            I => \N__6390\
        );

    \I__1125\ : Span12Mux_v
    port map (
            O => \N__6390\,
            I => \N__6387\
        );

    \I__1124\ : Span12Mux_h
    port map (
            O => \N__6387\,
            I => \N__6384\
        );

    \I__1123\ : Odrv12
    port map (
            O => \N__6384\,
            I => \A_c_2\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6381\,
            I => \N__6378\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6378\,
            I => \N__6374\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6377\,
            I => \N__6371\
        );

    \I__1119\ : Span4Mux_h
    port map (
            O => \N__6374\,
            I => \N__6368\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6371\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__6368\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6363\,
            I => \N__6360\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__6360\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6354\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__6354\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6351\,
            I => \N__6347\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6350\,
            I => \N__6344\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6347\,
            I => \N__6341\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6344\,
            I => \N__6337\
        );

    \I__1108\ : Span4Mux_h
    port map (
            O => \N__6341\,
            I => \N__6334\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6340\,
            I => \N__6331\
        );

    \I__1106\ : Odrv4
    port map (
            O => \N__6337\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1105\ : Odrv4
    port map (
            O => \N__6334\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6331\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__6324\,
            I => \N__6320\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__6323\,
            I => \N__6317\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6320\,
            I => \N__6314\
        );

    \I__1100\ : InMux
    port map (
            O => \N__6317\,
            I => \N__6311\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6314\,
            I => \N__6308\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__6311\,
            I => \N__6305\
        );

    \I__1097\ : Span4Mux_v
    port map (
            O => \N__6308\,
            I => \N__6302\
        );

    \I__1096\ : Span4Mux_h
    port map (
            O => \N__6305\,
            I => \N__6299\
        );

    \I__1095\ : Odrv4
    port map (
            O => \N__6302\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1094\ : Odrv4
    port map (
            O => \N__6299\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1093\ : InMux
    port map (
            O => \N__6294\,
            I => \N__6290\
        );

    \I__1092\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6287\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__6290\,
            I => \N__6281\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__6287\,
            I => \N__6281\
        );

    \I__1089\ : InMux
    port map (
            O => \N__6286\,
            I => \N__6278\
        );

    \I__1088\ : Span4Mux_h
    port map (
            O => \N__6281\,
            I => \N__6274\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__6278\,
            I => \N__6271\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6277\,
            I => \N__6268\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__6274\,
            I => \U712_CHIP_RAM.N_567\
        );

    \I__1084\ : Odrv4
    port map (
            O => \N__6271\,
            I => \U712_CHIP_RAM.N_567\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__6268\,
            I => \U712_CHIP_RAM.N_567\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6261\,
            I => \N__6256\
        );

    \I__1081\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6251\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6259\,
            I => \N__6251\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6256\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6251\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__6246\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_1_cascade_\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6240\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6240\,
            I => \N__6235\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6239\,
            I => \N__6232\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6238\,
            I => \N__6229\
        );

    \I__1072\ : Span4Mux_h
    port map (
            O => \N__6235\,
            I => \N__6219\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__6232\,
            I => \N__6219\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__6229\,
            I => \N__6219\
        );

    \I__1069\ : InMux
    port map (
            O => \N__6228\,
            I => \N__6216\
        );

    \I__1068\ : InMux
    port map (
            O => \N__6227\,
            I => \N__6213\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6226\,
            I => \N__6210\
        );

    \I__1066\ : Odrv4
    port map (
            O => \N__6219\,
            I => \U712_CHIP_RAM.N_562\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__6216\,
            I => \U712_CHIP_RAM.N_562\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__6213\,
            I => \U712_CHIP_RAM.N_562\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__6210\,
            I => \U712_CHIP_RAM.N_562\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6197\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6200\,
            I => \N__6194\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6197\,
            I => \N__6191\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6194\,
            I => \U712_CHIP_RAM.N_502\
        );

    \I__1058\ : Odrv4
    port map (
            O => \N__6191\,
            I => \U712_CHIP_RAM.N_502\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__6186\,
            I => \N__6182\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__6185\,
            I => \N__6179\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6182\,
            I => \N__6174\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6179\,
            I => \N__6171\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__6178\,
            I => \N__6168\
        );

    \I__1052\ : InMux
    port map (
            O => \N__6177\,
            I => \N__6165\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6174\,
            I => \N__6160\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6171\,
            I => \N__6157\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6168\,
            I => \N__6154\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__6165\,
            I => \N__6151\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6164\,
            I => \N__6148\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6163\,
            I => \N__6141\
        );

    \I__1045\ : Span4Mux_v
    port map (
            O => \N__6160\,
            I => \N__6136\
        );

    \I__1044\ : Span4Mux_v
    port map (
            O => \N__6157\,
            I => \N__6136\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6154\,
            I => \N__6129\
        );

    \I__1042\ : Span4Mux_v
    port map (
            O => \N__6151\,
            I => \N__6129\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__6148\,
            I => \N__6129\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6147\,
            I => \N__6126\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6146\,
            I => \N__6123\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6145\,
            I => \N__6120\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6144\,
            I => \N__6117\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6141\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1035\ : Odrv4
    port map (
            O => \N__6136\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1034\ : Odrv4
    port map (
            O => \N__6129\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6126\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6123\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6120\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6117\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1029\ : InMux
    port map (
            O => \N__6102\,
            I => \N__6098\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6101\,
            I => \N__6095\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__6098\,
            I => \N__6089\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__6095\,
            I => \N__6086\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6083\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__6093\,
            I => \N__6077\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6072\
        );

    \I__1022\ : Span4Mux_h
    port map (
            O => \N__6089\,
            I => \N__6069\
        );

    \I__1021\ : Span4Mux_h
    port map (
            O => \N__6086\,
            I => \N__6064\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6083\,
            I => \N__6064\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6061\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6058\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6080\,
            I => \N__6055\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6052\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6047\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6075\,
            I => \N__6047\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__6072\,
            I => \U712_CHIP_RAM.N_545\
        );

    \I__1012\ : Odrv4
    port map (
            O => \N__6069\,
            I => \U712_CHIP_RAM.N_545\
        );

    \I__1011\ : Odrv4
    port map (
            O => \N__6064\,
            I => \U712_CHIP_RAM.N_545\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__6061\,
            I => \U712_CHIP_RAM.N_545\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6058\,
            I => \U712_CHIP_RAM.N_545\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6055\,
            I => \U712_CHIP_RAM.N_545\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6052\,
            I => \U712_CHIP_RAM.N_545\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6047\,
            I => \U712_CHIP_RAM.N_545\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6030\,
            I => \N__6023\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6029\,
            I => \N__6023\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6019\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6023\,
            I => \N__6016\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6022\,
            I => \N__6013\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__6019\,
            I => \U712_CHIP_RAM.N_572\
        );

    \I__999\ : Odrv12
    port map (
            O => \N__6016\,
            I => \U712_CHIP_RAM.N_572\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__6013\,
            I => \U712_CHIP_RAM.N_572\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__6006\,
            I => \U712_CHIP_RAM.N_518_cascade_\
        );

    \I__996\ : InMux
    port map (
            O => \N__6003\,
            I => \N__5999\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__6002\,
            I => \N__5996\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5999\,
            I => \N__5993\
        );

    \I__993\ : InMux
    port map (
            O => \N__5996\,
            I => \N__5985\
        );

    \I__992\ : Span4Mux_v
    port map (
            O => \N__5993\,
            I => \N__5982\
        );

    \I__991\ : InMux
    port map (
            O => \N__5992\,
            I => \N__5979\
        );

    \I__990\ : InMux
    port map (
            O => \N__5991\,
            I => \N__5974\
        );

    \I__989\ : InMux
    port map (
            O => \N__5990\,
            I => \N__5974\
        );

    \I__988\ : InMux
    port map (
            O => \N__5989\,
            I => \N__5969\
        );

    \I__987\ : InMux
    port map (
            O => \N__5988\,
            I => \N__5969\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5985\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__985\ : Odrv4
    port map (
            O => \N__5982\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5979\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5974\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5969\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__981\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5955\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__5955\,
            I => \N__5952\
        );

    \I__979\ : Odrv4
    port map (
            O => \N__5952\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0\
        );

    \I__978\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5946\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5946\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\
        );

    \I__976\ : InMux
    port map (
            O => \N__5943\,
            I => \N__5940\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__5940\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__5937\,
            I => \U712_CHIP_RAM.N_379_cascade_\
        );

    \I__973\ : InMux
    port map (
            O => \N__5934\,
            I => \N__5931\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5931\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__971\ : InMux
    port map (
            O => \N__5928\,
            I => \N__5925\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5925\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__969\ : SRMux
    port map (
            O => \N__5922\,
            I => \N__5919\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5919\,
            I => \N__5916\
        );

    \I__967\ : Odrv12
    port map (
            O => \N__5916\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__5913\,
            I => \U712_CHIP_RAM.REFRESH_RST_cascade_\
        );

    \I__965\ : InMux
    port map (
            O => \N__5910\,
            I => \N__5907\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5907\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i\
        );

    \I__963\ : IoInMux
    port map (
            O => \N__5904\,
            I => \N__5901\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5901\,
            I => \N__5898\
        );

    \I__961\ : IoSpan4Mux
    port map (
            O => \N__5898\,
            I => \N__5895\
        );

    \I__960\ : Span4Mux_s2_v
    port map (
            O => \N__5895\,
            I => \N__5892\
        );

    \I__959\ : Sp12to4
    port map (
            O => \N__5892\,
            I => \N__5888\
        );

    \I__958\ : InMux
    port map (
            O => \N__5891\,
            I => \N__5885\
        );

    \I__957\ : Span12Mux_s8_v
    port map (
            O => \N__5888\,
            I => \N__5882\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__5885\,
            I => \N__5879\
        );

    \I__955\ : Span12Mux_v
    port map (
            O => \N__5882\,
            I => \N__5876\
        );

    \I__954\ : Span4Mux_v
    port map (
            O => \N__5879\,
            I => \N__5873\
        );

    \I__953\ : Span12Mux_h
    port map (
            O => \N__5876\,
            I => \N__5868\
        );

    \I__952\ : Sp12to4
    port map (
            O => \N__5873\,
            I => \N__5868\
        );

    \I__951\ : Span12Mux_h
    port map (
            O => \N__5868\,
            I => \N__5865\
        );

    \I__950\ : Odrv12
    port map (
            O => \N__5865\,
            I => \A_c_11\
        );

    \I__949\ : InMux
    port map (
            O => \N__5862\,
            I => \N__5859\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5859\,
            I => \N__5856\
        );

    \I__947\ : Span4Mux_v
    port map (
            O => \N__5856\,
            I => \N__5853\
        );

    \I__946\ : Span4Mux_v
    port map (
            O => \N__5853\,
            I => \N__5850\
        );

    \I__945\ : Sp12to4
    port map (
            O => \N__5850\,
            I => \N__5847\
        );

    \I__944\ : Span12Mux_h
    port map (
            O => \N__5847\,
            I => \N__5844\
        );

    \I__943\ : Odrv12
    port map (
            O => \N__5844\,
            I => \A_c_4\
        );

    \I__942\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5838\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5838\,
            I => \U712_CHIP_RAM.N_517\
        );

    \I__940\ : InMux
    port map (
            O => \N__5835\,
            I => \N__5830\
        );

    \I__939\ : InMux
    port map (
            O => \N__5834\,
            I => \N__5825\
        );

    \I__938\ : InMux
    port map (
            O => \N__5833\,
            I => \N__5825\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__5830\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5825\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__935\ : IoInMux
    port map (
            O => \N__5820\,
            I => \N__5817\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5817\,
            I => \N__5813\
        );

    \I__933\ : IoInMux
    port map (
            O => \N__5816\,
            I => \N__5810\
        );

    \I__932\ : Span4Mux_s0_v
    port map (
            O => \N__5813\,
            I => \N__5807\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5810\,
            I => \N__5804\
        );

    \I__930\ : Sp12to4
    port map (
            O => \N__5807\,
            I => \N__5801\
        );

    \I__929\ : IoSpan4Mux
    port map (
            O => \N__5804\,
            I => \N__5798\
        );

    \I__928\ : Span12Mux_s11_h
    port map (
            O => \N__5801\,
            I => \N__5795\
        );

    \I__927\ : Sp12to4
    port map (
            O => \N__5798\,
            I => \N__5792\
        );

    \I__926\ : Span12Mux_v
    port map (
            O => \N__5795\,
            I => \N__5786\
        );

    \I__925\ : Span12Mux_v
    port map (
            O => \N__5792\,
            I => \N__5786\
        );

    \I__924\ : InMux
    port map (
            O => \N__5791\,
            I => \N__5783\
        );

    \I__923\ : Odrv12
    port map (
            O => \N__5786\,
            I => \ASn_c\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__5783\,
            I => \ASn_c\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__5778\,
            I => \N__5774\
        );

    \I__920\ : InMux
    port map (
            O => \N__5777\,
            I => \N__5769\
        );

    \I__919\ : InMux
    port map (
            O => \N__5774\,
            I => \N__5766\
        );

    \I__918\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5763\
        );

    \I__917\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5760\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5769\,
            I => \N__5757\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__5766\,
            I => \REG_TACK\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__5763\,
            I => \REG_TACK\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5760\,
            I => \REG_TACK\
        );

    \I__912\ : Odrv4
    port map (
            O => \N__5757\,
            I => \REG_TACK\
        );

    \I__911\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5744\
        );

    \I__910\ : InMux
    port map (
            O => \N__5747\,
            I => \N__5741\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5744\,
            I => \N__5738\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__5741\,
            I => \N__5735\
        );

    \I__907\ : Span4Mux_v
    port map (
            O => \N__5738\,
            I => \N__5732\
        );

    \I__906\ : Span4Mux_v
    port map (
            O => \N__5735\,
            I => \N__5729\
        );

    \I__905\ : Sp12to4
    port map (
            O => \N__5732\,
            I => \N__5726\
        );

    \I__904\ : Span4Mux_h
    port map (
            O => \N__5729\,
            I => \N__5723\
        );

    \I__903\ : Span12Mux_h
    port map (
            O => \N__5726\,
            I => \N__5718\
        );

    \I__902\ : Sp12to4
    port map (
            O => \N__5723\,
            I => \N__5718\
        );

    \I__901\ : Odrv12
    port map (
            O => \N__5718\,
            I => \AWEn_c\
        );

    \I__900\ : InMux
    port map (
            O => \N__5715\,
            I => \N__5711\
        );

    \I__899\ : InMux
    port map (
            O => \N__5714\,
            I => \N__5708\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__5711\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5708\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__896\ : IoInMux
    port map (
            O => \N__5703\,
            I => \N__5700\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__5700\,
            I => \N__5697\
        );

    \I__894\ : IoSpan4Mux
    port map (
            O => \N__5697\,
            I => \N__5694\
        );

    \I__893\ : Span4Mux_s3_v
    port map (
            O => \N__5694\,
            I => \N__5691\
        );

    \I__892\ : Span4Mux_v
    port map (
            O => \N__5691\,
            I => \N__5688\
        );

    \I__891\ : Sp12to4
    port map (
            O => \N__5688\,
            I => \N__5685\
        );

    \I__890\ : Span12Mux_v
    port map (
            O => \N__5685\,
            I => \N__5681\
        );

    \I__889\ : InMux
    port map (
            O => \N__5684\,
            I => \N__5678\
        );

    \I__888\ : Odrv12
    port map (
            O => \N__5681\,
            I => \DBDIR_c\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5678\,
            I => \DBDIR_c\
        );

    \I__886\ : InMux
    port map (
            O => \N__5673\,
            I => \N__5670\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5670\,
            I => \N__5667\
        );

    \I__884\ : Span4Mux_v
    port map (
            O => \N__5667\,
            I => \N__5664\
        );

    \I__883\ : Odrv4
    port map (
            O => \N__5664\,
            I => \U712_REG_SM.N_447\
        );

    \I__882\ : CascadeMux
    port map (
            O => \N__5661\,
            I => \U712_REG_SM.N_447_cascade_\
        );

    \I__881\ : InMux
    port map (
            O => \N__5658\,
            I => \N__5655\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5655\,
            I => \U712_REG_SM.REG_TACK_RNOZ0Z_0\
        );

    \I__879\ : InMux
    port map (
            O => \N__5652\,
            I => \N__5649\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__5649\,
            I => \U712_REG_SM.N_478\
        );

    \I__877\ : IoInMux
    port map (
            O => \N__5646\,
            I => \N__5643\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5643\,
            I => \N__5640\
        );

    \I__875\ : IoSpan4Mux
    port map (
            O => \N__5640\,
            I => \N__5637\
        );

    \I__874\ : Span4Mux_s2_h
    port map (
            O => \N__5637\,
            I => \N__5634\
        );

    \I__873\ : Sp12to4
    port map (
            O => \N__5634\,
            I => \N__5631\
        );

    \I__872\ : Span12Mux_s11_h
    port map (
            O => \N__5631\,
            I => \N__5628\
        );

    \I__871\ : Span12Mux_v
    port map (
            O => \N__5628\,
            I => \N__5625\
        );

    \I__870\ : Odrv12
    port map (
            O => \N__5625\,
            I => \CMA_c_5\
        );

    \I__869\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5619\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5619\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__867\ : IoInMux
    port map (
            O => \N__5616\,
            I => \N__5613\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5613\,
            I => \N__5610\
        );

    \I__865\ : Span4Mux_s3_h
    port map (
            O => \N__5610\,
            I => \N__5607\
        );

    \I__864\ : Sp12to4
    port map (
            O => \N__5607\,
            I => \N__5604\
        );

    \I__863\ : Span12Mux_v
    port map (
            O => \N__5604\,
            I => \N__5601\
        );

    \I__862\ : Span12Mux_h
    port map (
            O => \N__5601\,
            I => \N__5598\
        );

    \I__861\ : Odrv12
    port map (
            O => \N__5598\,
            I => \CMA_c_7\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__5595\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\
        );

    \I__859\ : CEMux
    port map (
            O => \N__5592\,
            I => \N__5589\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5589\,
            I => \N__5586\
        );

    \I__857\ : Span4Mux_h
    port map (
            O => \N__5586\,
            I => \N__5583\
        );

    \I__856\ : Odrv4
    port map (
            O => \N__5583\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_1\
        );

    \I__855\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5576\
        );

    \I__854\ : InMux
    port map (
            O => \N__5579\,
            I => \N__5573\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5576\,
            I => \U712_CHIP_RAM.N_666\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5573\,
            I => \U712_CHIP_RAM.N_666\
        );

    \I__851\ : InMux
    port map (
            O => \N__5568\,
            I => \N__5565\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5565\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__5562\,
            I => \N__5559\
        );

    \I__848\ : InMux
    port map (
            O => \N__5559\,
            I => \N__5552\
        );

    \I__847\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5549\
        );

    \I__846\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5545\
        );

    \I__845\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5540\
        );

    \I__844\ : InMux
    port map (
            O => \N__5555\,
            I => \N__5540\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__5552\,
            I => \N__5535\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5549\,
            I => \N__5535\
        );

    \I__841\ : InMux
    port map (
            O => \N__5548\,
            I => \N__5532\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5545\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5540\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__5535\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5532\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__836\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5519\
        );

    \I__835\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5513\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5519\,
            I => \N__5510\
        );

    \I__833\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5507\
        );

    \I__832\ : InMux
    port map (
            O => \N__5517\,
            I => \N__5504\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__5516\,
            I => \N__5500\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5513\,
            I => \N__5497\
        );

    \I__829\ : Span4Mux_v
    port map (
            O => \N__5510\,
            I => \N__5494\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5507\,
            I => \N__5489\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5504\,
            I => \N__5489\
        );

    \I__826\ : InMux
    port map (
            O => \N__5503\,
            I => \N__5486\
        );

    \I__825\ : InMux
    port map (
            O => \N__5500\,
            I => \N__5483\
        );

    \I__824\ : Span4Mux_v
    port map (
            O => \N__5497\,
            I => \N__5480\
        );

    \I__823\ : Odrv4
    port map (
            O => \N__5494\,
            I => \U712_CHIP_RAM.N_557\
        );

    \I__822\ : Odrv4
    port map (
            O => \N__5489\,
            I => \U712_CHIP_RAM.N_557\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5486\,
            I => \U712_CHIP_RAM.N_557\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5483\,
            I => \U712_CHIP_RAM.N_557\
        );

    \I__819\ : Odrv4
    port map (
            O => \N__5480\,
            I => \U712_CHIP_RAM.N_557\
        );

    \I__818\ : InMux
    port map (
            O => \N__5469\,
            I => \N__5466\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5466\,
            I => \U712_CHIP_RAM.N_393\
        );

    \I__816\ : InMux
    port map (
            O => \N__5463\,
            I => \N__5459\
        );

    \I__815\ : InMux
    port map (
            O => \N__5462\,
            I => \N__5456\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__5459\,
            I => \N__5453\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5456\,
            I => \N__5450\
        );

    \I__812\ : Span4Mux_h
    port map (
            O => \N__5453\,
            I => \N__5445\
        );

    \I__811\ : Span4Mux_h
    port map (
            O => \N__5450\,
            I => \N__5445\
        );

    \I__810\ : Odrv4
    port map (
            O => \N__5445\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_0_a2_0\
        );

    \I__809\ : CascadeMux
    port map (
            O => \N__5442\,
            I => \U712_CHIP_RAM.N_557_cascade_\
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__5439\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\
        );

    \I__807\ : InMux
    port map (
            O => \N__5436\,
            I => \N__5433\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5433\,
            I => \N__5430\
        );

    \I__805\ : Odrv4
    port map (
            O => \N__5430\,
            I => \U712_CHIP_RAM.N_31\
        );

    \I__804\ : IoInMux
    port map (
            O => \N__5427\,
            I => \N__5424\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5424\,
            I => \N__5421\
        );

    \I__802\ : Span4Mux_s1_v
    port map (
            O => \N__5421\,
            I => \N__5418\
        );

    \I__801\ : Sp12to4
    port map (
            O => \N__5418\,
            I => \N__5415\
        );

    \I__800\ : Span12Mux_h
    port map (
            O => \N__5415\,
            I => \N__5412\
        );

    \I__799\ : Span12Mux_v
    port map (
            O => \N__5412\,
            I => \N__5408\
        );

    \I__798\ : InMux
    port map (
            O => \N__5411\,
            I => \N__5405\
        );

    \I__797\ : Odrv12
    port map (
            O => \N__5408\,
            I => \LATCH_CLK_c\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5405\,
            I => \LATCH_CLK_c\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__5400\,
            I => \N__5397\
        );

    \I__794\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5390\
        );

    \I__793\ : InMux
    port map (
            O => \N__5396\,
            I => \N__5387\
        );

    \I__792\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5381\
        );

    \I__791\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5381\
        );

    \I__790\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5373\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5390\,
            I => \N__5368\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5387\,
            I => \N__5368\
        );

    \I__787\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5365\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5381\,
            I => \N__5362\
        );

    \I__785\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5359\
        );

    \I__784\ : InMux
    port map (
            O => \N__5379\,
            I => \N__5354\
        );

    \I__783\ : InMux
    port map (
            O => \N__5378\,
            I => \N__5354\
        );

    \I__782\ : InMux
    port map (
            O => \N__5377\,
            I => \N__5349\
        );

    \I__781\ : InMux
    port map (
            O => \N__5376\,
            I => \N__5349\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5373\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__779\ : Odrv4
    port map (
            O => \N__5368\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5365\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__777\ : Odrv4
    port map (
            O => \N__5362\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__5359\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5354\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5349\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__773\ : InMux
    port map (
            O => \N__5334\,
            I => \N__5331\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5331\,
            I => \N__5327\
        );

    \I__771\ : InMux
    port map (
            O => \N__5330\,
            I => \N__5324\
        );

    \I__770\ : Odrv12
    port map (
            O => \N__5327\,
            I => \U712_CHIP_RAM.N_566\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5324\,
            I => \U712_CHIP_RAM.N_566\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__5319\,
            I => \N__5314\
        );

    \I__767\ : CascadeMux
    port map (
            O => \N__5318\,
            I => \N__5311\
        );

    \I__766\ : InMux
    port map (
            O => \N__5317\,
            I => \N__5307\
        );

    \I__765\ : InMux
    port map (
            O => \N__5314\,
            I => \N__5302\
        );

    \I__764\ : InMux
    port map (
            O => \N__5311\,
            I => \N__5302\
        );

    \I__763\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5299\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__5307\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__5302\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__5299\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__759\ : IoInMux
    port map (
            O => \N__5292\,
            I => \N__5288\
        );

    \I__758\ : IoInMux
    port map (
            O => \N__5291\,
            I => \N__5285\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__5288\,
            I => \N__5282\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__5285\,
            I => \N__5279\
        );

    \I__755\ : IoSpan4Mux
    port map (
            O => \N__5282\,
            I => \N__5276\
        );

    \I__754\ : IoSpan4Mux
    port map (
            O => \N__5279\,
            I => \N__5273\
        );

    \I__753\ : Sp12to4
    port map (
            O => \N__5276\,
            I => \N__5269\
        );

    \I__752\ : Span4Mux_s2_h
    port map (
            O => \N__5273\,
            I => \N__5266\
        );

    \I__751\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5263\
        );

    \I__750\ : Span12Mux_s7_v
    port map (
            O => \N__5269\,
            I => \N__5260\
        );

    \I__749\ : Sp12to4
    port map (
            O => \N__5266\,
            I => \N__5257\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5263\,
            I => \N__5254\
        );

    \I__747\ : Span12Mux_v
    port map (
            O => \N__5260\,
            I => \N__5250\
        );

    \I__746\ : Span12Mux_h
    port map (
            O => \N__5257\,
            I => \N__5247\
        );

    \I__745\ : Span4Mux_h
    port map (
            O => \N__5254\,
            I => \N__5244\
        );

    \I__744\ : InMux
    port map (
            O => \N__5253\,
            I => \N__5241\
        );

    \I__743\ : Odrv12
    port map (
            O => \N__5250\,
            I => \TACK_OUTn\
        );

    \I__742\ : Odrv12
    port map (
            O => \N__5247\,
            I => \TACK_OUTn\
        );

    \I__741\ : Odrv4
    port map (
            O => \N__5244\,
            I => \TACK_OUTn\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5241\,
            I => \TACK_OUTn\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__5232\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\
        );

    \I__738\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5226\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__5226\,
            I => \N__5223\
        );

    \I__736\ : Span12Mux_v
    port map (
            O => \N__5223\,
            I => \N__5220\
        );

    \I__735\ : Span12Mux_h
    port map (
            O => \N__5220\,
            I => \N__5217\
        );

    \I__734\ : Odrv12
    port map (
            O => \N__5217\,
            I => \A_c_20\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__5214\,
            I => \U712_CHIP_RAM.N_506_cascade_\
        );

    \I__732\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5207\
        );

    \I__731\ : InMux
    port map (
            O => \N__5210\,
            I => \N__5204\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__5207\,
            I => \N__5201\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__5204\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__728\ : Odrv12
    port map (
            O => \N__5201\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__727\ : InMux
    port map (
            O => \N__5196\,
            I => \N__5193\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5193\,
            I => \N__5190\
        );

    \I__725\ : Span4Mux_v
    port map (
            O => \N__5190\,
            I => \N__5187\
        );

    \I__724\ : Odrv4
    port map (
            O => \N__5187\,
            I => \U712_CHIP_RAM.N_375\
        );

    \I__723\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5177\
        );

    \I__722\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5172\
        );

    \I__721\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5172\
        );

    \I__720\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5169\
        );

    \I__719\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5166\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5177\,
            I => \U712_CHIP_RAM.N_547\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5172\,
            I => \U712_CHIP_RAM.N_547\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5169\,
            I => \U712_CHIP_RAM.N_547\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5166\,
            I => \U712_CHIP_RAM.N_547\
        );

    \I__714\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5154\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__5154\,
            I => \N__5149\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__5153\,
            I => \N__5146\
        );

    \I__711\ : InMux
    port map (
            O => \N__5152\,
            I => \N__5142\
        );

    \I__710\ : Span4Mux_h
    port map (
            O => \N__5149\,
            I => \N__5139\
        );

    \I__709\ : InMux
    port map (
            O => \N__5146\,
            I => \N__5136\
        );

    \I__708\ : InMux
    port map (
            O => \N__5145\,
            I => \N__5133\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__5142\,
            I => \N__5130\
        );

    \I__706\ : Odrv4
    port map (
            O => \N__5139\,
            I => \U712_CHIP_RAM.N_522\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5136\,
            I => \U712_CHIP_RAM.N_522\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5133\,
            I => \U712_CHIP_RAM.N_522\
        );

    \I__703\ : Odrv4
    port map (
            O => \N__5130\,
            I => \U712_CHIP_RAM.N_522\
        );

    \I__702\ : CascadeMux
    port map (
            O => \N__5121\,
            I => \U712_CHIP_RAM.N_523_cascade_\
        );

    \I__701\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5115\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__5115\,
            I => \U712_CHIP_RAM.BANK0_9\
        );

    \I__699\ : IoInMux
    port map (
            O => \N__5112\,
            I => \N__5109\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5109\,
            I => \N__5106\
        );

    \I__697\ : Span12Mux_s5_v
    port map (
            O => \N__5106\,
            I => \N__5103\
        );

    \I__696\ : Span12Mux_v
    port map (
            O => \N__5103\,
            I => \N__5099\
        );

    \I__695\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5096\
        );

    \I__694\ : Odrv12
    port map (
            O => \N__5099\,
            I => \BANK0_c\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__5096\,
            I => \BANK0_c\
        );

    \I__692\ : InMux
    port map (
            O => \N__5091\,
            I => \N__5087\
        );

    \I__691\ : InMux
    port map (
            O => \N__5090\,
            I => \N__5084\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__5087\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5084\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__688\ : InMux
    port map (
            O => \N__5079\,
            I => \N__5075\
        );

    \I__687\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5072\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5075\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__5072\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__684\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5063\
        );

    \I__683\ : InMux
    port map (
            O => \N__5066\,
            I => \N__5060\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5063\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5060\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__680\ : CascadeMux
    port map (
            O => \N__5055\,
            I => \U712_CHIP_RAM.N_545_cascade_\
        );

    \I__679\ : InMux
    port map (
            O => \N__5052\,
            I => \N__5046\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__5051\,
            I => \N__5043\
        );

    \I__677\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5036\
        );

    \I__676\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5036\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5046\,
            I => \N__5033\
        );

    \I__674\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5026\
        );

    \I__673\ : InMux
    port map (
            O => \N__5042\,
            I => \N__5026\
        );

    \I__672\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5026\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__5036\,
            I => \U712_CHIP_RAM.N_549\
        );

    \I__670\ : Odrv4
    port map (
            O => \N__5033\,
            I => \U712_CHIP_RAM.N_549\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5026\,
            I => \U712_CHIP_RAM.N_549\
        );

    \I__668\ : InMux
    port map (
            O => \N__5019\,
            I => \N__5010\
        );

    \I__667\ : InMux
    port map (
            O => \N__5018\,
            I => \N__5010\
        );

    \I__666\ : InMux
    port map (
            O => \N__5017\,
            I => \N__5010\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5010\,
            I => \N__5006\
        );

    \I__664\ : InMux
    port map (
            O => \N__5009\,
            I => \N__5002\
        );

    \I__663\ : Span4Mux_h
    port map (
            O => \N__5006\,
            I => \N__4999\
        );

    \I__662\ : InMux
    port map (
            O => \N__5005\,
            I => \N__4996\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5002\,
            I => \U712_CHIP_RAM.N_560\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__4999\,
            I => \U712_CHIP_RAM.N_560\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__4996\,
            I => \U712_CHIP_RAM.N_560\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__4989\,
            I => \N__4986\
        );

    \I__657\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4983\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__4983\,
            I => \U712_CHIP_RAM.N_501\
        );

    \I__655\ : InMux
    port map (
            O => \N__4980\,
            I => \N__4977\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4977\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1\
        );

    \I__653\ : InMux
    port map (
            O => \N__4974\,
            I => \N__4968\
        );

    \I__652\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4968\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__4968\,
            I => \U712_CHIP_RAM.N_515\
        );

    \I__650\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4962\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__4962\,
            I => \U712_CHIP_RAM.N_516\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__4959\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\
        );

    \I__647\ : InMux
    port map (
            O => \N__4956\,
            I => \N__4952\
        );

    \I__646\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4949\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4952\,
            I => \U712_CHIP_RAM.N_519\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4949\,
            I => \U712_CHIP_RAM.N_519\
        );

    \I__643\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4941\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__4941\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0\
        );

    \I__641\ : IoInMux
    port map (
            O => \N__4938\,
            I => \N__4935\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4935\,
            I => \N__4932\
        );

    \I__639\ : Span4Mux_s2_v
    port map (
            O => \N__4932\,
            I => \N__4929\
        );

    \I__638\ : Sp12to4
    port map (
            O => \N__4929\,
            I => \N__4925\
        );

    \I__637\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4922\
        );

    \I__636\ : Span12Mux_h
    port map (
            O => \N__4925\,
            I => \N__4919\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4922\,
            I => \N__4916\
        );

    \I__634\ : Odrv12
    port map (
            O => \N__4919\,
            I => \CONSTANT_ONE_NET\
        );

    \I__633\ : Odrv12
    port map (
            O => \N__4916\,
            I => \CONSTANT_ONE_NET\
        );

    \I__632\ : InMux
    port map (
            O => \N__4911\,
            I => \N__4908\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4908\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_0\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__4905\,
            I => \N__4899\
        );

    \I__629\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4890\
        );

    \I__628\ : InMux
    port map (
            O => \N__4903\,
            I => \N__4890\
        );

    \I__627\ : InMux
    port map (
            O => \N__4902\,
            I => \N__4887\
        );

    \I__626\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4884\
        );

    \I__625\ : InMux
    port map (
            O => \N__4898\,
            I => \N__4875\
        );

    \I__624\ : InMux
    port map (
            O => \N__4897\,
            I => \N__4875\
        );

    \I__623\ : InMux
    port map (
            O => \N__4896\,
            I => \N__4875\
        );

    \I__622\ : InMux
    port map (
            O => \N__4895\,
            I => \N__4875\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__4890\,
            I => \N__4872\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__4887\,
            I => \U712_CHIP_RAM.N_78\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4884\,
            I => \U712_CHIP_RAM.N_78\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__4875\,
            I => \U712_CHIP_RAM.N_78\
        );

    \I__617\ : Odrv4
    port map (
            O => \N__4872\,
            I => \U712_CHIP_RAM.N_78\
        );

    \I__616\ : CEMux
    port map (
            O => \N__4863\,
            I => \N__4858\
        );

    \I__615\ : CEMux
    port map (
            O => \N__4862\,
            I => \N__4855\
        );

    \I__614\ : CEMux
    port map (
            O => \N__4861\,
            I => \N__4852\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__4858\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4855\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__4852\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__610\ : CascadeMux
    port map (
            O => \N__4845\,
            I => \U712_CHIP_RAM.N_559_cascade_\
        );

    \I__609\ : InMux
    port map (
            O => \N__4842\,
            I => \N__4836\
        );

    \I__608\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4836\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__4836\,
            I => \U712_CHIP_RAM.N_665\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__4833\,
            I => \U712_CHIP_RAM.N_665_cascade_\
        );

    \I__605\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4827\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4827\,
            I => \U712_CHIP_RAM.N_471\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__4824\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\
        );

    \I__602\ : InMux
    port map (
            O => \N__4821\,
            I => \N__4817\
        );

    \I__601\ : InMux
    port map (
            O => \N__4820\,
            I => \N__4814\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__4817\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4814\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__598\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4805\
        );

    \I__597\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4802\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__4805\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4802\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__594\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4793\
        );

    \I__593\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4790\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4793\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4790\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__590\ : InMux
    port map (
            O => \N__4785\,
            I => \N__4782\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4782\,
            I => \N__4779\
        );

    \I__588\ : Span12Mux_v
    port map (
            O => \N__4779\,
            I => \N__4776\
        );

    \I__587\ : Span12Mux_h
    port map (
            O => \N__4776\,
            I => \N__4773\
        );

    \I__586\ : Odrv12
    port map (
            O => \N__4773\,
            I => \A_c_14\
        );

    \I__585\ : InMux
    port map (
            O => \N__4770\,
            I => \N__4767\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4767\,
            I => \N__4764\
        );

    \I__583\ : Span4Mux_v
    port map (
            O => \N__4764\,
            I => \N__4761\
        );

    \I__582\ : Sp12to4
    port map (
            O => \N__4761\,
            I => \N__4758\
        );

    \I__581\ : Span12Mux_h
    port map (
            O => \N__4758\,
            I => \N__4755\
        );

    \I__580\ : Odrv12
    port map (
            O => \N__4755\,
            I => \A_c_7\
        );

    \I__579\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4748\
        );

    \I__578\ : InMux
    port map (
            O => \N__4751\,
            I => \N__4745\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__4748\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__4745\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__575\ : InMux
    port map (
            O => \N__4740\,
            I => \N__4736\
        );

    \I__574\ : InMux
    port map (
            O => \N__4739\,
            I => \N__4733\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4736\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4733\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__4728\,
            I => \N__4724\
        );

    \I__570\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4721\
        );

    \I__569\ : InMux
    port map (
            O => \N__4724\,
            I => \N__4718\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4721\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4718\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__566\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4709\
        );

    \I__565\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4706\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4709\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4706\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__562\ : InMux
    port map (
            O => \N__4701\,
            I => \N__4698\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__4698\,
            I => \N__4695\
        );

    \I__560\ : Span4Mux_v
    port map (
            O => \N__4695\,
            I => \N__4692\
        );

    \I__559\ : Sp12to4
    port map (
            O => \N__4692\,
            I => \N__4689\
        );

    \I__558\ : Span12Mux_h
    port map (
            O => \N__4689\,
            I => \N__4686\
        );

    \I__557\ : Odrv12
    port map (
            O => \N__4686\,
            I => \A_c_8\
        );

    \I__556\ : InMux
    port map (
            O => \N__4683\,
            I => \N__4680\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4680\,
            I => \N__4677\
        );

    \I__554\ : Span4Mux_v
    port map (
            O => \N__4677\,
            I => \N__4674\
        );

    \I__553\ : Sp12to4
    port map (
            O => \N__4674\,
            I => \N__4671\
        );

    \I__552\ : Span12Mux_h
    port map (
            O => \N__4671\,
            I => \N__4668\
        );

    \I__551\ : Span12Mux_v
    port map (
            O => \N__4668\,
            I => \N__4665\
        );

    \I__550\ : Odrv12
    port map (
            O => \N__4665\,
            I => \A_c_15\
        );

    \I__549\ : CascadeMux
    port map (
            O => \N__4662\,
            I => \U712_CHIP_RAM.N_669_cascade_\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__4659\,
            I => \U712_CHIP_RAM.N_520_cascade_\
        );

    \I__547\ : CascadeMux
    port map (
            O => \N__4656\,
            I => \U712_CYCLE_TERM.N_539_cascade_\
        );

    \I__546\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4647\
        );

    \I__545\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4644\
        );

    \I__544\ : InMux
    port map (
            O => \N__4651\,
            I => \N__4639\
        );

    \I__543\ : InMux
    port map (
            O => \N__4650\,
            I => \N__4639\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4647\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__4644\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4639\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__539\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4624\
        );

    \I__538\ : InMux
    port map (
            O => \N__4631\,
            I => \N__4624\
        );

    \I__537\ : InMux
    port map (
            O => \N__4630\,
            I => \N__4621\
        );

    \I__536\ : InMux
    port map (
            O => \N__4629\,
            I => \N__4618\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4624\,
            I => \CPU_TACKm\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__4621\,
            I => \CPU_TACKm\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__4618\,
            I => \CPU_TACKm\
        );

    \I__532\ : InMux
    port map (
            O => \N__4611\,
            I => \N__4608\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__4608\,
            I => \N__4603\
        );

    \I__530\ : InMux
    port map (
            O => \N__4607\,
            I => \N__4600\
        );

    \I__529\ : InMux
    port map (
            O => \N__4606\,
            I => \N__4597\
        );

    \I__528\ : Span4Mux_h
    port map (
            O => \N__4603\,
            I => \N__4594\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4600\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4597\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__525\ : Odrv4
    port map (
            O => \N__4594\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__524\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4584\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4584\,
            I => \N__4581\
        );

    \I__522\ : Span4Mux_v
    port map (
            O => \N__4581\,
            I => \N__4578\
        );

    \I__521\ : Span4Mux_v
    port map (
            O => \N__4578\,
            I => \N__4575\
        );

    \I__520\ : Span4Mux_h
    port map (
            O => \N__4575\,
            I => \N__4572\
        );

    \I__519\ : Sp12to4
    port map (
            O => \N__4572\,
            I => \N__4569\
        );

    \I__518\ : Odrv12
    port map (
            O => \N__4569\,
            I => \A_c_6\
        );

    \I__517\ : InMux
    port map (
            O => \N__4566\,
            I => \N__4563\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4563\,
            I => \N__4560\
        );

    \I__515\ : Span4Mux_v
    port map (
            O => \N__4560\,
            I => \N__4557\
        );

    \I__514\ : Sp12to4
    port map (
            O => \N__4557\,
            I => \N__4554\
        );

    \I__513\ : Span12Mux_h
    port map (
            O => \N__4554\,
            I => \N__4551\
        );

    \I__512\ : Odrv12
    port map (
            O => \N__4551\,
            I => \A_c_13\
        );

    \I__511\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4545\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__4545\,
            I => \N__4542\
        );

    \I__509\ : Span12Mux_v
    port map (
            O => \N__4542\,
            I => \N__4539\
        );

    \I__508\ : Span12Mux_h
    port map (
            O => \N__4539\,
            I => \N__4536\
        );

    \I__507\ : Odrv12
    port map (
            O => \N__4536\,
            I => \A_c_18\
        );

    \I__506\ : InMux
    port map (
            O => \N__4533\,
            I => \N__4530\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4530\,
            I => \N__4527\
        );

    \I__504\ : Span12Mux_v
    port map (
            O => \N__4527\,
            I => \N__4524\
        );

    \I__503\ : Span12Mux_h
    port map (
            O => \N__4524\,
            I => \N__4521\
        );

    \I__502\ : Odrv12
    port map (
            O => \N__4521\,
            I => \A_c_16\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__4518\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\
        );

    \I__500\ : InMux
    port map (
            O => \N__4515\,
            I => \N__4512\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4512\,
            I => \N__4509\
        );

    \I__498\ : Span4Mux_h
    port map (
            O => \N__4509\,
            I => \N__4506\
        );

    \I__497\ : Sp12to4
    port map (
            O => \N__4506\,
            I => \N__4503\
        );

    \I__496\ : Span12Mux_v
    port map (
            O => \N__4503\,
            I => \N__4500\
        );

    \I__495\ : Odrv12
    port map (
            O => \N__4500\,
            I => \A_c_5\
        );

    \I__494\ : InMux
    port map (
            O => \N__4497\,
            I => \N__4494\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__4494\,
            I => \N__4491\
        );

    \I__492\ : Span12Mux_v
    port map (
            O => \N__4491\,
            I => \N__4488\
        );

    \I__491\ : Span12Mux_h
    port map (
            O => \N__4488\,
            I => \N__4485\
        );

    \I__490\ : Odrv12
    port map (
            O => \N__4485\,
            I => \A_c_12\
        );

    \I__489\ : InMux
    port map (
            O => \N__4482\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__488\ : CascadeMux
    port map (
            O => \N__4479\,
            I => \U712_CHIP_RAM.N_666_cascade_\
        );

    \I__487\ : CascadeMux
    port map (
            O => \N__4476\,
            I => \U712_CHIP_RAM.N_393_cascade_\
        );

    \I__486\ : CascadeMux
    port map (
            O => \N__4473\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_\
        );

    \I__485\ : CEMux
    port map (
            O => \N__4470\,
            I => \N__4467\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4467\,
            I => \N__4464\
        );

    \I__483\ : Span4Mux_h
    port map (
            O => \N__4464\,
            I => \N__4461\
        );

    \I__482\ : Span4Mux_h
    port map (
            O => \N__4461\,
            I => \N__4458\
        );

    \I__481\ : Odrv4
    port map (
            O => \N__4458\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\
        );

    \I__480\ : InMux
    port map (
            O => \N__4455\,
            I => \N__4452\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4452\,
            I => \N__4449\
        );

    \I__478\ : Odrv4
    port map (
            O => \N__4449\,
            I => \U712_CHIP_RAM.CLK_EN_6_0\
        );

    \I__477\ : CascadeMux
    port map (
            O => \N__4446\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0_cascade_\
        );

    \I__476\ : IoInMux
    port map (
            O => \N__4443\,
            I => \N__4440\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__4440\,
            I => \N__4437\
        );

    \I__474\ : IoSpan4Mux
    port map (
            O => \N__4437\,
            I => \N__4434\
        );

    \I__473\ : IoSpan4Mux
    port map (
            O => \N__4434\,
            I => \N__4431\
        );

    \I__472\ : Sp12to4
    port map (
            O => \N__4431\,
            I => \N__4428\
        );

    \I__471\ : Span12Mux_s7_h
    port map (
            O => \N__4428\,
            I => \N__4425\
        );

    \I__470\ : Span12Mux_h
    port map (
            O => \N__4425\,
            I => \N__4421\
        );

    \I__469\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4418\
        );

    \I__468\ : Odrv12
    port map (
            O => \N__4421\,
            I => \CLK_EN_c\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4418\,
            I => \CLK_EN_c\
        );

    \I__466\ : InMux
    port map (
            O => \N__4413\,
            I => \N__4410\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4410\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\
        );

    \I__464\ : InMux
    port map (
            O => \N__4407\,
            I => \N__4404\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4404\,
            I => \U712_CHIP_RAM.N_504\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__4401\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_a2_0_cascade_\
        );

    \I__461\ : InMux
    port map (
            O => \N__4398\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__460\ : InMux
    port map (
            O => \N__4395\,
            I => \N__4392\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__4392\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__458\ : InMux
    port map (
            O => \N__4389\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__457\ : InMux
    port map (
            O => \N__4386\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__456\ : InMux
    port map (
            O => \N__4383\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__455\ : InMux
    port map (
            O => \N__4380\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__454\ : InMux
    port map (
            O => \N__4377\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__4374\,
            I => \U712_CHIP_RAM.N_375_cascade_\
        );

    \I__452\ : CascadeMux
    port map (
            O => \N__4371\,
            I => \N__4367\
        );

    \I__451\ : InMux
    port map (
            O => \N__4370\,
            I => \N__4364\
        );

    \I__450\ : InMux
    port map (
            O => \N__4367\,
            I => \N__4361\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__4364\,
            I => \N__4358\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4361\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__447\ : Odrv4
    port map (
            O => \N__4358\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__4353\,
            I => \N__4350\
        );

    \I__445\ : InMux
    port map (
            O => \N__4350\,
            I => \N__4347\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__4347\,
            I => \U712_CHIP_RAM.N_498\
        );

    \I__443\ : CascadeMux
    port map (
            O => \N__4344\,
            I => \U712_CHIP_RAM.N_547_cascade_\
        );

    \I__442\ : CascadeMux
    port map (
            O => \N__4341\,
            I => \U712_CHIP_RAM.N_501_cascade_\
        );

    \I__441\ : InMux
    port map (
            O => \N__4338\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__440\ : InMux
    port map (
            O => \N__4335\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__439\ : InMux
    port map (
            O => \N__4332\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__438\ : InMux
    port map (
            O => \N__4329\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__437\ : InMux
    port map (
            O => \N__4326\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__436\ : InMux
    port map (
            O => \N__4323\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__435\ : ClkMux
    port map (
            O => \N__4320\,
            I => \N__4296\
        );

    \I__434\ : ClkMux
    port map (
            O => \N__4319\,
            I => \N__4296\
        );

    \I__433\ : ClkMux
    port map (
            O => \N__4318\,
            I => \N__4296\
        );

    \I__432\ : ClkMux
    port map (
            O => \N__4317\,
            I => \N__4296\
        );

    \I__431\ : ClkMux
    port map (
            O => \N__4316\,
            I => \N__4296\
        );

    \I__430\ : ClkMux
    port map (
            O => \N__4315\,
            I => \N__4296\
        );

    \I__429\ : ClkMux
    port map (
            O => \N__4314\,
            I => \N__4296\
        );

    \I__428\ : ClkMux
    port map (
            O => \N__4313\,
            I => \N__4296\
        );

    \I__427\ : GlobalMux
    port map (
            O => \N__4296\,
            I => \N__4293\
        );

    \I__426\ : gio2CtrlBuf
    port map (
            O => \N__4293\,
            I => \C1_c_g\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__4290\,
            I => \U712_CHIP_RAM.N_371_cascade_\
        );

    \I__424\ : CascadeMux
    port map (
            O => \N__4287\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_2_cascade_\
        );

    \I__423\ : InMux
    port map (
            O => \N__4284\,
            I => \N__4281\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4281\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1\
        );

    \I__421\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4274\
        );

    \I__420\ : InMux
    port map (
            O => \N__4277\,
            I => \N__4271\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__4274\,
            I => \N__4268\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__4271\,
            I => \U712_CYCLE_TERM.N_565\
        );

    \I__417\ : Odrv4
    port map (
            O => \N__4268\,
            I => \U712_CYCLE_TERM.N_565\
        );

    \I__416\ : InMux
    port map (
            O => \N__4263\,
            I => \N__4259\
        );

    \I__415\ : InMux
    port map (
            O => \N__4262\,
            I => \N__4256\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__4259\,
            I => \N__4253\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__4256\,
            I => \U712_CYCLE_TERM.N_407\
        );

    \I__412\ : Odrv4
    port map (
            O => \N__4253\,
            I => \U712_CYCLE_TERM.N_407\
        );

    \I__411\ : InMux
    port map (
            O => \N__4248\,
            I => \N__4245\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__4245\,
            I => \N__4242\
        );

    \I__409\ : Odrv4
    port map (
            O => \N__4242\,
            I => \U712_CYCLE_TERM.N_534\
        );

    \I__408\ : InMux
    port map (
            O => \N__4239\,
            I => \bfn_9_9_0_\
        );

    \I__407\ : InMux
    port map (
            O => \N__4236\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__406\ : InMux
    port map (
            O => \N__4233\,
            I => \N__4227\
        );

    \I__405\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4227\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4227\,
            I => \U712_CHIP_RAM.N_373\
        );

    \I__403\ : InMux
    port map (
            O => \N__4224\,
            I => \N__4221\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__4221\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0\
        );

    \I__401\ : InMux
    port map (
            O => \N__4218\,
            I => \N__4215\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__4215\,
            I => \N__4212\
        );

    \I__399\ : Odrv4
    port map (
            O => \N__4212\,
            I => \U712_CHIP_RAM.N_409\
        );

    \I__398\ : CascadeMux
    port map (
            O => \N__4209\,
            I => \U712_REG_SM.N_486_cascade_\
        );

    \I__397\ : InMux
    port map (
            O => \N__4206\,
            I => \N__4203\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__4203\,
            I => \U712_CHIP_RAM.CLK_EN_6_0_a3_0_a2_1\
        );

    \I__395\ : IoInMux
    port map (
            O => \N__4200\,
            I => \N__4197\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__4197\,
            I => \N__4194\
        );

    \I__393\ : Span12Mux_s9_v
    port map (
            O => \N__4194\,
            I => \N__4191\
        );

    \I__392\ : Odrv12
    port map (
            O => \N__4191\,
            I => \N_490\
        );

    \I__391\ : CEMux
    port map (
            O => \N__4188\,
            I => \N__4185\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__4185\,
            I => \N__4182\
        );

    \I__389\ : Span4Mux_v
    port map (
            O => \N__4182\,
            I => \N__4179\
        );

    \I__388\ : Odrv4
    port map (
            O => \N__4179\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0\
        );

    \I__387\ : CascadeMux
    port map (
            O => \N__4176\,
            I => \U712_CHIP_RAM.N_554_cascade_\
        );

    \I__386\ : CascadeMux
    port map (
            O => \N__4173\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_a2_0_cascade_\
        );

    \I__385\ : IoInMux
    port map (
            O => \N__4170\,
            I => \N__4167\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__4167\,
            I => \N__4164\
        );

    \I__383\ : IoSpan4Mux
    port map (
            O => \N__4164\,
            I => \N__4161\
        );

    \I__382\ : Span4Mux_s3_v
    port map (
            O => \N__4161\,
            I => \N__4158\
        );

    \I__381\ : Odrv4
    port map (
            O => \N__4158\,
            I => \CLK80_PLL_i_i\
        );

    \I__380\ : CascadeMux
    port map (
            O => \N__4155\,
            I => \DBRn_c_i_cascade_\
        );

    \I__379\ : IoInMux
    port map (
            O => \N__4152\,
            I => \N__4149\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__4149\,
            I => \N__4146\
        );

    \I__377\ : IoSpan4Mux
    port map (
            O => \N__4146\,
            I => \N__4143\
        );

    \I__376\ : Sp12to4
    port map (
            O => \N__4143\,
            I => \N__4140\
        );

    \I__375\ : Odrv12
    port map (
            O => \N__4140\,
            I => \DBRn_c_i_0\
        );

    \I__374\ : CascadeMux
    port map (
            O => \N__4137\,
            I => \N__4134\
        );

    \I__373\ : InMux
    port map (
            O => \N__4134\,
            I => \N__4131\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__4131\,
            I => \DBRn_c_i\
        );

    \I__371\ : IoInMux
    port map (
            O => \N__4128\,
            I => \N__4125\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__4125\,
            I => \N__4122\
        );

    \I__369\ : IoSpan4Mux
    port map (
            O => \N__4122\,
            I => \N__4119\
        );

    \I__368\ : Span4Mux_s2_v
    port map (
            O => \N__4119\,
            I => \N__4116\
        );

    \I__367\ : Sp12to4
    port map (
            O => \N__4116\,
            I => \N__4113\
        );

    \I__366\ : Span12Mux_v
    port map (
            O => \N__4113\,
            I => \N__4110\
        );

    \I__365\ : Span12Mux_h
    port map (
            O => \N__4110\,
            I => \N__4107\
        );

    \I__364\ : Odrv12
    port map (
            O => \N__4107\,
            I => \U712_CYCLE_TERM_TCIn_0_i\
        );

    \I__363\ : CascadeMux
    port map (
            O => \N__4104\,
            I => \N__4100\
        );

    \I__362\ : InMux
    port map (
            O => \N__4103\,
            I => \N__4097\
        );

    \I__361\ : InMux
    port map (
            O => \N__4100\,
            I => \N__4094\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__4097\,
            I => \U712_CYCLE_TERM.RAM_CYCLEZ0\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__4094\,
            I => \U712_CYCLE_TERM.RAM_CYCLEZ0\
        );

    \I__358\ : IoInMux
    port map (
            O => \N__4089\,
            I => \N__4086\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__4086\,
            I => \N__4083\
        );

    \I__356\ : IoSpan4Mux
    port map (
            O => \N__4083\,
            I => \N__4080\
        );

    \I__355\ : Span4Mux_s2_v
    port map (
            O => \N__4080\,
            I => \N__4077\
        );

    \I__354\ : Sp12to4
    port map (
            O => \N__4077\,
            I => \N__4074\
        );

    \I__353\ : Span12Mux_v
    port map (
            O => \N__4074\,
            I => \N__4071\
        );

    \I__352\ : Odrv12
    port map (
            O => \N__4071\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__4314\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__4317\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__4318\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__4313\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__4315\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__4316\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__4319\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6962\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7959\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4152\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7011\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9042\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7499\,
            lcout => \DBRn_c_i\,
            ltout => \DBRn_c_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4155\,
            in3 => \N__10293\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_A20_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__10416\,
            in1 => \N__10629\,
            in2 => \N__4137\,
            in3 => \N__5210\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__10254\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10292\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4224\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.RAM_CYCLE_RNILITE_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__5272\,
            in1 => \N__4103\,
            in2 => \_gnd_net_\,
            in3 => \N__7396\,
            lcout => \U712_CYCLE_TERM_TCIn_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.RAM_CYCLE_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__8516\,
            in1 => \N__4248\,
            in2 => \N__4104\,
            in3 => \N__7442\,
            lcout => \U712_CYCLE_TERM.RAM_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__9932\,
            in1 => \N__11216\,
            in2 => \_gnd_net_\,
            in3 => \N__6774\,
            lcout => \U712_CHIP_RAM.CLK_EN_6_0_a3_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8097\,
            in2 => \_gnd_net_\,
            in3 => \N__7898\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_486_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011100100"
        )
    port map (
            in0 => \N__8518\,
            in1 => \N__10117\,
            in2 => \N__4209\,
            in3 => \N__5673\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9035\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4206\,
            in1 => \N__5334\,
            in2 => \N__6186\,
            in3 => \N__6101\,
            lcout => \U712_CHIP_RAM.CLK_EN_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_i_i_a2_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__10130\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9946\,
            lcout => \N_490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6903\,
            in1 => \N__6294\,
            in2 => \_gnd_net_\,
            in3 => \N__6003\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9019\,
            ce => \N__4188\,
            sr => \N__10255\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6766\,
            in1 => \N__6579\,
            in2 => \_gnd_net_\,
            in3 => \N__8628\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_554_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOJRU2_1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__4232\,
            in1 => \N__6657\,
            in2 => \N__4176\,
            in3 => \N__5380\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4173\,
            in3 => \N__5180\,
            lcout => \U712_CHIP_RAM.N_522\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__11213\,
            in1 => \N__6765\,
            in2 => \_gnd_net_\,
            in3 => \N__6578\,
            lcout => \U712_CHIP_RAM.N_373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6767\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8431\,
            lcout => \U712_CHIP_RAM.N_560\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8430\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5557\,
            lcout => \U712_CHIP_RAM.N_572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__4218\,
            in1 => \N__11214\,
            in2 => \N__4371\,
            in3 => \N__8432\,
            lcout => \WRITE_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9023\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__4233\,
            in1 => \N__5522\,
            in2 => \N__4353\,
            in3 => \N__6658\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__4395\,
            in1 => \N__8482\,
            in2 => \N__4905\,
            in3 => \N__4370\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9027\,
            ce => \N__4863\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_0_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11215\,
            in1 => \N__6768\,
            in2 => \_gnd_net_\,
            in3 => \N__6594\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNIDG0M2_4_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101110"
        )
    port map (
            in0 => \N__4611\,
            in1 => \N__4278\,
            in2 => \N__6323\,
            in3 => \N__4263\,
            lcout => \U712_CYCLE_TERM.un13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6901\,
            in2 => \_gnd_net_\,
            in3 => \N__6243\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9032\,
            ce => \N__4470\,
            sr => \N__10243\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8620\,
            in2 => \_gnd_net_\,
            in3 => \N__5393\,
            lcout => \U712_CHIP_RAM.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__10068\,
            in1 => \N__5747\,
            in2 => \_gnd_net_\,
            in3 => \N__6900\,
            lcout => \U712_CHIP_RAM.N_409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4284\,
            in1 => \N__11231\,
            in2 => \_gnd_net_\,
            in3 => \N__6807\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6177\,
            in1 => \N__6102\,
            in2 => \N__4287\,
            in3 => \N__5396\,
            lcout => \U712_CHIP_RAM.N_504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_0_a2_1_0_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4629\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5777\,
            lcout => \U712_CYCLE_TERM.N_565\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_5_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__9895\,
            in1 => \N__6690\,
            in2 => \_gnd_net_\,
            in3 => \N__6595\,
            lcout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNI05SV_3_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6340\,
            in2 => \_gnd_net_\,
            in3 => \N__5310\,
            lcout => \U712_CYCLE_TERM.N_407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4606\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8517\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9036\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101000001010100"
        )
    port map (
            in0 => \N__4607\,
            in1 => \N__4277\,
            in2 => \N__6324\,
            in3 => \N__4262\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9038\,
            ce => 'H',
            sr => \N__10231\
        );

    \U712_CYCLE_TERM.RAM_CYCLE_RNO_0_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4652\,
            in2 => \_gnd_net_\,
            in3 => \N__4630\,
            lcout => \U712_CYCLE_TERM.N_534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4713\,
            in2 => \_gnd_net_\,
            in3 => \N__4239\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__4320\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4740\,
            in2 => \_gnd_net_\,
            in3 => \N__4236\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__4320\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4752\,
            in2 => \_gnd_net_\,
            in3 => \N__4338\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__4320\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6377\,
            in2 => \_gnd_net_\,
            in3 => \N__4335\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__4320\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4727\,
            in2 => \_gnd_net_\,
            in3 => \N__4332\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__4320\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4797\,
            in2 => \_gnd_net_\,
            in3 => \N__4329\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__4320\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4809\,
            in2 => \_gnd_net_\,
            in3 => \N__4326\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__4320\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4821\,
            in2 => \_gnd_net_\,
            in3 => \N__4323\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4320\,
            ce => 'H',
            sr => \N__5922\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001001000100"
        )
    port map (
            in0 => \N__6806\,
            in1 => \N__5394\,
            in2 => \N__6692\,
            in3 => \N__6566\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_371_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_4_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6164\,
            in1 => \N__6022\,
            in2 => \N__4290\,
            in3 => \N__6094\,
            lcout => \U712_CHIP_RAM.N_519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__8520\,
            in1 => \_gnd_net_\,
            in2 => \N__5153\,
            in3 => \N__4830\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5009\,
            in1 => \N__5517\,
            in2 => \N__6587\,
            in3 => \N__6687\,
            lcout => \U712_CHIP_RAM.N_516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_1_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010000000"
        )
    port map (
            in0 => \N__8519\,
            in1 => \N__5395\,
            in2 => \N__6693\,
            in3 => \N__6567\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIR9VE1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6897\,
            in2 => \_gnd_net_\,
            in3 => \N__6293\,
            lcout => \U712_CHIP_RAM.N_375\,
            ltout => \U712_CHIP_RAM.N_375_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIPCS25_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4374\,
            in3 => \N__6238\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__5556\,
            in1 => \N__8427\,
            in2 => \N__6808\,
            in3 => \N__4842\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9020\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6896\,
            in1 => \N__6286\,
            in2 => \_gnd_net_\,
            in3 => \N__6227\,
            lcout => \U712_CHIP_RAM.N_498\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__5990\,
            in1 => \N__6028\,
            in2 => \N__6178\,
            in3 => \N__6201\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6144\,
            in1 => \N__5555\,
            in2 => \_gnd_net_\,
            in3 => \N__6075\,
            lcout => \U712_CHIP_RAM.N_547\,
            ltout => \U712_CHIP_RAM.N_547_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_4_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__5005\,
            in1 => \N__4841\,
            in2 => \N__4344\,
            in3 => \N__5049\,
            lcout => \U712_CHIP_RAM.N_501\,
            ltout => \U712_CHIP_RAM.N_501_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIG9KPG_2_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__8428\,
            in1 => \N__5145\,
            in2 => \N__4341\,
            in3 => \N__5991\,
            lcout => \U712_CHIP_RAM.N_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVTLS1_7_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6076\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8429\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIE24B8_2_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__5050\,
            in1 => \N__4955\,
            in2 => \N__4401\,
            in3 => \N__6785\,
            lcout => \U712_CHIP_RAM.N_515\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_cry_c_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6571\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4895\,
            in1 => \N__5386\,
            in2 => \_gnd_net_\,
            in3 => \N__4398\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__9024\,
            ce => \N__4861\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6784\,
            in2 => \_gnd_net_\,
            in3 => \N__4389\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4896\,
            in1 => \N__6678\,
            in2 => \_gnd_net_\,
            in3 => \N__4386\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__9024\,
            ce => \N__4861\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4903\,
            in1 => \N__6163\,
            in2 => \_gnd_net_\,
            in3 => \N__4383\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__9024\,
            ce => \N__4861\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4897\,
            in1 => \N__5067\,
            in2 => \_gnd_net_\,
            in3 => \N__4380\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__9024\,
            ce => \N__4861\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4904\,
            in1 => \N__5079\,
            in2 => \_gnd_net_\,
            in3 => \N__4377\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__9024\,
            ce => \N__4861\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4898\,
            in1 => \N__5091\,
            in2 => \_gnd_net_\,
            in3 => \N__4482\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9024\,
            ce => \N__4861\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6146\,
            in1 => \N__5330\,
            in2 => \N__5562\,
            in3 => \N__6080\,
            lcout => \U712_CHIP_RAM.N_666\,
            ltout => \U712_CHIP_RAM.N_666_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNIJH788_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__6810\,
            in1 => \N__8618\,
            in2 => \N__4479\,
            in3 => \N__5714\,
            lcout => \U712_CHIP_RAM.N_393\,
            ltout => \U712_CHIP_RAM.N_393_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIFS4TD_2_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6811\,
            in2 => \N__4476\,
            in3 => \N__5152\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4473\,
            in3 => \N__10290\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__8619\,
            in1 => \N__6812\,
            in2 => \_gnd_net_\,
            in3 => \N__5580\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101111101010000"
        )
    port map (
            in0 => \N__4455\,
            in1 => \_gnd_net_\,
            in2 => \N__4446\,
            in3 => \N__4424\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9028\,
            ce => 'H',
            sr => \N__10236\
        );

    \U712_CHIP_RAM.DBENn_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010111011101110"
        )
    port map (
            in0 => \N__8679\,
            in1 => \N__4413\,
            in2 => \N__6002\,
            in3 => \N__9516\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9028\,
            ce => 'H',
            sr => \N__10236\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101010"
        )
    port map (
            in0 => \N__4407\,
            in1 => \N__11235\,
            in2 => \N__5400\,
            in3 => \N__9964\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9033\,
            ce => \N__5592\,
            sr => \N__10232\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001111"
        )
    port map (
            in0 => \N__4632\,
            in1 => \N__5773\,
            in2 => \N__5318\,
            in3 => \N__4651\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_539_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__8047\,
            in1 => \N__4653\,
            in2 => \N__4656\,
            in3 => \N__8521\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__4650\,
            in1 => \N__5772\,
            in2 => \_gnd_net_\,
            in3 => \N__4631\,
            lcout => \U712_CYCLE_TERM.TACK_EN_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__8522\,
            in1 => \_gnd_net_\,
            in2 => \N__5319\,
            in3 => \N__8048\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4587\,
            in1 => \N__4566\,
            in2 => \_gnd_net_\,
            in3 => \N__9739\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4548\,
            in1 => \N__4533\,
            in2 => \_gnd_net_\,
            in3 => \N__9740\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9741\,
            in1 => \N__9965\,
            in2 => \N__4518\,
            in3 => \N__7920\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4515\,
            in1 => \N__4497\,
            in2 => \_gnd_net_\,
            in3 => \N__9742\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9743\,
            in1 => \N__9950\,
            in2 => \N__4824\,
            in3 => \N__7935\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4820\,
            in1 => \N__4808\,
            in2 => \_gnd_net_\,
            in3 => \N__4796\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4785\,
            in1 => \N__4770\,
            in2 => \_gnd_net_\,
            in3 => \N__9698\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__4751\,
            in1 => \N__4739\,
            in2 => \N__4728\,
            in3 => \N__4712\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4701\,
            in1 => \N__4683\,
            in2 => \_gnd_net_\,
            in3 => \N__9697\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5523\,
            in1 => \N__6688\,
            in2 => \_gnd_net_\,
            in3 => \N__5019\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_669_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001011"
        )
    port map (
            in0 => \N__7216\,
            in1 => \N__5834\,
            in2 => \N__4662\,
            in3 => \N__4974\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9012\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5183\,
            in1 => \N__6689\,
            in2 => \N__6597\,
            in3 => \N__5018\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_520_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110100000001"
        )
    port map (
            in0 => \N__4944\,
            in1 => \N__5833\,
            in2 => \N__4659\,
            in3 => \N__9738\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9012\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__11242\,
            in1 => \N__5017\,
            in2 => \N__6596\,
            in3 => \N__5518\,
            lcout => \U712_CHIP_RAM.N_517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__6200\,
            in1 => \N__5182\,
            in2 => \N__4989\,
            in3 => \N__4980\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000001"
        )
    port map (
            in0 => \N__4973\,
            in1 => \N__4965\,
            in2 => \N__4959\,
            in3 => \N__7120\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9012\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__6435\,
            in1 => \N__4956\,
            in2 => \N__6902\,
            in3 => \N__6239\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101011010"
        )
    port map (
            in0 => \N__4928\,
            in1 => \N__4911\,
            in2 => \N__6577\,
            in3 => \N__4902\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9015\,
            ce => \N__4862\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_1_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5376\,
            in1 => \N__6651\,
            in2 => \_gnd_net_\,
            in3 => \N__6546\,
            lcout => \U712_CHIP_RAM.N_549\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_0_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6547\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6659\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_559_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_4_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5377\,
            in1 => \N__6147\,
            in2 => \N__4845\,
            in3 => \N__6081\,
            lcout => \U712_CHIP_RAM.N_665\,
            ltout => \U712_CHIP_RAM.N_665_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__6813\,
            in1 => \N__5181\,
            in2 => \N__4833\,
            in3 => \N__5052\,
            lcout => \U712_CHIP_RAM.N_471\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6277\,
            in1 => \N__6898\,
            in2 => \_gnd_net_\,
            in3 => \N__5988\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_2_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__10624\,
            in1 => \_gnd_net_\,
            in2 => \N__5232\,
            in3 => \N__5229\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_1_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__6881\,
            in1 => \N__5989\,
            in2 => \N__5214\,
            in3 => \N__5211\,
            lcout => \U712_CHIP_RAM.BANK0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_2_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6790\,
            in1 => \N__6082\,
            in2 => \_gnd_net_\,
            in3 => \N__5042\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_0_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5196\,
            in1 => \N__6791\,
            in2 => \N__5051\,
            in3 => \N__5184\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_523_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__5102\,
            in1 => \N__5157\,
            in2 => \N__5121\,
            in3 => \N__5118\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9021\,
            ce => 'H',
            sr => \N__10237\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5090\,
            in1 => \N__5078\,
            in2 => \_gnd_net_\,
            in3 => \N__5066\,
            lcout => \U712_CHIP_RAM.N_545\,
            ltout => \U712_CHIP_RAM.N_545_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5548\,
            in1 => \N__6789\,
            in2 => \N__5055\,
            in3 => \N__5041\,
            lcout => \U712_CHIP_RAM.N_562\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__5462\,
            in1 => \N__5503\,
            in2 => \N__6680\,
            in3 => \N__5568\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10289\,
            in1 => \_gnd_net_\,
            in2 => \N__5595\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__6653\,
            in1 => \N__5579\,
            in2 => \N__5516\,
            in3 => \N__6809\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5379\,
            in1 => \N__6145\,
            in2 => \N__6093\,
            in3 => \N__5558\,
            lcout => \U712_CHIP_RAM.N_557\,
            ltout => \U712_CHIP_RAM.N_557_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__5469\,
            in1 => \N__5463\,
            in2 => \N__5442\,
            in3 => \N__6679\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010101000"
        )
    port map (
            in0 => \N__8505\,
            in1 => \N__5411\,
            in2 => \N__5439\,
            in3 => \N__5436\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9025\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_1_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6652\,
            in1 => \N__5378\,
            in2 => \_gnd_net_\,
            in3 => \N__6586\,
            lcout => \U712_CHIP_RAM.N_566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6861\,
            in2 => \_gnd_net_\,
            in3 => \N__6226\,
            lcout => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__5253\,
            in1 => \N__6350\,
            in2 => \N__8049\,
            in3 => \N__5317\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9029\,
            ce => 'H',
            sr => \N__10228\
        );

    \U712_REG_SM.ASn_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__7017\,
            in1 => \N__8194\,
            in2 => \N__7728\,
            in3 => \N__5791\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9029\,
            ce => 'H',
            sr => \N__10228\
        );

    \U712_REG_SM.REG_TACK_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__7880\,
            in1 => \N__5652\,
            in2 => \N__5778\,
            in3 => \N__5658\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9029\,
            ce => 'H',
            sr => \N__10228\
        );

    \U712_CHIP_RAM.DBDIR_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__5748\,
            in1 => \N__5684\,
            in2 => \_gnd_net_\,
            in3 => \N__5715\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9029\,
            ce => 'H',
            sr => \N__10228\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__8124\,
            in1 => \N__7688\,
            in2 => \_gnd_net_\,
            in3 => \N__8178\,
            lcout => \U712_REG_SM.N_447\,
            ltout => \U712_REG_SM.N_447_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__10082\,
            in1 => \_gnd_net_\,
            in2 => \N__5661\,
            in3 => \N__7778\,
            lcout => \U712_REG_SM.REG_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__7779\,
            in1 => \N__7689\,
            in2 => \_gnd_net_\,
            in3 => \N__8179\,
            lcout => \U712_REG_SM.N_478\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5928\,
            in1 => \N__5934\,
            in2 => \_gnd_net_\,
            in3 => \N__5943\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9001\,
            ce => \N__8891\,
            sr => \N__10256\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__9095\,
            in1 => \N__10641\,
            in2 => \N__9192\,
            in3 => \N__5622\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9001\,
            ce => \N__8891\,
            sr => \N__10256\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__10291\,
            in1 => \N__5910\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__9953\,
            in1 => \N__5949\,
            in2 => \N__9612\,
            in3 => \N__9759\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7113\,
            in2 => \_gnd_net_\,
            in3 => \N__7065\,
            lcout => \U712_CHIP_RAM.N_379\,
            ltout => \U712_CHIP_RAM.N_379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001111"
        )
    port map (
            in0 => \N__9951\,
            in1 => \N__8858\,
            in2 => \N__5937\,
            in3 => \N__9758\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110001111"
        )
    port map (
            in0 => \N__8859\,
            in1 => \N__9094\,
            in2 => \N__9779\,
            in3 => \N__9952\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9694\,
            in1 => \N__7052\,
            in2 => \N__7212\,
            in3 => \N__7099\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => \U712_CHIP_RAM.REFRESH_RST_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__9695\,
            in1 => \N__7202\,
            in2 => \N__5913\,
            in3 => \N__7100\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9696\,
            in1 => \N__5891\,
            in2 => \_gnd_net_\,
            in3 => \N__5862\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__5841\,
            in1 => \N__5835\,
            in2 => \N__7070\,
            in3 => \N__5958\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9009\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8515\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6261\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6422\,
            in1 => \N__6399\,
            in2 => \_gnd_net_\,
            in3 => \N__9717\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010110000"
        )
    port map (
            in0 => \N__6381\,
            in1 => \N__6363\,
            in2 => \N__8523\,
            in3 => \N__6357\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9009\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8426\,
            in2 => \_gnd_net_\,
            in3 => \N__6351\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9013\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6259\,
            in1 => \N__6457\,
            in2 => \_gnd_net_\,
            in3 => \N__7797\,
            lcout => \U712_CHIP_RAM.N_567\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIHSHE1_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__8425\,
            in1 => \N__6862\,
            in2 => \_gnd_net_\,
            in3 => \N__6260\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__7808\,
            in1 => \N__6458\,
            in2 => \N__6246\,
            in3 => \N__6228\,
            lcout => \U712_CHIP_RAM.N_502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6029\,
            in1 => \N__6498\,
            in2 => \N__6185\,
            in3 => \N__6092\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_518_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6030\,
            in2 => \N__6006\,
            in3 => \N__5992\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011111000"
        )
    port map (
            in0 => \N__8541\,
            in1 => \N__8504\,
            in2 => \N__6899\,
            in3 => \N__8640\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6792\,
            in1 => \N__6691\,
            in2 => \_gnd_net_\,
            in3 => \N__6565\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9938\,
            in2 => \_gnd_net_\,
            in3 => \N__6459\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_492_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__6492\,
            in1 => \N__7640\,
            in2 => \N__6462\,
            in3 => \N__8503\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7839\,
            in1 => \N__7770\,
            in2 => \_gnd_net_\,
            in3 => \N__8132\,
            lcout => OPEN,
            ltout => \U712_REG_SM.STATE_COUNT_srsts_i_0_0_a2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011110001"
        )
    port map (
            in0 => \N__7771\,
            in1 => \N__6441\,
            in2 => \N__6444\,
            in3 => \N__7881\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9022\,
            ce => 'H',
            sr => \N__10229\
        );

    \U712_REG_SM.C3_SYNC_RNI347S_1_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7701\,
            in1 => \N__8195\,
            in2 => \_gnd_net_\,
            in3 => \N__7807\,
            lcout => \U712_REG_SM.N_661\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__10072\,
            in1 => \N__8089\,
            in2 => \_gnd_net_\,
            in3 => \N__8127\,
            lcout => \U712_REG_SM.DS_EN_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__8125\,
            in1 => \N__7695\,
            in2 => \_gnd_net_\,
            in3 => \N__8188\,
            lcout => \U712_REG_SM.N_374\,
            ltout => \U712_REG_SM.N_374_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__8506\,
            in1 => \N__7772\,
            in2 => \N__7020\,
            in3 => \N__8128\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9026\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8088\,
            in2 => \_gnd_net_\,
            in3 => \N__8224\,
            lcout => \U712_REG_SM.N_389\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_RNO_0_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8187\,
            in1 => \N__8225\,
            in2 => \_gnd_net_\,
            in3 => \N__8126\,
            lcout => \U712_REG_SM.N_417\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_1_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6927\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9030\,
            ce => 'H',
            sr => \N__10226\
        );

    \U712_REG_SM.C3_SYNC_0_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6992\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9030\,
            ce => 'H',
            sr => \N__10226\
        );

    \U712_REG_SM.DS_EN_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100000001"
        )
    port map (
            in0 => \N__7647\,
            in1 => \N__6975\,
            in2 => \N__8058\,
            in3 => \N__11054\,
            lcout => \DS_ENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9030\,
            ce => 'H',
            sr => \N__10226\
        );

    \U712_REG_SM.C3_SYNC_1_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6969\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9030\,
            ce => 'H',
            sr => \N__10226\
        );

    \U712_REG_SM.C1_SYNC_0_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6963\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9034\,
            ce => 'H',
            sr => \N__10225\
        );

    \U712_CHIP_RAM.RASn_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7128\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8997\,
            ce => 'H',
            sr => \N__10270\
        );

    \U712_CHIP_RAM.WEn_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7071\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8998\,
            ce => 'H',
            sr => \N__10253\
        );

    \U712_CHIP_RAM.CRCSn_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7221\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8998\,
            ce => 'H',
            sr => \N__10253\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__7029\,
            in1 => \N__10374\,
            in2 => \N__9975\,
            in3 => \N__7314\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8999\,
            ce => \N__8912\,
            sr => \N__10247\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__7028\,
            in1 => \N__7272\,
            in2 => \N__9974\,
            in3 => \N__7947\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8999\,
            ce => \N__8912\,
            sr => \N__10247\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__9121\,
            in1 => \N__7545\,
            in2 => \N__9789\,
            in3 => \N__7515\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8999\,
            ce => \N__8912\,
            sr => \N__10247\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__9782\,
            in1 => \_gnd_net_\,
            in2 => \N__9131\,
            in3 => \N__7220\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8999\,
            ce => \N__8912\,
            sr => \N__10247\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__7941\,
            in1 => \N__9125\,
            in2 => \N__9193\,
            in3 => \N__7134\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8999\,
            ce => \N__8912\,
            sr => \N__10247\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__7140\,
            in1 => \N__9781\,
            in2 => \N__9967\,
            in3 => \N__8550\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__7121\,
            in1 => \N__9780\,
            in2 => \_gnd_net_\,
            in3 => \N__7066\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7470\,
            in2 => \_gnd_net_\,
            in3 => \N__7831\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_477_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__8497\,
            in1 => \N__7641\,
            in2 => \N__7611\,
            in3 => \N__7608\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9004\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7577\,
            in1 => \N__9936\,
            in2 => \_gnd_net_\,
            in3 => \N__8772\,
            lcout => \U712_CHIP_RAM.N_422\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7536\,
            in1 => \N__9937\,
            in2 => \_gnd_net_\,
            in3 => \N__7926\,
            lcout => \U712_CHIP_RAM.N_445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_0_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7506\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9005\,
            ce => 'H',
            sr => \N__10230\
        );

    \DBR_SYNC_1_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7476\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9005\,
            ce => 'H',
            sr => \N__10230\
        );

    \U712_REG_SM.START_RST_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__7469\,
            in1 => \N__7742\,
            in2 => \_gnd_net_\,
            in3 => \N__8232\,
            lcout => \U712_REG_SM.START_RSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9011\,
            ce => 'H',
            sr => \N__10227\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__7372\,
            in1 => \N__7455\,
            in2 => \_gnd_net_\,
            in3 => \N__7443\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9011\,
            ce => 'H',
            sr => \N__10227\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8093\,
            in2 => \N__7724\,
            in3 => \N__8197\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_475_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__7899\,
            in1 => \N__7879\,
            in2 => \N__7863\,
            in3 => \N__8494\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9014\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_57_i_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000101"
        )
    port map (
            in0 => \N__8565\,
            in1 => \N__11174\,
            in2 => \N__8662\,
            in3 => \N__8689\,
            lcout => \N_57_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7838\,
            in1 => \N__8196\,
            in2 => \N__7723\,
            in3 => \N__7818\,
            lcout => \U712_REG_SM.START_RST_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101110111011"
        )
    port map (
            in0 => \N__8094\,
            in1 => \N__7769\,
            in2 => \N__7812\,
            in3 => \N__7716\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_449_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__8495\,
            in1 => \N__7712\,
            in2 => \N__7782\,
            in3 => \N__8198\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9014\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7700\,
            in2 => \_gnd_net_\,
            in3 => \N__8193\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_396_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__8231\,
            in1 => \N__7743\,
            in2 => \N__7731\,
            in3 => \N__8496\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_2_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__8095\,
            in1 => \N__8226\,
            in2 => \N__8199\,
            in3 => \N__7696\,
            lcout => \U712_REG_SM.un1_STATE_COUNT_4_i_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__8227\,
            in1 => \N__8192\,
            in2 => \N__8133\,
            in3 => \N__8096\,
            lcout => \U712_REG_SM.N_479\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_RNI8MQ3_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8043\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8481\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10736\,
            in1 => \_gnd_net_\,
            in2 => \N__10623\,
            in3 => \N__10434\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10365\,
            ce => \N__10331\,
            sr => \N__10257\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10603\,
            in1 => \N__8280\,
            in2 => \_gnd_net_\,
            in3 => \N__8820\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10365\,
            ce => \N__10331\,
            sr => \N__10257\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9435\,
            in1 => \N__10602\,
            in2 => \_gnd_net_\,
            in3 => \N__9387\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__10330\,
            sr => \N__10248\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8816\,
            in1 => \N__10598\,
            in2 => \_gnd_net_\,
            in3 => \N__8279\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10329\,
            sr => \N__10245\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10728\,
            in1 => \N__10599\,
            in2 => \_gnd_net_\,
            in3 => \N__10429\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__10329\,
            sr => \N__10245\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9745\,
            in1 => \N__7908\,
            in2 => \N__9959\,
            in3 => \N__8556\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9744\,
            in2 => \_gnd_net_\,
            in3 => \N__9918\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9588\,
            in1 => \N__10608\,
            in2 => \_gnd_net_\,
            in3 => \N__8809\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10326\,
            sr => \N__10238\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9382\,
            in1 => \N__10609\,
            in2 => \_gnd_net_\,
            in3 => \N__8272\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10326\,
            sr => \N__10238\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__8492\,
            in1 => \N__10029\,
            in2 => \_gnd_net_\,
            in3 => \N__11170\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8331\,
            in2 => \_gnd_net_\,
            in3 => \N__8531\,
            lcout => \U712_CHIP_RAM.un3_DMA_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8532\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8493\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9945\,
            in1 => \N__8325\,
            in2 => \N__9787\,
            in3 => \N__9627\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__9112\,
            in1 => \N__8238\,
            in2 => \N__9194\,
            in3 => \N__8313\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9002\,
            ce => \N__8908\,
            sr => \N__10260\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9386\,
            in1 => \N__10600\,
            in2 => \_gnd_net_\,
            in3 => \N__8271\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10364\,
            ce => \N__10332\,
            sr => \N__10258\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10601\,
            in1 => \N__9495\,
            in2 => \_gnd_net_\,
            in3 => \N__9431\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10364\,
            ce => \N__10332\,
            sr => \N__10258\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__9132\,
            in1 => \N__9597\,
            in2 => \N__9173\,
            in3 => \N__8847\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9010\,
            ce => \N__8907\,
            sr => \N__10249\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9587\,
            in1 => \N__10545\,
            in2 => \_gnd_net_\,
            in3 => \N__8795\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10363\,
            ce => \N__10327\,
            sr => \N__10244\
        );

    \U712_BYTE_ENABLE.N_295_i_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__8574\,
            in1 => \N__8706\,
            in2 => \N__10028\,
            in3 => \N__8655\,
            lcout => \N_295_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_299_i_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100011"
        )
    port map (
            in0 => \N__10024\,
            in1 => \N__9309\,
            in2 => \N__8664\,
            in3 => \N__8708\,
            lcout => \N_299_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_297_i_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__8707\,
            in1 => \N__9315\,
            in2 => \N__8663\,
            in3 => \N__11169\,
            lcout => \N_297_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000101010"
        )
    port map (
            in0 => \N__9963\,
            in1 => \N__10950\,
            in2 => \N__9300\,
            in3 => \N__10873\,
            lcout => \U712_BYTE_ENABLE.N_528\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_o2_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10874\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10781\,
            lcout => \U712_BYTE_ENABLE.N_377\,
            ltout => \U712_BYTE_ENABLE.N_377_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010101010"
        )
    port map (
            in0 => \N__9961\,
            in1 => \N__10948\,
            in2 => \N__8568\,
            in3 => \N__9295\,
            lcout => \U712_BYTE_ENABLE.N_508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010101010"
        )
    port map (
            in0 => \N__9962\,
            in1 => \N__10949\,
            in2 => \N__9324\,
            in3 => \N__9296\,
            lcout => \U712_BYTE_ENABLE.N_530\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000000"
        )
    port map (
            in0 => \N__9294\,
            in1 => \N__10947\,
            in2 => \N__10882\,
            in3 => \N__9966\,
            lcout => \U712_BYTE_ENABLE.N_532\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_i_x2_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11023\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10780\,
            lcout => \U712_BYTE_ENABLE.N_364_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DMA_LATCH_EN_0_a2_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__10020\,
            in1 => \N__11178\,
            in2 => \_gnd_net_\,
            in3 => \N__11255\,
            lcout => \DMA_LATCH_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_403_i_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011100000"
        )
    port map (
            in0 => \N__10935\,
            in1 => \N__10883\,
            in2 => \N__11014\,
            in3 => \N__10779\,
            lcout => \N_403_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9788\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9000\,
            ce => 'H',
            sr => \N__10272\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__9333\,
            in1 => \N__9127\,
            in2 => \N__9195\,
            in3 => \N__9633\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9003\,
            ce => \N__8913\,
            sr => \N__10269\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__9191\,
            in1 => \N__9126\,
            in2 => \N__9447\,
            in3 => \N__9069\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9003\,
            ce => \N__8913\,
            sr => \N__10269\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9960\,
            in1 => \N__9798\,
            in2 => \N__9786\,
            in3 => \N__9618\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10611\,
            in1 => \N__10737\,
            in2 => \_gnd_net_\,
            in3 => \N__10685\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__10335\,
            sr => \N__10261\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10612\,
            in1 => \N__9494\,
            in2 => \_gnd_net_\,
            in3 => \N__9430\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__10335\,
            sr => \N__10261\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10684\,
            in1 => \N__10610\,
            in2 => \_gnd_net_\,
            in3 => \N__9486\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__10333\,
            sr => \N__10259\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9543\,
            in1 => \N__10572\,
            in2 => \_gnd_net_\,
            in3 => \N__9586\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10360\,
            ce => \N__10328\,
            sr => \N__10246\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9582\,
            in1 => \N__10607\,
            in2 => \_gnd_net_\,
            in3 => \N__9539\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10334\,
            sr => \N__10239\
        );

    \U712_BYTE_ENABLE.N_402_i_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111010000"
        )
    port map (
            in0 => \N__10936\,
            in1 => \N__10884\,
            in2 => \N__11024\,
            in3 => \N__10802\,
            lcout => \N_402_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9493\,
            in1 => \_gnd_net_\,
            in2 => \N__10628\,
            in3 => \N__10680\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10361\,
            ce => \N__10336\,
            sr => \N__10268\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10619\,
            in1 => \N__9429\,
            in2 => \_gnd_net_\,
            in3 => \N__9369\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10361\,
            ce => \N__10336\,
            sr => \N__10268\
        );

    \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100011111111"
        )
    port map (
            in0 => \N__10864\,
            in1 => \N__10986\,
            in2 => \N__10815\,
            in3 => \N__11069\,
            lcout => \N_291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_400_i_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110100000"
        )
    port map (
            in0 => \N__10933\,
            in1 => \N__10865\,
            in2 => \N__10811\,
            in3 => \N__11018\,
            lcout => \N_400_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011111111"
        )
    port map (
            in0 => \N__10869\,
            in1 => \N__10807\,
            in2 => \N__11025\,
            in3 => \N__11073\,
            lcout => \N_293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_401_i_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100101010"
        )
    port map (
            in0 => \N__11019\,
            in1 => \N__10934\,
            in2 => \N__10881\,
            in3 => \N__10806\,
            lcout => \N_401_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10550\,
            in1 => \N__10729\,
            in2 => \_gnd_net_\,
            in3 => \N__10686\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10362\,
            ce => \N__10337\,
            sr => \N__10271\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10549\,
            in1 => \N__10449\,
            in2 => \_gnd_net_\,
            in3 => \N__10433\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10359\,
            ce => \N__10338\,
            sr => \N__10273\
        );

    \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000100000"
        )
    port map (
            in0 => \N__11156\,
            in1 => \N__10140\,
            in2 => \N__10019\,
            in3 => \_gnd_net_\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_0_m2_LC_24_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100001111"
        )
    port map (
            in0 => \N__10086\,
            in1 => \N__10004\,
            in2 => \N__11262\,
            in3 => \N__11155\,
            lcout => \N_450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
